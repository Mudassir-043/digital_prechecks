magic
tech sky130B
magscale 1 2
timestamp 1667543118
<< locali >>
rect -5892 9472 28954 10488
rect -5892 8532 28978 9472
rect -5818 -7669 -3777 8532
rect -2834 7181 25461 7315
rect -2834 6715 285 7181
rect 5863 7155 25461 7181
rect 5863 6761 16853 7155
rect 21927 6761 25461 7155
rect 5863 6715 25461 6761
rect -2834 6609 25461 6715
rect -5831 -10604 -3752 -7669
rect -2834 -8378 -717 6609
rect 152 6204 6039 6224
rect 152 6170 162 6204
rect 196 6170 234 6204
rect 268 6170 306 6204
rect 340 6170 378 6204
rect 412 6170 450 6204
rect 484 6170 522 6204
rect 556 6170 594 6204
rect 628 6170 666 6204
rect 700 6170 738 6204
rect 772 6170 810 6204
rect 844 6170 882 6204
rect 916 6170 954 6204
rect 988 6170 1026 6204
rect 1060 6170 1098 6204
rect 1132 6170 1170 6204
rect 1204 6170 1242 6204
rect 1276 6170 1314 6204
rect 1348 6170 1386 6204
rect 1420 6170 1458 6204
rect 1492 6170 1530 6204
rect 1564 6170 1602 6204
rect 1636 6170 1674 6204
rect 1708 6170 1746 6204
rect 1780 6170 1818 6204
rect 1852 6170 1890 6204
rect 1924 6170 1962 6204
rect 1996 6170 2034 6204
rect 2068 6170 2106 6204
rect 2140 6170 2178 6204
rect 2212 6170 2250 6204
rect 2284 6170 2322 6204
rect 2356 6170 2394 6204
rect 2428 6170 2466 6204
rect 2500 6170 2538 6204
rect 2572 6170 2610 6204
rect 2644 6170 2682 6204
rect 2716 6170 2754 6204
rect 2788 6170 2826 6204
rect 2860 6170 2898 6204
rect 2932 6170 2970 6204
rect 3004 6170 3042 6204
rect 3076 6170 3114 6204
rect 3148 6170 3186 6204
rect 3220 6170 3258 6204
rect 3292 6170 3330 6204
rect 3364 6170 3402 6204
rect 3436 6170 3474 6204
rect 3508 6170 3546 6204
rect 3580 6170 3618 6204
rect 3652 6170 3690 6204
rect 3724 6170 3762 6204
rect 3796 6170 3834 6204
rect 3868 6170 3906 6204
rect 3940 6170 3978 6204
rect 4012 6170 4050 6204
rect 4084 6170 4122 6204
rect 4156 6170 4194 6204
rect 4228 6170 4266 6204
rect 4300 6170 4338 6204
rect 4372 6170 4410 6204
rect 4444 6170 4482 6204
rect 4516 6170 4554 6204
rect 4588 6170 4626 6204
rect 4660 6170 4698 6204
rect 4732 6170 4770 6204
rect 4804 6170 4842 6204
rect 4876 6170 4914 6204
rect 4948 6170 4986 6204
rect 5020 6170 5058 6204
rect 5092 6170 5130 6204
rect 5164 6170 5202 6204
rect 5236 6170 5274 6204
rect 5308 6170 5346 6204
rect 5380 6170 5418 6204
rect 5452 6170 5490 6204
rect 5524 6170 5562 6204
rect 5596 6170 5634 6204
rect 5668 6170 5706 6204
rect 5740 6170 5778 6204
rect 5812 6170 5850 6204
rect 5884 6170 5922 6204
rect 5956 6170 5994 6204
rect 6028 6170 6039 6204
rect 152 6150 6039 6170
rect 16426 6207 22162 6225
rect 16426 6173 16433 6207
rect 16467 6173 16505 6207
rect 16539 6173 16577 6207
rect 16611 6173 16649 6207
rect 16683 6173 16721 6207
rect 16755 6173 16793 6207
rect 16827 6173 16865 6207
rect 16899 6173 16937 6207
rect 16971 6173 17009 6207
rect 17043 6173 17081 6207
rect 17115 6173 17153 6207
rect 17187 6173 17225 6207
rect 17259 6173 17297 6207
rect 17331 6173 17369 6207
rect 17403 6173 17441 6207
rect 17475 6173 17513 6207
rect 17547 6173 17585 6207
rect 17619 6173 17657 6207
rect 17691 6173 17729 6207
rect 17763 6173 17801 6207
rect 17835 6173 17873 6207
rect 17907 6173 17945 6207
rect 17979 6173 18017 6207
rect 18051 6173 18089 6207
rect 18123 6173 18161 6207
rect 18195 6173 18233 6207
rect 18267 6173 18305 6207
rect 18339 6173 18377 6207
rect 18411 6173 18449 6207
rect 18483 6173 18521 6207
rect 18555 6173 18593 6207
rect 18627 6173 18665 6207
rect 18699 6173 18737 6207
rect 18771 6173 18809 6207
rect 18843 6173 18881 6207
rect 18915 6173 18953 6207
rect 18987 6173 19025 6207
rect 19059 6173 19097 6207
rect 19131 6173 19169 6207
rect 19203 6173 19241 6207
rect 19275 6173 19313 6207
rect 19347 6173 19385 6207
rect 19419 6173 19457 6207
rect 19491 6173 19529 6207
rect 19563 6173 19601 6207
rect 19635 6173 19673 6207
rect 19707 6173 19745 6207
rect 19779 6173 19817 6207
rect 19851 6173 19889 6207
rect 19923 6173 19961 6207
rect 19995 6173 20033 6207
rect 20067 6173 20105 6207
rect 20139 6173 20177 6207
rect 20211 6173 20249 6207
rect 20283 6173 20321 6207
rect 20355 6173 20393 6207
rect 20427 6173 20465 6207
rect 20499 6173 20537 6207
rect 20571 6173 20609 6207
rect 20643 6173 20681 6207
rect 20715 6173 20753 6207
rect 20787 6173 20825 6207
rect 20859 6173 20897 6207
rect 20931 6173 20969 6207
rect 21003 6173 21041 6207
rect 21075 6173 21113 6207
rect 21147 6173 21185 6207
rect 21219 6173 21257 6207
rect 21291 6173 21329 6207
rect 21363 6173 21401 6207
rect 21435 6173 21473 6207
rect 21507 6173 21545 6207
rect 21579 6173 21617 6207
rect 21651 6173 21689 6207
rect 21723 6173 21761 6207
rect 21795 6173 21833 6207
rect 21867 6173 21905 6207
rect 21939 6173 21977 6207
rect 22011 6173 22049 6207
rect 22083 6173 22121 6207
rect 22155 6173 22162 6207
rect 16426 6155 22162 6173
rect 6297 2269 15884 2538
rect 6297 1227 10568 2269
rect 12258 1227 15884 2269
rect 6297 557 15884 1227
rect 651 -1018 6052 -115
rect 16380 -1045 22087 -125
rect 6272 -4837 15879 -4296
rect 6272 -7031 10086 -4837
rect 11848 -7031 15879 -4837
rect 869 -7325 6010 -7309
rect 869 -7359 902 -7325
rect 936 -7359 974 -7325
rect 1008 -7359 1046 -7325
rect 1080 -7359 1118 -7325
rect 1152 -7359 1190 -7325
rect 1224 -7359 1262 -7325
rect 1296 -7359 1334 -7325
rect 1368 -7359 1406 -7325
rect 1440 -7359 1478 -7325
rect 1512 -7359 1550 -7325
rect 1584 -7359 1622 -7325
rect 1656 -7359 1694 -7325
rect 1728 -7359 1766 -7325
rect 1800 -7359 1838 -7325
rect 1872 -7359 1910 -7325
rect 1944 -7359 1982 -7325
rect 2016 -7359 2054 -7325
rect 2088 -7359 2126 -7325
rect 2160 -7359 2198 -7325
rect 2232 -7359 2270 -7325
rect 2304 -7359 2342 -7325
rect 2376 -7359 2414 -7325
rect 2448 -7359 2486 -7325
rect 2520 -7359 2558 -7325
rect 2592 -7359 2630 -7325
rect 2664 -7359 2702 -7325
rect 2736 -7359 2774 -7325
rect 2808 -7359 2846 -7325
rect 2880 -7359 2918 -7325
rect 2952 -7359 2990 -7325
rect 3024 -7359 3062 -7325
rect 3096 -7359 3134 -7325
rect 3168 -7359 3206 -7325
rect 3240 -7359 3278 -7325
rect 3312 -7359 3350 -7325
rect 3384 -7359 3422 -7325
rect 3456 -7359 3494 -7325
rect 3528 -7359 3566 -7325
rect 3600 -7359 3638 -7325
rect 3672 -7359 3710 -7325
rect 3744 -7359 3782 -7325
rect 3816 -7359 3854 -7325
rect 3888 -7359 3926 -7325
rect 3960 -7359 3998 -7325
rect 4032 -7359 4070 -7325
rect 4104 -7359 4142 -7325
rect 4176 -7359 4214 -7325
rect 4248 -7359 4286 -7325
rect 4320 -7359 4358 -7325
rect 4392 -7359 4430 -7325
rect 4464 -7359 4502 -7325
rect 4536 -7359 4574 -7325
rect 4608 -7359 4646 -7325
rect 4680 -7359 4718 -7325
rect 4752 -7359 4790 -7325
rect 4824 -7359 4862 -7325
rect 4896 -7359 4934 -7325
rect 4968 -7359 5006 -7325
rect 5040 -7359 5078 -7325
rect 5112 -7359 5150 -7325
rect 5184 -7359 5222 -7325
rect 5256 -7359 5294 -7325
rect 5328 -7359 5366 -7325
rect 5400 -7359 5438 -7325
rect 5472 -7359 5510 -7325
rect 5544 -7359 5582 -7325
rect 5616 -7359 5654 -7325
rect 5688 -7359 5726 -7325
rect 5760 -7359 5798 -7325
rect 5832 -7359 5870 -7325
rect 5904 -7359 5942 -7325
rect 5976 -7359 6010 -7325
rect 869 -7375 6010 -7359
rect 6272 -7406 15879 -7031
rect 16434 -7308 21937 -7305
rect 16434 -7342 16468 -7308
rect 16502 -7342 16540 -7308
rect 16574 -7342 16612 -7308
rect 16646 -7342 16684 -7308
rect 16718 -7342 16756 -7308
rect 16790 -7342 16828 -7308
rect 16862 -7342 16900 -7308
rect 16934 -7342 16972 -7308
rect 17006 -7342 17044 -7308
rect 17078 -7342 17116 -7308
rect 17150 -7342 17188 -7308
rect 17222 -7342 17260 -7308
rect 17294 -7342 17332 -7308
rect 17366 -7342 17404 -7308
rect 17438 -7342 17476 -7308
rect 17510 -7342 17548 -7308
rect 17582 -7342 17620 -7308
rect 17654 -7342 17692 -7308
rect 17726 -7342 17764 -7308
rect 17798 -7342 17836 -7308
rect 17870 -7342 17908 -7308
rect 17942 -7342 17980 -7308
rect 18014 -7342 18052 -7308
rect 18086 -7342 18124 -7308
rect 18158 -7342 18196 -7308
rect 18230 -7342 18268 -7308
rect 18302 -7342 18340 -7308
rect 18374 -7342 18412 -7308
rect 18446 -7342 18484 -7308
rect 18518 -7342 18556 -7308
rect 18590 -7342 18628 -7308
rect 18662 -7342 18700 -7308
rect 18734 -7342 18772 -7308
rect 18806 -7342 18844 -7308
rect 18878 -7342 18916 -7308
rect 18950 -7342 18988 -7308
rect 19022 -7342 19060 -7308
rect 19094 -7342 19132 -7308
rect 19166 -7342 19204 -7308
rect 19238 -7342 19276 -7308
rect 19310 -7342 19348 -7308
rect 19382 -7342 19420 -7308
rect 19454 -7342 19492 -7308
rect 19526 -7342 19564 -7308
rect 19598 -7342 19636 -7308
rect 19670 -7342 19708 -7308
rect 19742 -7342 19780 -7308
rect 19814 -7342 19852 -7308
rect 19886 -7342 19924 -7308
rect 19958 -7342 19996 -7308
rect 20030 -7342 20068 -7308
rect 20102 -7342 20140 -7308
rect 20174 -7342 20212 -7308
rect 20246 -7342 20284 -7308
rect 20318 -7342 20356 -7308
rect 20390 -7342 20428 -7308
rect 20462 -7342 20500 -7308
rect 20534 -7342 20572 -7308
rect 20606 -7342 20644 -7308
rect 20678 -7342 20716 -7308
rect 20750 -7342 20788 -7308
rect 20822 -7342 20860 -7308
rect 20894 -7342 20932 -7308
rect 20966 -7342 21004 -7308
rect 21038 -7342 21076 -7308
rect 21110 -7342 21148 -7308
rect 21182 -7342 21220 -7308
rect 21254 -7342 21292 -7308
rect 21326 -7342 21364 -7308
rect 21398 -7342 21436 -7308
rect 21470 -7342 21508 -7308
rect 21542 -7342 21580 -7308
rect 21614 -7342 21652 -7308
rect 21686 -7342 21724 -7308
rect 21758 -7342 21796 -7308
rect 21830 -7342 21868 -7308
rect 21902 -7342 21937 -7308
rect 16434 -7344 21937 -7342
rect 6292 -7436 15879 -7406
rect 23344 -8378 25461 6609
rect -2835 -8522 25461 -8378
rect -2835 -8588 16582 -8522
rect -2835 -8910 1087 -8588
rect 5729 -8910 16582 -8588
rect -2835 -8988 16582 -8910
rect 21800 -8959 25461 -8522
rect 21800 -8988 25460 -8959
rect -2835 -9084 25460 -8988
rect 26937 -10604 28978 8532
rect -5831 -12560 29015 -10604
<< viali >>
rect 285 6715 5863 7181
rect 16853 6761 21927 7155
rect 162 6170 196 6204
rect 234 6170 268 6204
rect 306 6170 340 6204
rect 378 6170 412 6204
rect 450 6170 484 6204
rect 522 6170 556 6204
rect 594 6170 628 6204
rect 666 6170 700 6204
rect 738 6170 772 6204
rect 810 6170 844 6204
rect 882 6170 916 6204
rect 954 6170 988 6204
rect 1026 6170 1060 6204
rect 1098 6170 1132 6204
rect 1170 6170 1204 6204
rect 1242 6170 1276 6204
rect 1314 6170 1348 6204
rect 1386 6170 1420 6204
rect 1458 6170 1492 6204
rect 1530 6170 1564 6204
rect 1602 6170 1636 6204
rect 1674 6170 1708 6204
rect 1746 6170 1780 6204
rect 1818 6170 1852 6204
rect 1890 6170 1924 6204
rect 1962 6170 1996 6204
rect 2034 6170 2068 6204
rect 2106 6170 2140 6204
rect 2178 6170 2212 6204
rect 2250 6170 2284 6204
rect 2322 6170 2356 6204
rect 2394 6170 2428 6204
rect 2466 6170 2500 6204
rect 2538 6170 2572 6204
rect 2610 6170 2644 6204
rect 2682 6170 2716 6204
rect 2754 6170 2788 6204
rect 2826 6170 2860 6204
rect 2898 6170 2932 6204
rect 2970 6170 3004 6204
rect 3042 6170 3076 6204
rect 3114 6170 3148 6204
rect 3186 6170 3220 6204
rect 3258 6170 3292 6204
rect 3330 6170 3364 6204
rect 3402 6170 3436 6204
rect 3474 6170 3508 6204
rect 3546 6170 3580 6204
rect 3618 6170 3652 6204
rect 3690 6170 3724 6204
rect 3762 6170 3796 6204
rect 3834 6170 3868 6204
rect 3906 6170 3940 6204
rect 3978 6170 4012 6204
rect 4050 6170 4084 6204
rect 4122 6170 4156 6204
rect 4194 6170 4228 6204
rect 4266 6170 4300 6204
rect 4338 6170 4372 6204
rect 4410 6170 4444 6204
rect 4482 6170 4516 6204
rect 4554 6170 4588 6204
rect 4626 6170 4660 6204
rect 4698 6170 4732 6204
rect 4770 6170 4804 6204
rect 4842 6170 4876 6204
rect 4914 6170 4948 6204
rect 4986 6170 5020 6204
rect 5058 6170 5092 6204
rect 5130 6170 5164 6204
rect 5202 6170 5236 6204
rect 5274 6170 5308 6204
rect 5346 6170 5380 6204
rect 5418 6170 5452 6204
rect 5490 6170 5524 6204
rect 5562 6170 5596 6204
rect 5634 6170 5668 6204
rect 5706 6170 5740 6204
rect 5778 6170 5812 6204
rect 5850 6170 5884 6204
rect 5922 6170 5956 6204
rect 5994 6170 6028 6204
rect 16433 6173 16467 6207
rect 16505 6173 16539 6207
rect 16577 6173 16611 6207
rect 16649 6173 16683 6207
rect 16721 6173 16755 6207
rect 16793 6173 16827 6207
rect 16865 6173 16899 6207
rect 16937 6173 16971 6207
rect 17009 6173 17043 6207
rect 17081 6173 17115 6207
rect 17153 6173 17187 6207
rect 17225 6173 17259 6207
rect 17297 6173 17331 6207
rect 17369 6173 17403 6207
rect 17441 6173 17475 6207
rect 17513 6173 17547 6207
rect 17585 6173 17619 6207
rect 17657 6173 17691 6207
rect 17729 6173 17763 6207
rect 17801 6173 17835 6207
rect 17873 6173 17907 6207
rect 17945 6173 17979 6207
rect 18017 6173 18051 6207
rect 18089 6173 18123 6207
rect 18161 6173 18195 6207
rect 18233 6173 18267 6207
rect 18305 6173 18339 6207
rect 18377 6173 18411 6207
rect 18449 6173 18483 6207
rect 18521 6173 18555 6207
rect 18593 6173 18627 6207
rect 18665 6173 18699 6207
rect 18737 6173 18771 6207
rect 18809 6173 18843 6207
rect 18881 6173 18915 6207
rect 18953 6173 18987 6207
rect 19025 6173 19059 6207
rect 19097 6173 19131 6207
rect 19169 6173 19203 6207
rect 19241 6173 19275 6207
rect 19313 6173 19347 6207
rect 19385 6173 19419 6207
rect 19457 6173 19491 6207
rect 19529 6173 19563 6207
rect 19601 6173 19635 6207
rect 19673 6173 19707 6207
rect 19745 6173 19779 6207
rect 19817 6173 19851 6207
rect 19889 6173 19923 6207
rect 19961 6173 19995 6207
rect 20033 6173 20067 6207
rect 20105 6173 20139 6207
rect 20177 6173 20211 6207
rect 20249 6173 20283 6207
rect 20321 6173 20355 6207
rect 20393 6173 20427 6207
rect 20465 6173 20499 6207
rect 20537 6173 20571 6207
rect 20609 6173 20643 6207
rect 20681 6173 20715 6207
rect 20753 6173 20787 6207
rect 20825 6173 20859 6207
rect 20897 6173 20931 6207
rect 20969 6173 21003 6207
rect 21041 6173 21075 6207
rect 21113 6173 21147 6207
rect 21185 6173 21219 6207
rect 21257 6173 21291 6207
rect 21329 6173 21363 6207
rect 21401 6173 21435 6207
rect 21473 6173 21507 6207
rect 21545 6173 21579 6207
rect 21617 6173 21651 6207
rect 21689 6173 21723 6207
rect 21761 6173 21795 6207
rect 21833 6173 21867 6207
rect 21905 6173 21939 6207
rect 21977 6173 22011 6207
rect 22049 6173 22083 6207
rect 22121 6173 22155 6207
rect 10568 1227 12258 2269
rect 10086 -7031 11848 -4837
rect 902 -7359 936 -7325
rect 974 -7359 1008 -7325
rect 1046 -7359 1080 -7325
rect 1118 -7359 1152 -7325
rect 1190 -7359 1224 -7325
rect 1262 -7359 1296 -7325
rect 1334 -7359 1368 -7325
rect 1406 -7359 1440 -7325
rect 1478 -7359 1512 -7325
rect 1550 -7359 1584 -7325
rect 1622 -7359 1656 -7325
rect 1694 -7359 1728 -7325
rect 1766 -7359 1800 -7325
rect 1838 -7359 1872 -7325
rect 1910 -7359 1944 -7325
rect 1982 -7359 2016 -7325
rect 2054 -7359 2088 -7325
rect 2126 -7359 2160 -7325
rect 2198 -7359 2232 -7325
rect 2270 -7359 2304 -7325
rect 2342 -7359 2376 -7325
rect 2414 -7359 2448 -7325
rect 2486 -7359 2520 -7325
rect 2558 -7359 2592 -7325
rect 2630 -7359 2664 -7325
rect 2702 -7359 2736 -7325
rect 2774 -7359 2808 -7325
rect 2846 -7359 2880 -7325
rect 2918 -7359 2952 -7325
rect 2990 -7359 3024 -7325
rect 3062 -7359 3096 -7325
rect 3134 -7359 3168 -7325
rect 3206 -7359 3240 -7325
rect 3278 -7359 3312 -7325
rect 3350 -7359 3384 -7325
rect 3422 -7359 3456 -7325
rect 3494 -7359 3528 -7325
rect 3566 -7359 3600 -7325
rect 3638 -7359 3672 -7325
rect 3710 -7359 3744 -7325
rect 3782 -7359 3816 -7325
rect 3854 -7359 3888 -7325
rect 3926 -7359 3960 -7325
rect 3998 -7359 4032 -7325
rect 4070 -7359 4104 -7325
rect 4142 -7359 4176 -7325
rect 4214 -7359 4248 -7325
rect 4286 -7359 4320 -7325
rect 4358 -7359 4392 -7325
rect 4430 -7359 4464 -7325
rect 4502 -7359 4536 -7325
rect 4574 -7359 4608 -7325
rect 4646 -7359 4680 -7325
rect 4718 -7359 4752 -7325
rect 4790 -7359 4824 -7325
rect 4862 -7359 4896 -7325
rect 4934 -7359 4968 -7325
rect 5006 -7359 5040 -7325
rect 5078 -7359 5112 -7325
rect 5150 -7359 5184 -7325
rect 5222 -7359 5256 -7325
rect 5294 -7359 5328 -7325
rect 5366 -7359 5400 -7325
rect 5438 -7359 5472 -7325
rect 5510 -7359 5544 -7325
rect 5582 -7359 5616 -7325
rect 5654 -7359 5688 -7325
rect 5726 -7359 5760 -7325
rect 5798 -7359 5832 -7325
rect 5870 -7359 5904 -7325
rect 5942 -7359 5976 -7325
rect 16468 -7342 16502 -7308
rect 16540 -7342 16574 -7308
rect 16612 -7342 16646 -7308
rect 16684 -7342 16718 -7308
rect 16756 -7342 16790 -7308
rect 16828 -7342 16862 -7308
rect 16900 -7342 16934 -7308
rect 16972 -7342 17006 -7308
rect 17044 -7342 17078 -7308
rect 17116 -7342 17150 -7308
rect 17188 -7342 17222 -7308
rect 17260 -7342 17294 -7308
rect 17332 -7342 17366 -7308
rect 17404 -7342 17438 -7308
rect 17476 -7342 17510 -7308
rect 17548 -7342 17582 -7308
rect 17620 -7342 17654 -7308
rect 17692 -7342 17726 -7308
rect 17764 -7342 17798 -7308
rect 17836 -7342 17870 -7308
rect 17908 -7342 17942 -7308
rect 17980 -7342 18014 -7308
rect 18052 -7342 18086 -7308
rect 18124 -7342 18158 -7308
rect 18196 -7342 18230 -7308
rect 18268 -7342 18302 -7308
rect 18340 -7342 18374 -7308
rect 18412 -7342 18446 -7308
rect 18484 -7342 18518 -7308
rect 18556 -7342 18590 -7308
rect 18628 -7342 18662 -7308
rect 18700 -7342 18734 -7308
rect 18772 -7342 18806 -7308
rect 18844 -7342 18878 -7308
rect 18916 -7342 18950 -7308
rect 18988 -7342 19022 -7308
rect 19060 -7342 19094 -7308
rect 19132 -7342 19166 -7308
rect 19204 -7342 19238 -7308
rect 19276 -7342 19310 -7308
rect 19348 -7342 19382 -7308
rect 19420 -7342 19454 -7308
rect 19492 -7342 19526 -7308
rect 19564 -7342 19598 -7308
rect 19636 -7342 19670 -7308
rect 19708 -7342 19742 -7308
rect 19780 -7342 19814 -7308
rect 19852 -7342 19886 -7308
rect 19924 -7342 19958 -7308
rect 19996 -7342 20030 -7308
rect 20068 -7342 20102 -7308
rect 20140 -7342 20174 -7308
rect 20212 -7342 20246 -7308
rect 20284 -7342 20318 -7308
rect 20356 -7342 20390 -7308
rect 20428 -7342 20462 -7308
rect 20500 -7342 20534 -7308
rect 20572 -7342 20606 -7308
rect 20644 -7342 20678 -7308
rect 20716 -7342 20750 -7308
rect 20788 -7342 20822 -7308
rect 20860 -7342 20894 -7308
rect 20932 -7342 20966 -7308
rect 21004 -7342 21038 -7308
rect 21076 -7342 21110 -7308
rect 21148 -7342 21182 -7308
rect 21220 -7342 21254 -7308
rect 21292 -7342 21326 -7308
rect 21364 -7342 21398 -7308
rect 21436 -7342 21470 -7308
rect 21508 -7342 21542 -7308
rect 21580 -7342 21614 -7308
rect 21652 -7342 21686 -7308
rect 21724 -7342 21758 -7308
rect 21796 -7342 21830 -7308
rect 21868 -7342 21902 -7308
rect 1087 -8910 5729 -8588
rect 16582 -8988 21800 -8522
<< metal1 >>
rect 140 7181 6055 7301
rect 140 6715 285 7181
rect 5863 6715 6055 7181
rect 140 6204 6055 6715
rect 140 6170 162 6204
rect 196 6170 234 6204
rect 268 6170 306 6204
rect 340 6170 378 6204
rect 412 6170 450 6204
rect 484 6170 522 6204
rect 556 6170 594 6204
rect 628 6170 666 6204
rect 700 6170 738 6204
rect 772 6170 810 6204
rect 844 6170 882 6204
rect 916 6170 954 6204
rect 988 6170 1026 6204
rect 1060 6170 1098 6204
rect 1132 6170 1170 6204
rect 1204 6170 1242 6204
rect 1276 6170 1314 6204
rect 1348 6170 1386 6204
rect 1420 6170 1458 6204
rect 1492 6170 1530 6204
rect 1564 6170 1602 6204
rect 1636 6170 1674 6204
rect 1708 6170 1746 6204
rect 1780 6170 1818 6204
rect 1852 6170 1890 6204
rect 1924 6170 1962 6204
rect 1996 6170 2034 6204
rect 2068 6170 2106 6204
rect 2140 6170 2178 6204
rect 2212 6170 2250 6204
rect 2284 6170 2322 6204
rect 2356 6170 2394 6204
rect 2428 6170 2466 6204
rect 2500 6170 2538 6204
rect 2572 6170 2610 6204
rect 2644 6170 2682 6204
rect 2716 6170 2754 6204
rect 2788 6170 2826 6204
rect 2860 6170 2898 6204
rect 2932 6170 2970 6204
rect 3004 6170 3042 6204
rect 3076 6170 3114 6204
rect 3148 6170 3186 6204
rect 3220 6170 3258 6204
rect 3292 6170 3330 6204
rect 3364 6170 3402 6204
rect 3436 6170 3474 6204
rect 3508 6170 3546 6204
rect 3580 6170 3618 6204
rect 3652 6170 3690 6204
rect 3724 6170 3762 6204
rect 3796 6170 3834 6204
rect 3868 6170 3906 6204
rect 3940 6170 3978 6204
rect 4012 6170 4050 6204
rect 4084 6170 4122 6204
rect 4156 6170 4194 6204
rect 4228 6170 4266 6204
rect 4300 6170 4338 6204
rect 4372 6170 4410 6204
rect 4444 6170 4482 6204
rect 4516 6170 4554 6204
rect 4588 6170 4626 6204
rect 4660 6170 4698 6204
rect 4732 6170 4770 6204
rect 4804 6170 4842 6204
rect 4876 6170 4914 6204
rect 4948 6170 4986 6204
rect 5020 6170 5058 6204
rect 5092 6170 5130 6204
rect 5164 6170 5202 6204
rect 5236 6170 5274 6204
rect 5308 6170 5346 6204
rect 5380 6170 5418 6204
rect 5452 6170 5490 6204
rect 5524 6170 5562 6204
rect 5596 6170 5634 6204
rect 5668 6170 5706 6204
rect 5740 6170 5778 6204
rect 5812 6170 5850 6204
rect 5884 6170 5922 6204
rect 5956 6170 5994 6204
rect 6028 6170 6055 6204
rect 140 6136 6055 6170
rect 266 2002 5862 5338
rect -8163 8 5862 2002
rect 10064 2269 12587 10493
rect 16402 7155 22219 7601
rect 16402 6761 16853 7155
rect 21927 6761 22219 7155
rect 16402 6207 22219 6761
rect 16402 6173 16433 6207
rect 16467 6173 16505 6207
rect 16539 6173 16577 6207
rect 16611 6173 16649 6207
rect 16683 6173 16721 6207
rect 16755 6173 16793 6207
rect 16827 6173 16865 6207
rect 16899 6173 16937 6207
rect 16971 6173 17009 6207
rect 17043 6173 17081 6207
rect 17115 6173 17153 6207
rect 17187 6173 17225 6207
rect 17259 6173 17297 6207
rect 17331 6173 17369 6207
rect 17403 6173 17441 6207
rect 17475 6173 17513 6207
rect 17547 6173 17585 6207
rect 17619 6173 17657 6207
rect 17691 6173 17729 6207
rect 17763 6173 17801 6207
rect 17835 6173 17873 6207
rect 17907 6173 17945 6207
rect 17979 6173 18017 6207
rect 18051 6173 18089 6207
rect 18123 6173 18161 6207
rect 18195 6173 18233 6207
rect 18267 6173 18305 6207
rect 18339 6173 18377 6207
rect 18411 6173 18449 6207
rect 18483 6173 18521 6207
rect 18555 6173 18593 6207
rect 18627 6173 18665 6207
rect 18699 6173 18737 6207
rect 18771 6173 18809 6207
rect 18843 6173 18881 6207
rect 18915 6173 18953 6207
rect 18987 6173 19025 6207
rect 19059 6173 19097 6207
rect 19131 6173 19169 6207
rect 19203 6173 19241 6207
rect 19275 6173 19313 6207
rect 19347 6173 19385 6207
rect 19419 6173 19457 6207
rect 19491 6173 19529 6207
rect 19563 6173 19601 6207
rect 19635 6173 19673 6207
rect 19707 6173 19745 6207
rect 19779 6173 19817 6207
rect 19851 6173 19889 6207
rect 19923 6173 19961 6207
rect 19995 6173 20033 6207
rect 20067 6173 20105 6207
rect 20139 6173 20177 6207
rect 20211 6173 20249 6207
rect 20283 6173 20321 6207
rect 20355 6173 20393 6207
rect 20427 6173 20465 6207
rect 20499 6173 20537 6207
rect 20571 6173 20609 6207
rect 20643 6173 20681 6207
rect 20715 6173 20753 6207
rect 20787 6173 20825 6207
rect 20859 6173 20897 6207
rect 20931 6173 20969 6207
rect 21003 6173 21041 6207
rect 21075 6173 21113 6207
rect 21147 6173 21185 6207
rect 21219 6173 21257 6207
rect 21291 6173 21329 6207
rect 21363 6173 21401 6207
rect 21435 6173 21473 6207
rect 21507 6173 21545 6207
rect 21579 6173 21617 6207
rect 21651 6173 21689 6207
rect 21723 6173 21761 6207
rect 21795 6173 21833 6207
rect 21867 6173 21905 6207
rect 21939 6173 21977 6207
rect 22011 6173 22049 6207
rect 22083 6173 22121 6207
rect 22155 6173 22219 6207
rect 16402 6145 22219 6173
rect 10064 1227 10568 2269
rect 12258 1227 12587 2269
rect 10064 831 12587 1227
rect 16266 2404 21862 5338
rect -8163 -1263 8508 8
rect 16266 -167 31050 2404
rect 14557 -866 31050 -167
rect 14563 -940 31050 -866
rect -8163 -2081 5862 -1263
rect 266 -6677 5862 -2081
rect 16266 -2451 31050 -940
rect 9571 -4837 12402 -4461
rect 9571 -7031 10086 -4837
rect 11848 -7031 12402 -4837
rect 16266 -6677 21862 -2451
rect 830 -7325 6035 -7286
rect 830 -7359 902 -7325
rect 936 -7359 974 -7325
rect 1008 -7359 1046 -7325
rect 1080 -7359 1118 -7325
rect 1152 -7359 1190 -7325
rect 1224 -7359 1262 -7325
rect 1296 -7359 1334 -7325
rect 1368 -7359 1406 -7325
rect 1440 -7359 1478 -7325
rect 1512 -7359 1550 -7325
rect 1584 -7359 1622 -7325
rect 1656 -7359 1694 -7325
rect 1728 -7359 1766 -7325
rect 1800 -7359 1838 -7325
rect 1872 -7359 1910 -7325
rect 1944 -7359 1982 -7325
rect 2016 -7359 2054 -7325
rect 2088 -7359 2126 -7325
rect 2160 -7359 2198 -7325
rect 2232 -7359 2270 -7325
rect 2304 -7359 2342 -7325
rect 2376 -7359 2414 -7325
rect 2448 -7359 2486 -7325
rect 2520 -7359 2558 -7325
rect 2592 -7359 2630 -7325
rect 2664 -7359 2702 -7325
rect 2736 -7359 2774 -7325
rect 2808 -7359 2846 -7325
rect 2880 -7359 2918 -7325
rect 2952 -7359 2990 -7325
rect 3024 -7359 3062 -7325
rect 3096 -7359 3134 -7325
rect 3168 -7359 3206 -7325
rect 3240 -7359 3278 -7325
rect 3312 -7359 3350 -7325
rect 3384 -7359 3422 -7325
rect 3456 -7359 3494 -7325
rect 3528 -7359 3566 -7325
rect 3600 -7359 3638 -7325
rect 3672 -7359 3710 -7325
rect 3744 -7359 3782 -7325
rect 3816 -7359 3854 -7325
rect 3888 -7359 3926 -7325
rect 3960 -7359 3998 -7325
rect 4032 -7359 4070 -7325
rect 4104 -7359 4142 -7325
rect 4176 -7359 4214 -7325
rect 4248 -7359 4286 -7325
rect 4320 -7359 4358 -7325
rect 4392 -7359 4430 -7325
rect 4464 -7359 4502 -7325
rect 4536 -7359 4574 -7325
rect 4608 -7359 4646 -7325
rect 4680 -7359 4718 -7325
rect 4752 -7359 4790 -7325
rect 4824 -7359 4862 -7325
rect 4896 -7359 4934 -7325
rect 4968 -7359 5006 -7325
rect 5040 -7359 5078 -7325
rect 5112 -7359 5150 -7325
rect 5184 -7359 5222 -7325
rect 5256 -7359 5294 -7325
rect 5328 -7359 5366 -7325
rect 5400 -7359 5438 -7325
rect 5472 -7359 5510 -7325
rect 5544 -7359 5582 -7325
rect 5616 -7359 5654 -7325
rect 5688 -7359 5726 -7325
rect 5760 -7359 5798 -7325
rect 5832 -7359 5870 -7325
rect 5904 -7359 5942 -7325
rect 5976 -7359 6035 -7325
rect 830 -8588 6035 -7359
rect 830 -8910 1087 -8588
rect 5729 -8910 6035 -8588
rect 830 -9170 6035 -8910
rect 9571 -12584 12402 -7031
rect 16409 -7308 21985 -7286
rect 16409 -7342 16468 -7308
rect 16502 -7342 16540 -7308
rect 16574 -7342 16612 -7308
rect 16646 -7342 16684 -7308
rect 16718 -7342 16756 -7308
rect 16790 -7342 16828 -7308
rect 16862 -7342 16900 -7308
rect 16934 -7342 16972 -7308
rect 17006 -7342 17044 -7308
rect 17078 -7342 17116 -7308
rect 17150 -7342 17188 -7308
rect 17222 -7342 17260 -7308
rect 17294 -7342 17332 -7308
rect 17366 -7342 17404 -7308
rect 17438 -7342 17476 -7308
rect 17510 -7342 17548 -7308
rect 17582 -7342 17620 -7308
rect 17654 -7342 17692 -7308
rect 17726 -7342 17764 -7308
rect 17798 -7342 17836 -7308
rect 17870 -7342 17908 -7308
rect 17942 -7342 17980 -7308
rect 18014 -7342 18052 -7308
rect 18086 -7342 18124 -7308
rect 18158 -7342 18196 -7308
rect 18230 -7342 18268 -7308
rect 18302 -7342 18340 -7308
rect 18374 -7342 18412 -7308
rect 18446 -7342 18484 -7308
rect 18518 -7342 18556 -7308
rect 18590 -7342 18628 -7308
rect 18662 -7342 18700 -7308
rect 18734 -7342 18772 -7308
rect 18806 -7342 18844 -7308
rect 18878 -7342 18916 -7308
rect 18950 -7342 18988 -7308
rect 19022 -7342 19060 -7308
rect 19094 -7342 19132 -7308
rect 19166 -7342 19204 -7308
rect 19238 -7342 19276 -7308
rect 19310 -7342 19348 -7308
rect 19382 -7342 19420 -7308
rect 19454 -7342 19492 -7308
rect 19526 -7342 19564 -7308
rect 19598 -7342 19636 -7308
rect 19670 -7342 19708 -7308
rect 19742 -7342 19780 -7308
rect 19814 -7342 19852 -7308
rect 19886 -7342 19924 -7308
rect 19958 -7342 19996 -7308
rect 20030 -7342 20068 -7308
rect 20102 -7342 20140 -7308
rect 20174 -7342 20212 -7308
rect 20246 -7342 20284 -7308
rect 20318 -7342 20356 -7308
rect 20390 -7342 20428 -7308
rect 20462 -7342 20500 -7308
rect 20534 -7342 20572 -7308
rect 20606 -7342 20644 -7308
rect 20678 -7342 20716 -7308
rect 20750 -7342 20788 -7308
rect 20822 -7342 20860 -7308
rect 20894 -7342 20932 -7308
rect 20966 -7342 21004 -7308
rect 21038 -7342 21076 -7308
rect 21110 -7342 21148 -7308
rect 21182 -7342 21220 -7308
rect 21254 -7342 21292 -7308
rect 21326 -7342 21364 -7308
rect 21398 -7342 21436 -7308
rect 21470 -7342 21508 -7308
rect 21542 -7342 21580 -7308
rect 21614 -7342 21652 -7308
rect 21686 -7342 21724 -7308
rect 21758 -7342 21796 -7308
rect 21830 -7342 21868 -7308
rect 21902 -7342 21985 -7308
rect 16409 -8522 21985 -7342
rect 16409 -8988 16582 -8522
rect 21800 -8988 21985 -8522
rect 16409 -9062 21985 -8988
use sky130_fd_pr__diode_pd2nw_05v5_4V93LZ  sky130_fd_pr__diode_pd2nw_05v5_4V93LZ_0
timestamp 1667543118
transform 1 0 19085 0 1 3085
box -3266 -3266 3266 3266
use sky130_fd_pr__diode_pd2nw_05v5_4V93LZ  sky130_fd_pr__diode_pd2nw_05v5_4V93LZ_1
timestamp 1667543118
transform 1 0 19086 0 1 -4236
box -3266 -3266 3266 3266
use sky130_fd_pr__diode_pd2nw_05v5_4V93LZ  sky130_fd_pr__diode_pd2nw_05v5_4V93LZ_2
timestamp 1667543118
transform 1 0 3086 0 1 -4236
box -3266 -3266 3266 3266
use sky130_fd_pr__diode_pd2nw_05v5_4V93LZ  sky130_fd_pr__diode_pd2nw_05v5_4V93LZ_3
timestamp 1667543118
transform 1 0 3085 0 1 3085
box -3266 -3266 3266 3266
use sky130_fd_pr__res_xhigh_po_5p73_BN6JD5  sky130_fd_pr__res_xhigh_po_5p73_BN6JD5_0
timestamp 1667543118
transform 0 1 11426 -1 0 -623
box -729 -3588 729 3588
<< end >>
