magic
tech sky130B
magscale 1 2
timestamp 1667544806
<< nwell >>
rect -6932 15844 -5270 17704
rect -3192 15796 -154 18390
rect 22964 17450 28112 19044
rect 24480 16850 28112 17450
rect 16862 15064 18378 15074
rect 12782 15058 18378 15064
rect 12782 11470 19842 15058
rect 38660 16594 40322 18454
rect 42400 16546 45438 19140
rect 14742 11464 19842 11470
rect 14742 7950 19840 11464
rect 17266 7924 19840 7950
rect 22912 13562 24506 13568
rect 22912 12052 26066 13562
rect 24472 8872 26066 12052
<< pwell >>
rect 22978 16776 24414 17384
rect 22978 16690 27710 16776
rect 22978 15888 24520 16690
rect 23084 15725 24520 15888
rect -7912 15355 -4401 15541
rect -7912 12302 -7727 15355
rect -7497 12809 -4807 14861
rect -4571 12302 -4401 15355
rect -7912 12108 -4401 12302
rect -4036 14975 -3654 15061
rect -4036 12371 -3950 14975
rect -3740 12371 -3654 14975
rect -4036 12285 -3654 12371
rect -9145 11464 -3249 11634
rect 23084 14691 23237 15725
rect 24271 15208 24520 15725
rect 27624 15208 27710 16690
rect 37680 16105 41191 16291
rect 24271 15122 27710 15208
rect 28808 15332 29826 15418
rect 24271 14691 24424 15122
rect -9145 11190 -8979 11464
rect -3428 11190 -3249 11464
rect 20356 14540 21692 14626
rect -9145 10138 -3249 11190
rect -9145 8466 -8979 10138
rect -7818 8773 -4662 9825
rect -3428 8466 -3249 10138
rect -9145 8300 -3249 8466
rect 12756 11207 14096 11360
rect 12756 10173 12909 11207
rect 13943 10173 14096 11207
rect 12756 9717 14096 10173
rect 12756 8683 12909 9717
rect 13943 8683 14096 9717
rect 12756 8530 14096 8683
rect 12756 8460 14086 8530
rect 12746 8307 14086 8460
rect -8018 7780 -3372 7908
rect -8018 7564 -7884 7780
rect -3506 7564 -3372 7780
rect -8018 5512 -3372 7564
rect -8018 5326 -7884 5512
rect -3506 5326 -3372 5512
rect -8018 5200 -3372 5326
rect 12746 7273 12899 8307
rect 13933 7273 14086 8307
rect 12746 6957 14086 7273
rect 16054 7180 17072 7266
rect 12746 5923 12899 6957
rect 13933 5923 14086 6957
rect 12746 5607 14086 5923
rect 12746 4573 12899 5607
rect 13933 4573 14086 5607
rect 12746 4420 14086 4573
rect 14396 6987 15736 7140
rect 14396 5953 14549 6987
rect 15583 5953 15736 6987
rect 14396 5627 15736 5953
rect 14396 4593 14549 5627
rect 15583 4593 15736 5627
rect 14396 4440 15736 4593
rect 16054 4576 16140 7180
rect 16986 4576 17072 7180
rect 16054 4490 17072 4576
rect 17262 4300 20148 7796
rect 20356 4650 20442 14540
rect 21606 4650 21692 14540
rect 23084 14538 24424 14691
rect 28808 13688 28894 15332
rect 29740 13688 29826 15332
rect 22882 10552 24378 11988
rect 26372 13484 27390 13500
rect 28808 13484 29826 13688
rect 26372 13414 29834 13484
rect 26372 8052 26458 13414
rect 20356 4564 21692 4650
rect 23362 3442 26458 8052
rect 26372 3010 26458 3442
rect 27304 13398 29834 13414
rect 27304 6394 27630 13398
rect 29748 6394 29834 13398
rect 37680 13052 37865 16105
rect 38095 13559 40785 15611
rect 41021 13052 41191 16105
rect 37680 12858 41191 13052
rect 41556 15725 41938 15811
rect 41556 13121 41642 15725
rect 41852 13121 41938 15725
rect 41556 13035 41938 13121
rect 36447 12214 42343 12384
rect 36447 11940 36613 12214
rect 42164 11940 42343 12214
rect 36447 10888 42343 11940
rect 36447 9216 36613 10888
rect 37774 9523 40930 10575
rect 42164 9216 42343 10888
rect 36447 9050 42343 9216
rect 27304 6308 29834 6394
rect 37574 8530 42220 8658
rect 37574 8314 37708 8530
rect 42086 8314 42220 8530
rect 27304 3010 27390 6308
rect 37574 6262 42220 8314
rect 37574 6076 37708 6262
rect 42086 6076 42220 6262
rect 37574 5950 42220 6076
rect 26372 2924 27390 3010
<< nbase >>
rect 23237 14691 24271 15725
rect 12909 10173 13943 11207
rect 12909 8683 13943 9717
rect 12899 7273 13933 8307
rect 12899 5923 13933 6957
rect 12899 4573 13933 5607
rect 14549 5953 15583 6987
rect 14549 4593 15583 5627
<< mvnmos >>
rect 23196 16136 24196 17136
rect -7413 12835 -7213 14835
rect -7155 12835 -6955 14835
rect -6897 12835 -6697 14835
rect -6639 12835 -6439 14835
rect -6381 12835 -6181 14835
rect -6123 12835 -5923 14835
rect -5865 12835 -5665 14835
rect -5607 12835 -5407 14835
rect -5349 12835 -5149 14835
rect -5091 12835 -4891 14835
rect -8769 10164 -8569 11164
rect -8511 10164 -8311 11164
rect -8253 10164 -8053 11164
rect -7995 10164 -7795 11164
rect -7737 10164 -7537 11164
rect -7479 10164 -7279 11164
rect -7221 10164 -7021 11164
rect -6963 10164 -6763 11164
rect -6705 10164 -6505 11164
rect -6447 10164 -6247 11164
rect -6189 10164 -5989 11164
rect -5931 10164 -5731 11164
rect -5673 10164 -5473 11164
rect -5415 10164 -5215 11164
rect -5157 10164 -4957 11164
rect -4899 10164 -4699 11164
rect -4641 10164 -4441 11164
rect -4383 10164 -4183 11164
rect -4125 10164 -3925 11164
rect -3867 10164 -3667 11164
rect -7734 8799 -7534 9799
rect -7268 8799 -7068 9799
rect -7010 8799 -6810 9799
rect -6752 8799 -6552 9799
rect -6494 8799 -6294 9799
rect -6236 8799 -6036 9799
rect -5978 8799 -5778 9799
rect -5720 8799 -5520 9799
rect -5462 8799 -5262 9799
rect -5204 8799 -5004 9799
rect -4946 8799 -4746 9799
rect -7734 5538 -7534 7538
rect -7476 5538 -7276 7538
rect -7218 5538 -7018 7538
rect -6960 5538 -6760 7538
rect -6702 5538 -6502 7538
rect -6444 5538 -6244 7538
rect -6186 5538 -5986 7538
rect -5928 5538 -5728 7538
rect -5670 5538 -5470 7538
rect -5412 5538 -5212 7538
rect -5154 5538 -4954 7538
rect -4896 5538 -4696 7538
rect -4638 5538 -4438 7538
rect -4380 5538 -4180 7538
rect -4122 5538 -3922 7538
rect -3864 5538 -3664 7538
rect 17480 4548 18480 7548
rect 18930 4548 19930 7548
rect 38179 13585 38379 15585
rect 38437 13585 38637 15585
rect 38695 13585 38895 15585
rect 38953 13585 39153 15585
rect 39211 13585 39411 15585
rect 39469 13585 39669 15585
rect 39727 13585 39927 15585
rect 39985 13585 40185 15585
rect 40243 13585 40443 15585
rect 40501 13585 40701 15585
rect 23130 10770 24130 11770
rect 23610 6834 24610 7834
rect 23610 5776 24610 6776
rect 23610 4718 24610 5718
rect 23610 3660 24610 4660
rect 25110 6834 26110 7834
rect 25110 5776 26110 6776
rect 25110 4718 26110 5718
rect 25110 3660 26110 4660
rect 36823 10914 37023 11914
rect 37081 10914 37281 11914
rect 37339 10914 37539 11914
rect 37597 10914 37797 11914
rect 37855 10914 38055 11914
rect 38113 10914 38313 11914
rect 38371 10914 38571 11914
rect 38629 10914 38829 11914
rect 38887 10914 39087 11914
rect 39145 10914 39345 11914
rect 39403 10914 39603 11914
rect 39661 10914 39861 11914
rect 39919 10914 40119 11914
rect 40177 10914 40377 11914
rect 40435 10914 40635 11914
rect 40693 10914 40893 11914
rect 40951 10914 41151 11914
rect 41209 10914 41409 11914
rect 41467 10914 41667 11914
rect 41725 10914 41925 11914
rect 37858 9549 38058 10549
rect 38324 9549 38524 10549
rect 38582 9549 38782 10549
rect 38840 9549 39040 10549
rect 39098 9549 39298 10549
rect 39356 9549 39556 10549
rect 39614 9549 39814 10549
rect 39872 9549 40072 10549
rect 40130 9549 40330 10549
rect 40388 9549 40588 10549
rect 40646 9549 40846 10549
rect 37858 6288 38058 8288
rect 38116 6288 38316 8288
rect 38374 6288 38574 8288
rect 38632 6288 38832 8288
rect 38890 6288 39090 8288
rect 39148 6288 39348 8288
rect 39406 6288 39606 8288
rect 39664 6288 39864 8288
rect 39922 6288 40122 8288
rect 40180 6288 40380 8288
rect 40438 6288 40638 8288
rect 40696 6288 40896 8288
rect 40954 6288 41154 8288
rect 41212 6288 41412 8288
rect 41470 6288 41670 8288
rect 41728 6288 41928 8288
<< mvpmos >>
rect -6402 16224 -6202 17224
rect -6144 16224 -5944 17224
rect -2934 16093 -2734 18093
rect -2676 16093 -2476 18093
rect -2418 16093 -2218 18093
rect -2160 16093 -1960 18093
rect -1902 16093 -1702 18093
rect -1644 16093 -1444 18093
rect -1386 16093 -1186 18093
rect -1128 16093 -928 18093
rect -870 16093 -670 18093
rect -612 16093 -412 18093
rect 23222 17747 24222 18747
rect 24738 17147 25738 18747
rect 25796 17147 26796 18747
rect 26854 17147 27854 18747
rect 39190 16974 39390 17974
rect 39448 16974 39648 17974
rect 42658 16843 42858 18843
rect 42916 16843 43116 18843
rect 43174 16843 43374 18843
rect 43432 16843 43632 18843
rect 43690 16843 43890 18843
rect 43948 16843 44148 18843
rect 44206 16843 44406 18843
rect 44464 16843 44664 18843
rect 44722 16843 44922 18843
rect 44980 16843 45180 18843
rect 13040 11767 14040 14767
rect 14098 11767 15098 14767
rect 15610 11767 16610 14767
rect 17120 11777 18120 14777
rect 18584 11761 19584 14761
rect 15000 8247 16000 11247
rect 16058 8247 17058 11247
rect 17524 8221 18524 11221
rect 18582 8221 19582 11221
rect 23209 12310 24209 13310
rect 24769 12304 25769 13304
rect 24769 11246 25769 12246
rect 24769 10188 25769 11188
rect 24769 9130 25769 10130
<< pdiff >>
rect 23414 15496 24094 15548
rect 23414 15462 23468 15496
rect 23502 15462 23558 15496
rect 23592 15462 23648 15496
rect 23682 15462 23738 15496
rect 23772 15462 23828 15496
rect 23862 15462 23918 15496
rect 23952 15462 24008 15496
rect 24042 15462 24094 15496
rect 23414 15406 24094 15462
rect 23414 15372 23468 15406
rect 23502 15372 23558 15406
rect 23592 15372 23648 15406
rect 23682 15372 23738 15406
rect 23772 15372 23828 15406
rect 23862 15372 23918 15406
rect 23952 15372 24008 15406
rect 24042 15372 24094 15406
rect 23414 15316 24094 15372
rect 23414 15282 23468 15316
rect 23502 15282 23558 15316
rect 23592 15282 23648 15316
rect 23682 15282 23738 15316
rect 23772 15282 23828 15316
rect 23862 15282 23918 15316
rect 23952 15282 24008 15316
rect 24042 15282 24094 15316
rect 23414 15226 24094 15282
rect 23414 15192 23468 15226
rect 23502 15192 23558 15226
rect 23592 15192 23648 15226
rect 23682 15192 23738 15226
rect 23772 15192 23828 15226
rect 23862 15192 23918 15226
rect 23952 15192 24008 15226
rect 24042 15192 24094 15226
rect 23414 15136 24094 15192
rect 23414 15102 23468 15136
rect 23502 15102 23558 15136
rect 23592 15102 23648 15136
rect 23682 15102 23738 15136
rect 23772 15102 23828 15136
rect 23862 15102 23918 15136
rect 23952 15102 24008 15136
rect 24042 15102 24094 15136
rect 23414 15046 24094 15102
rect 23414 15012 23468 15046
rect 23502 15012 23558 15046
rect 23592 15012 23648 15046
rect 23682 15012 23738 15046
rect 23772 15012 23828 15046
rect 23862 15012 23918 15046
rect 23952 15012 24008 15046
rect 24042 15012 24094 15046
rect 23414 14956 24094 15012
rect 23414 14922 23468 14956
rect 23502 14922 23558 14956
rect 23592 14922 23648 14956
rect 23682 14922 23738 14956
rect 23772 14922 23828 14956
rect 23862 14922 23918 14956
rect 23952 14922 24008 14956
rect 24042 14922 24094 14956
rect 23414 14868 24094 14922
rect 13086 10978 13766 11030
rect 13086 10944 13140 10978
rect 13174 10944 13230 10978
rect 13264 10944 13320 10978
rect 13354 10944 13410 10978
rect 13444 10944 13500 10978
rect 13534 10944 13590 10978
rect 13624 10944 13680 10978
rect 13714 10944 13766 10978
rect 13086 10888 13766 10944
rect 13086 10854 13140 10888
rect 13174 10854 13230 10888
rect 13264 10854 13320 10888
rect 13354 10854 13410 10888
rect 13444 10854 13500 10888
rect 13534 10854 13590 10888
rect 13624 10854 13680 10888
rect 13714 10854 13766 10888
rect 13086 10798 13766 10854
rect 13086 10764 13140 10798
rect 13174 10764 13230 10798
rect 13264 10764 13320 10798
rect 13354 10764 13410 10798
rect 13444 10764 13500 10798
rect 13534 10764 13590 10798
rect 13624 10764 13680 10798
rect 13714 10764 13766 10798
rect 13086 10708 13766 10764
rect 13086 10674 13140 10708
rect 13174 10674 13230 10708
rect 13264 10674 13320 10708
rect 13354 10674 13410 10708
rect 13444 10674 13500 10708
rect 13534 10674 13590 10708
rect 13624 10674 13680 10708
rect 13714 10674 13766 10708
rect 13086 10618 13766 10674
rect 13086 10584 13140 10618
rect 13174 10584 13230 10618
rect 13264 10584 13320 10618
rect 13354 10584 13410 10618
rect 13444 10584 13500 10618
rect 13534 10584 13590 10618
rect 13624 10584 13680 10618
rect 13714 10584 13766 10618
rect 13086 10528 13766 10584
rect 13086 10494 13140 10528
rect 13174 10494 13230 10528
rect 13264 10494 13320 10528
rect 13354 10494 13410 10528
rect 13444 10494 13500 10528
rect 13534 10494 13590 10528
rect 13624 10494 13680 10528
rect 13714 10494 13766 10528
rect 13086 10438 13766 10494
rect 13086 10404 13140 10438
rect 13174 10404 13230 10438
rect 13264 10404 13320 10438
rect 13354 10404 13410 10438
rect 13444 10404 13500 10438
rect 13534 10404 13590 10438
rect 13624 10404 13680 10438
rect 13714 10404 13766 10438
rect 13086 10350 13766 10404
rect 13086 9488 13766 9540
rect 13086 9454 13140 9488
rect 13174 9454 13230 9488
rect 13264 9454 13320 9488
rect 13354 9454 13410 9488
rect 13444 9454 13500 9488
rect 13534 9454 13590 9488
rect 13624 9454 13680 9488
rect 13714 9454 13766 9488
rect 13086 9398 13766 9454
rect 13086 9364 13140 9398
rect 13174 9364 13230 9398
rect 13264 9364 13320 9398
rect 13354 9364 13410 9398
rect 13444 9364 13500 9398
rect 13534 9364 13590 9398
rect 13624 9364 13680 9398
rect 13714 9364 13766 9398
rect 13086 9308 13766 9364
rect 13086 9274 13140 9308
rect 13174 9274 13230 9308
rect 13264 9274 13320 9308
rect 13354 9274 13410 9308
rect 13444 9274 13500 9308
rect 13534 9274 13590 9308
rect 13624 9274 13680 9308
rect 13714 9274 13766 9308
rect 13086 9218 13766 9274
rect 13086 9184 13140 9218
rect 13174 9184 13230 9218
rect 13264 9184 13320 9218
rect 13354 9184 13410 9218
rect 13444 9184 13500 9218
rect 13534 9184 13590 9218
rect 13624 9184 13680 9218
rect 13714 9184 13766 9218
rect 13086 9128 13766 9184
rect 13086 9094 13140 9128
rect 13174 9094 13230 9128
rect 13264 9094 13320 9128
rect 13354 9094 13410 9128
rect 13444 9094 13500 9128
rect 13534 9094 13590 9128
rect 13624 9094 13680 9128
rect 13714 9094 13766 9128
rect 13086 9038 13766 9094
rect 13086 9004 13140 9038
rect 13174 9004 13230 9038
rect 13264 9004 13320 9038
rect 13354 9004 13410 9038
rect 13444 9004 13500 9038
rect 13534 9004 13590 9038
rect 13624 9004 13680 9038
rect 13714 9004 13766 9038
rect 13086 8948 13766 9004
rect 13086 8914 13140 8948
rect 13174 8914 13230 8948
rect 13264 8914 13320 8948
rect 13354 8914 13410 8948
rect 13444 8914 13500 8948
rect 13534 8914 13590 8948
rect 13624 8914 13680 8948
rect 13714 8914 13766 8948
rect 13086 8860 13766 8914
rect 13076 8078 13756 8130
rect 13076 8044 13130 8078
rect 13164 8044 13220 8078
rect 13254 8044 13310 8078
rect 13344 8044 13400 8078
rect 13434 8044 13490 8078
rect 13524 8044 13580 8078
rect 13614 8044 13670 8078
rect 13704 8044 13756 8078
rect 13076 7988 13756 8044
rect 13076 7954 13130 7988
rect 13164 7954 13220 7988
rect 13254 7954 13310 7988
rect 13344 7954 13400 7988
rect 13434 7954 13490 7988
rect 13524 7954 13580 7988
rect 13614 7954 13670 7988
rect 13704 7954 13756 7988
rect 13076 7898 13756 7954
rect 13076 7864 13130 7898
rect 13164 7864 13220 7898
rect 13254 7864 13310 7898
rect 13344 7864 13400 7898
rect 13434 7864 13490 7898
rect 13524 7864 13580 7898
rect 13614 7864 13670 7898
rect 13704 7864 13756 7898
rect 13076 7808 13756 7864
rect 13076 7774 13130 7808
rect 13164 7774 13220 7808
rect 13254 7774 13310 7808
rect 13344 7774 13400 7808
rect 13434 7774 13490 7808
rect 13524 7774 13580 7808
rect 13614 7774 13670 7808
rect 13704 7774 13756 7808
rect 13076 7718 13756 7774
rect 13076 7684 13130 7718
rect 13164 7684 13220 7718
rect 13254 7684 13310 7718
rect 13344 7684 13400 7718
rect 13434 7684 13490 7718
rect 13524 7684 13580 7718
rect 13614 7684 13670 7718
rect 13704 7684 13756 7718
rect 13076 7628 13756 7684
rect 13076 7594 13130 7628
rect 13164 7594 13220 7628
rect 13254 7594 13310 7628
rect 13344 7594 13400 7628
rect 13434 7594 13490 7628
rect 13524 7594 13580 7628
rect 13614 7594 13670 7628
rect 13704 7594 13756 7628
rect 13076 7538 13756 7594
rect 13076 7504 13130 7538
rect 13164 7504 13220 7538
rect 13254 7504 13310 7538
rect 13344 7504 13400 7538
rect 13434 7504 13490 7538
rect 13524 7504 13580 7538
rect 13614 7504 13670 7538
rect 13704 7504 13756 7538
rect 13076 7450 13756 7504
rect 13076 6728 13756 6780
rect 13076 6694 13130 6728
rect 13164 6694 13220 6728
rect 13254 6694 13310 6728
rect 13344 6694 13400 6728
rect 13434 6694 13490 6728
rect 13524 6694 13580 6728
rect 13614 6694 13670 6728
rect 13704 6694 13756 6728
rect 13076 6638 13756 6694
rect 13076 6604 13130 6638
rect 13164 6604 13220 6638
rect 13254 6604 13310 6638
rect 13344 6604 13400 6638
rect 13434 6604 13490 6638
rect 13524 6604 13580 6638
rect 13614 6604 13670 6638
rect 13704 6604 13756 6638
rect 13076 6548 13756 6604
rect 13076 6514 13130 6548
rect 13164 6514 13220 6548
rect 13254 6514 13310 6548
rect 13344 6514 13400 6548
rect 13434 6514 13490 6548
rect 13524 6514 13580 6548
rect 13614 6514 13670 6548
rect 13704 6514 13756 6548
rect 13076 6458 13756 6514
rect 13076 6424 13130 6458
rect 13164 6424 13220 6458
rect 13254 6424 13310 6458
rect 13344 6424 13400 6458
rect 13434 6424 13490 6458
rect 13524 6424 13580 6458
rect 13614 6424 13670 6458
rect 13704 6424 13756 6458
rect 13076 6368 13756 6424
rect 13076 6334 13130 6368
rect 13164 6334 13220 6368
rect 13254 6334 13310 6368
rect 13344 6334 13400 6368
rect 13434 6334 13490 6368
rect 13524 6334 13580 6368
rect 13614 6334 13670 6368
rect 13704 6334 13756 6368
rect 13076 6278 13756 6334
rect 13076 6244 13130 6278
rect 13164 6244 13220 6278
rect 13254 6244 13310 6278
rect 13344 6244 13400 6278
rect 13434 6244 13490 6278
rect 13524 6244 13580 6278
rect 13614 6244 13670 6278
rect 13704 6244 13756 6278
rect 13076 6188 13756 6244
rect 13076 6154 13130 6188
rect 13164 6154 13220 6188
rect 13254 6154 13310 6188
rect 13344 6154 13400 6188
rect 13434 6154 13490 6188
rect 13524 6154 13580 6188
rect 13614 6154 13670 6188
rect 13704 6154 13756 6188
rect 13076 6100 13756 6154
rect 14726 6758 15406 6810
rect 14726 6724 14780 6758
rect 14814 6724 14870 6758
rect 14904 6724 14960 6758
rect 14994 6724 15050 6758
rect 15084 6724 15140 6758
rect 15174 6724 15230 6758
rect 15264 6724 15320 6758
rect 15354 6724 15406 6758
rect 14726 6668 15406 6724
rect 14726 6634 14780 6668
rect 14814 6634 14870 6668
rect 14904 6634 14960 6668
rect 14994 6634 15050 6668
rect 15084 6634 15140 6668
rect 15174 6634 15230 6668
rect 15264 6634 15320 6668
rect 15354 6634 15406 6668
rect 14726 6578 15406 6634
rect 14726 6544 14780 6578
rect 14814 6544 14870 6578
rect 14904 6544 14960 6578
rect 14994 6544 15050 6578
rect 15084 6544 15140 6578
rect 15174 6544 15230 6578
rect 15264 6544 15320 6578
rect 15354 6544 15406 6578
rect 14726 6488 15406 6544
rect 14726 6454 14780 6488
rect 14814 6454 14870 6488
rect 14904 6454 14960 6488
rect 14994 6454 15050 6488
rect 15084 6454 15140 6488
rect 15174 6454 15230 6488
rect 15264 6454 15320 6488
rect 15354 6454 15406 6488
rect 14726 6398 15406 6454
rect 14726 6364 14780 6398
rect 14814 6364 14870 6398
rect 14904 6364 14960 6398
rect 14994 6364 15050 6398
rect 15084 6364 15140 6398
rect 15174 6364 15230 6398
rect 15264 6364 15320 6398
rect 15354 6364 15406 6398
rect 14726 6308 15406 6364
rect 14726 6274 14780 6308
rect 14814 6274 14870 6308
rect 14904 6274 14960 6308
rect 14994 6274 15050 6308
rect 15084 6274 15140 6308
rect 15174 6274 15230 6308
rect 15264 6274 15320 6308
rect 15354 6274 15406 6308
rect 14726 6218 15406 6274
rect 14726 6184 14780 6218
rect 14814 6184 14870 6218
rect 14904 6184 14960 6218
rect 14994 6184 15050 6218
rect 15084 6184 15140 6218
rect 15174 6184 15230 6218
rect 15264 6184 15320 6218
rect 15354 6184 15406 6218
rect 14726 6130 15406 6184
rect 13076 5378 13756 5430
rect 13076 5344 13130 5378
rect 13164 5344 13220 5378
rect 13254 5344 13310 5378
rect 13344 5344 13400 5378
rect 13434 5344 13490 5378
rect 13524 5344 13580 5378
rect 13614 5344 13670 5378
rect 13704 5344 13756 5378
rect 13076 5288 13756 5344
rect 13076 5254 13130 5288
rect 13164 5254 13220 5288
rect 13254 5254 13310 5288
rect 13344 5254 13400 5288
rect 13434 5254 13490 5288
rect 13524 5254 13580 5288
rect 13614 5254 13670 5288
rect 13704 5254 13756 5288
rect 13076 5198 13756 5254
rect 13076 5164 13130 5198
rect 13164 5164 13220 5198
rect 13254 5164 13310 5198
rect 13344 5164 13400 5198
rect 13434 5164 13490 5198
rect 13524 5164 13580 5198
rect 13614 5164 13670 5198
rect 13704 5164 13756 5198
rect 13076 5108 13756 5164
rect 13076 5074 13130 5108
rect 13164 5074 13220 5108
rect 13254 5074 13310 5108
rect 13344 5074 13400 5108
rect 13434 5074 13490 5108
rect 13524 5074 13580 5108
rect 13614 5074 13670 5108
rect 13704 5074 13756 5108
rect 13076 5018 13756 5074
rect 13076 4984 13130 5018
rect 13164 4984 13220 5018
rect 13254 4984 13310 5018
rect 13344 4984 13400 5018
rect 13434 4984 13490 5018
rect 13524 4984 13580 5018
rect 13614 4984 13670 5018
rect 13704 4984 13756 5018
rect 13076 4928 13756 4984
rect 13076 4894 13130 4928
rect 13164 4894 13220 4928
rect 13254 4894 13310 4928
rect 13344 4894 13400 4928
rect 13434 4894 13490 4928
rect 13524 4894 13580 4928
rect 13614 4894 13670 4928
rect 13704 4894 13756 4928
rect 13076 4838 13756 4894
rect 13076 4804 13130 4838
rect 13164 4804 13220 4838
rect 13254 4804 13310 4838
rect 13344 4804 13400 4838
rect 13434 4804 13490 4838
rect 13524 4804 13580 4838
rect 13614 4804 13670 4838
rect 13704 4804 13756 4838
rect 13076 4750 13756 4804
rect 14726 5398 15406 5450
rect 14726 5364 14780 5398
rect 14814 5364 14870 5398
rect 14904 5364 14960 5398
rect 14994 5364 15050 5398
rect 15084 5364 15140 5398
rect 15174 5364 15230 5398
rect 15264 5364 15320 5398
rect 15354 5364 15406 5398
rect 14726 5308 15406 5364
rect 14726 5274 14780 5308
rect 14814 5274 14870 5308
rect 14904 5274 14960 5308
rect 14994 5274 15050 5308
rect 15084 5274 15140 5308
rect 15174 5274 15230 5308
rect 15264 5274 15320 5308
rect 15354 5274 15406 5308
rect 14726 5218 15406 5274
rect 14726 5184 14780 5218
rect 14814 5184 14870 5218
rect 14904 5184 14960 5218
rect 14994 5184 15050 5218
rect 15084 5184 15140 5218
rect 15174 5184 15230 5218
rect 15264 5184 15320 5218
rect 15354 5184 15406 5218
rect 14726 5128 15406 5184
rect 14726 5094 14780 5128
rect 14814 5094 14870 5128
rect 14904 5094 14960 5128
rect 14994 5094 15050 5128
rect 15084 5094 15140 5128
rect 15174 5094 15230 5128
rect 15264 5094 15320 5128
rect 15354 5094 15406 5128
rect 14726 5038 15406 5094
rect 14726 5004 14780 5038
rect 14814 5004 14870 5038
rect 14904 5004 14960 5038
rect 14994 5004 15050 5038
rect 15084 5004 15140 5038
rect 15174 5004 15230 5038
rect 15264 5004 15320 5038
rect 15354 5004 15406 5038
rect 14726 4948 15406 5004
rect 14726 4914 14780 4948
rect 14814 4914 14870 4948
rect 14904 4914 14960 4948
rect 14994 4914 15050 4948
rect 15084 4914 15140 4948
rect 15174 4914 15230 4948
rect 15264 4914 15320 4948
rect 15354 4914 15406 4948
rect 14726 4858 15406 4914
rect 14726 4824 14780 4858
rect 14814 4824 14870 4858
rect 14904 4824 14960 4858
rect 14994 4824 15050 4858
rect 15084 4824 15140 4858
rect 15174 4824 15230 4858
rect 15264 4824 15320 4858
rect 15354 4824 15406 4858
rect 14726 4770 15406 4824
<< mvndiff >>
rect 23138 17095 23196 17136
rect 23138 17061 23150 17095
rect 23184 17061 23196 17095
rect 23138 17027 23196 17061
rect 23138 16993 23150 17027
rect 23184 16993 23196 17027
rect 23138 16959 23196 16993
rect 23138 16925 23150 16959
rect 23184 16925 23196 16959
rect 23138 16891 23196 16925
rect 23138 16857 23150 16891
rect 23184 16857 23196 16891
rect 23138 16823 23196 16857
rect 23138 16789 23150 16823
rect 23184 16789 23196 16823
rect 23138 16755 23196 16789
rect 23138 16721 23150 16755
rect 23184 16721 23196 16755
rect 23138 16687 23196 16721
rect 23138 16653 23150 16687
rect 23184 16653 23196 16687
rect 23138 16619 23196 16653
rect 23138 16585 23150 16619
rect 23184 16585 23196 16619
rect 23138 16551 23196 16585
rect 23138 16517 23150 16551
rect 23184 16517 23196 16551
rect 23138 16483 23196 16517
rect 23138 16449 23150 16483
rect 23184 16449 23196 16483
rect 23138 16415 23196 16449
rect 23138 16381 23150 16415
rect 23184 16381 23196 16415
rect 23138 16347 23196 16381
rect 23138 16313 23150 16347
rect 23184 16313 23196 16347
rect 23138 16279 23196 16313
rect 23138 16245 23150 16279
rect 23184 16245 23196 16279
rect 23138 16211 23196 16245
rect 23138 16177 23150 16211
rect 23184 16177 23196 16211
rect 23138 16136 23196 16177
rect 24196 17095 24254 17136
rect 24196 17061 24208 17095
rect 24242 17061 24254 17095
rect 24196 17027 24254 17061
rect 24196 16993 24208 17027
rect 24242 16993 24254 17027
rect 24196 16959 24254 16993
rect 24196 16925 24208 16959
rect 24242 16925 24254 16959
rect 24196 16891 24254 16925
rect 24196 16857 24208 16891
rect 24242 16857 24254 16891
rect 24196 16823 24254 16857
rect 24196 16789 24208 16823
rect 24242 16789 24254 16823
rect 24196 16755 24254 16789
rect 24196 16721 24208 16755
rect 24242 16721 24254 16755
rect 24196 16687 24254 16721
rect 24196 16653 24208 16687
rect 24242 16653 24254 16687
rect 24196 16619 24254 16653
rect 24196 16585 24208 16619
rect 24242 16585 24254 16619
rect 24196 16551 24254 16585
rect 24196 16517 24208 16551
rect 24242 16517 24254 16551
rect 24196 16483 24254 16517
rect 24196 16449 24208 16483
rect 24242 16449 24254 16483
rect 24196 16415 24254 16449
rect 24196 16381 24208 16415
rect 24242 16381 24254 16415
rect 24196 16347 24254 16381
rect 24196 16313 24208 16347
rect 24242 16313 24254 16347
rect 24196 16279 24254 16313
rect 24196 16245 24208 16279
rect 24242 16245 24254 16279
rect 24196 16211 24254 16245
rect 24196 16177 24208 16211
rect 24242 16177 24254 16211
rect 24196 16136 24254 16177
rect -7471 14804 -7413 14835
rect -7471 14770 -7459 14804
rect -7425 14770 -7413 14804
rect -7471 14736 -7413 14770
rect -7471 14702 -7459 14736
rect -7425 14702 -7413 14736
rect -7471 14668 -7413 14702
rect -7471 14634 -7459 14668
rect -7425 14634 -7413 14668
rect -7471 14600 -7413 14634
rect -7471 14566 -7459 14600
rect -7425 14566 -7413 14600
rect -7471 14532 -7413 14566
rect -7471 14498 -7459 14532
rect -7425 14498 -7413 14532
rect -7471 14464 -7413 14498
rect -7471 14430 -7459 14464
rect -7425 14430 -7413 14464
rect -7471 14396 -7413 14430
rect -7471 14362 -7459 14396
rect -7425 14362 -7413 14396
rect -7471 14328 -7413 14362
rect -7471 14294 -7459 14328
rect -7425 14294 -7413 14328
rect -7471 14260 -7413 14294
rect -7471 14226 -7459 14260
rect -7425 14226 -7413 14260
rect -7471 14192 -7413 14226
rect -7471 14158 -7459 14192
rect -7425 14158 -7413 14192
rect -7471 14124 -7413 14158
rect -7471 14090 -7459 14124
rect -7425 14090 -7413 14124
rect -7471 14056 -7413 14090
rect -7471 14022 -7459 14056
rect -7425 14022 -7413 14056
rect -7471 13988 -7413 14022
rect -7471 13954 -7459 13988
rect -7425 13954 -7413 13988
rect -7471 13920 -7413 13954
rect -7471 13886 -7459 13920
rect -7425 13886 -7413 13920
rect -7471 13852 -7413 13886
rect -7471 13818 -7459 13852
rect -7425 13818 -7413 13852
rect -7471 13784 -7413 13818
rect -7471 13750 -7459 13784
rect -7425 13750 -7413 13784
rect -7471 13716 -7413 13750
rect -7471 13682 -7459 13716
rect -7425 13682 -7413 13716
rect -7471 13648 -7413 13682
rect -7471 13614 -7459 13648
rect -7425 13614 -7413 13648
rect -7471 13580 -7413 13614
rect -7471 13546 -7459 13580
rect -7425 13546 -7413 13580
rect -7471 13512 -7413 13546
rect -7471 13478 -7459 13512
rect -7425 13478 -7413 13512
rect -7471 13444 -7413 13478
rect -7471 13410 -7459 13444
rect -7425 13410 -7413 13444
rect -7471 13376 -7413 13410
rect -7471 13342 -7459 13376
rect -7425 13342 -7413 13376
rect -7471 13308 -7413 13342
rect -7471 13274 -7459 13308
rect -7425 13274 -7413 13308
rect -7471 13240 -7413 13274
rect -7471 13206 -7459 13240
rect -7425 13206 -7413 13240
rect -7471 13172 -7413 13206
rect -7471 13138 -7459 13172
rect -7425 13138 -7413 13172
rect -7471 13104 -7413 13138
rect -7471 13070 -7459 13104
rect -7425 13070 -7413 13104
rect -7471 13036 -7413 13070
rect -7471 13002 -7459 13036
rect -7425 13002 -7413 13036
rect -7471 12968 -7413 13002
rect -7471 12934 -7459 12968
rect -7425 12934 -7413 12968
rect -7471 12900 -7413 12934
rect -7471 12866 -7459 12900
rect -7425 12866 -7413 12900
rect -7471 12835 -7413 12866
rect -7213 14804 -7155 14835
rect -7213 14770 -7201 14804
rect -7167 14770 -7155 14804
rect -7213 14736 -7155 14770
rect -7213 14702 -7201 14736
rect -7167 14702 -7155 14736
rect -7213 14668 -7155 14702
rect -7213 14634 -7201 14668
rect -7167 14634 -7155 14668
rect -7213 14600 -7155 14634
rect -7213 14566 -7201 14600
rect -7167 14566 -7155 14600
rect -7213 14532 -7155 14566
rect -7213 14498 -7201 14532
rect -7167 14498 -7155 14532
rect -7213 14464 -7155 14498
rect -7213 14430 -7201 14464
rect -7167 14430 -7155 14464
rect -7213 14396 -7155 14430
rect -7213 14362 -7201 14396
rect -7167 14362 -7155 14396
rect -7213 14328 -7155 14362
rect -7213 14294 -7201 14328
rect -7167 14294 -7155 14328
rect -7213 14260 -7155 14294
rect -7213 14226 -7201 14260
rect -7167 14226 -7155 14260
rect -7213 14192 -7155 14226
rect -7213 14158 -7201 14192
rect -7167 14158 -7155 14192
rect -7213 14124 -7155 14158
rect -7213 14090 -7201 14124
rect -7167 14090 -7155 14124
rect -7213 14056 -7155 14090
rect -7213 14022 -7201 14056
rect -7167 14022 -7155 14056
rect -7213 13988 -7155 14022
rect -7213 13954 -7201 13988
rect -7167 13954 -7155 13988
rect -7213 13920 -7155 13954
rect -7213 13886 -7201 13920
rect -7167 13886 -7155 13920
rect -7213 13852 -7155 13886
rect -7213 13818 -7201 13852
rect -7167 13818 -7155 13852
rect -7213 13784 -7155 13818
rect -7213 13750 -7201 13784
rect -7167 13750 -7155 13784
rect -7213 13716 -7155 13750
rect -7213 13682 -7201 13716
rect -7167 13682 -7155 13716
rect -7213 13648 -7155 13682
rect -7213 13614 -7201 13648
rect -7167 13614 -7155 13648
rect -7213 13580 -7155 13614
rect -7213 13546 -7201 13580
rect -7167 13546 -7155 13580
rect -7213 13512 -7155 13546
rect -7213 13478 -7201 13512
rect -7167 13478 -7155 13512
rect -7213 13444 -7155 13478
rect -7213 13410 -7201 13444
rect -7167 13410 -7155 13444
rect -7213 13376 -7155 13410
rect -7213 13342 -7201 13376
rect -7167 13342 -7155 13376
rect -7213 13308 -7155 13342
rect -7213 13274 -7201 13308
rect -7167 13274 -7155 13308
rect -7213 13240 -7155 13274
rect -7213 13206 -7201 13240
rect -7167 13206 -7155 13240
rect -7213 13172 -7155 13206
rect -7213 13138 -7201 13172
rect -7167 13138 -7155 13172
rect -7213 13104 -7155 13138
rect -7213 13070 -7201 13104
rect -7167 13070 -7155 13104
rect -7213 13036 -7155 13070
rect -7213 13002 -7201 13036
rect -7167 13002 -7155 13036
rect -7213 12968 -7155 13002
rect -7213 12934 -7201 12968
rect -7167 12934 -7155 12968
rect -7213 12900 -7155 12934
rect -7213 12866 -7201 12900
rect -7167 12866 -7155 12900
rect -7213 12835 -7155 12866
rect -6955 14804 -6897 14835
rect -6955 14770 -6943 14804
rect -6909 14770 -6897 14804
rect -6955 14736 -6897 14770
rect -6955 14702 -6943 14736
rect -6909 14702 -6897 14736
rect -6955 14668 -6897 14702
rect -6955 14634 -6943 14668
rect -6909 14634 -6897 14668
rect -6955 14600 -6897 14634
rect -6955 14566 -6943 14600
rect -6909 14566 -6897 14600
rect -6955 14532 -6897 14566
rect -6955 14498 -6943 14532
rect -6909 14498 -6897 14532
rect -6955 14464 -6897 14498
rect -6955 14430 -6943 14464
rect -6909 14430 -6897 14464
rect -6955 14396 -6897 14430
rect -6955 14362 -6943 14396
rect -6909 14362 -6897 14396
rect -6955 14328 -6897 14362
rect -6955 14294 -6943 14328
rect -6909 14294 -6897 14328
rect -6955 14260 -6897 14294
rect -6955 14226 -6943 14260
rect -6909 14226 -6897 14260
rect -6955 14192 -6897 14226
rect -6955 14158 -6943 14192
rect -6909 14158 -6897 14192
rect -6955 14124 -6897 14158
rect -6955 14090 -6943 14124
rect -6909 14090 -6897 14124
rect -6955 14056 -6897 14090
rect -6955 14022 -6943 14056
rect -6909 14022 -6897 14056
rect -6955 13988 -6897 14022
rect -6955 13954 -6943 13988
rect -6909 13954 -6897 13988
rect -6955 13920 -6897 13954
rect -6955 13886 -6943 13920
rect -6909 13886 -6897 13920
rect -6955 13852 -6897 13886
rect -6955 13818 -6943 13852
rect -6909 13818 -6897 13852
rect -6955 13784 -6897 13818
rect -6955 13750 -6943 13784
rect -6909 13750 -6897 13784
rect -6955 13716 -6897 13750
rect -6955 13682 -6943 13716
rect -6909 13682 -6897 13716
rect -6955 13648 -6897 13682
rect -6955 13614 -6943 13648
rect -6909 13614 -6897 13648
rect -6955 13580 -6897 13614
rect -6955 13546 -6943 13580
rect -6909 13546 -6897 13580
rect -6955 13512 -6897 13546
rect -6955 13478 -6943 13512
rect -6909 13478 -6897 13512
rect -6955 13444 -6897 13478
rect -6955 13410 -6943 13444
rect -6909 13410 -6897 13444
rect -6955 13376 -6897 13410
rect -6955 13342 -6943 13376
rect -6909 13342 -6897 13376
rect -6955 13308 -6897 13342
rect -6955 13274 -6943 13308
rect -6909 13274 -6897 13308
rect -6955 13240 -6897 13274
rect -6955 13206 -6943 13240
rect -6909 13206 -6897 13240
rect -6955 13172 -6897 13206
rect -6955 13138 -6943 13172
rect -6909 13138 -6897 13172
rect -6955 13104 -6897 13138
rect -6955 13070 -6943 13104
rect -6909 13070 -6897 13104
rect -6955 13036 -6897 13070
rect -6955 13002 -6943 13036
rect -6909 13002 -6897 13036
rect -6955 12968 -6897 13002
rect -6955 12934 -6943 12968
rect -6909 12934 -6897 12968
rect -6955 12900 -6897 12934
rect -6955 12866 -6943 12900
rect -6909 12866 -6897 12900
rect -6955 12835 -6897 12866
rect -6697 14804 -6639 14835
rect -6697 14770 -6685 14804
rect -6651 14770 -6639 14804
rect -6697 14736 -6639 14770
rect -6697 14702 -6685 14736
rect -6651 14702 -6639 14736
rect -6697 14668 -6639 14702
rect -6697 14634 -6685 14668
rect -6651 14634 -6639 14668
rect -6697 14600 -6639 14634
rect -6697 14566 -6685 14600
rect -6651 14566 -6639 14600
rect -6697 14532 -6639 14566
rect -6697 14498 -6685 14532
rect -6651 14498 -6639 14532
rect -6697 14464 -6639 14498
rect -6697 14430 -6685 14464
rect -6651 14430 -6639 14464
rect -6697 14396 -6639 14430
rect -6697 14362 -6685 14396
rect -6651 14362 -6639 14396
rect -6697 14328 -6639 14362
rect -6697 14294 -6685 14328
rect -6651 14294 -6639 14328
rect -6697 14260 -6639 14294
rect -6697 14226 -6685 14260
rect -6651 14226 -6639 14260
rect -6697 14192 -6639 14226
rect -6697 14158 -6685 14192
rect -6651 14158 -6639 14192
rect -6697 14124 -6639 14158
rect -6697 14090 -6685 14124
rect -6651 14090 -6639 14124
rect -6697 14056 -6639 14090
rect -6697 14022 -6685 14056
rect -6651 14022 -6639 14056
rect -6697 13988 -6639 14022
rect -6697 13954 -6685 13988
rect -6651 13954 -6639 13988
rect -6697 13920 -6639 13954
rect -6697 13886 -6685 13920
rect -6651 13886 -6639 13920
rect -6697 13852 -6639 13886
rect -6697 13818 -6685 13852
rect -6651 13818 -6639 13852
rect -6697 13784 -6639 13818
rect -6697 13750 -6685 13784
rect -6651 13750 -6639 13784
rect -6697 13716 -6639 13750
rect -6697 13682 -6685 13716
rect -6651 13682 -6639 13716
rect -6697 13648 -6639 13682
rect -6697 13614 -6685 13648
rect -6651 13614 -6639 13648
rect -6697 13580 -6639 13614
rect -6697 13546 -6685 13580
rect -6651 13546 -6639 13580
rect -6697 13512 -6639 13546
rect -6697 13478 -6685 13512
rect -6651 13478 -6639 13512
rect -6697 13444 -6639 13478
rect -6697 13410 -6685 13444
rect -6651 13410 -6639 13444
rect -6697 13376 -6639 13410
rect -6697 13342 -6685 13376
rect -6651 13342 -6639 13376
rect -6697 13308 -6639 13342
rect -6697 13274 -6685 13308
rect -6651 13274 -6639 13308
rect -6697 13240 -6639 13274
rect -6697 13206 -6685 13240
rect -6651 13206 -6639 13240
rect -6697 13172 -6639 13206
rect -6697 13138 -6685 13172
rect -6651 13138 -6639 13172
rect -6697 13104 -6639 13138
rect -6697 13070 -6685 13104
rect -6651 13070 -6639 13104
rect -6697 13036 -6639 13070
rect -6697 13002 -6685 13036
rect -6651 13002 -6639 13036
rect -6697 12968 -6639 13002
rect -6697 12934 -6685 12968
rect -6651 12934 -6639 12968
rect -6697 12900 -6639 12934
rect -6697 12866 -6685 12900
rect -6651 12866 -6639 12900
rect -6697 12835 -6639 12866
rect -6439 14804 -6381 14835
rect -6439 14770 -6427 14804
rect -6393 14770 -6381 14804
rect -6439 14736 -6381 14770
rect -6439 14702 -6427 14736
rect -6393 14702 -6381 14736
rect -6439 14668 -6381 14702
rect -6439 14634 -6427 14668
rect -6393 14634 -6381 14668
rect -6439 14600 -6381 14634
rect -6439 14566 -6427 14600
rect -6393 14566 -6381 14600
rect -6439 14532 -6381 14566
rect -6439 14498 -6427 14532
rect -6393 14498 -6381 14532
rect -6439 14464 -6381 14498
rect -6439 14430 -6427 14464
rect -6393 14430 -6381 14464
rect -6439 14396 -6381 14430
rect -6439 14362 -6427 14396
rect -6393 14362 -6381 14396
rect -6439 14328 -6381 14362
rect -6439 14294 -6427 14328
rect -6393 14294 -6381 14328
rect -6439 14260 -6381 14294
rect -6439 14226 -6427 14260
rect -6393 14226 -6381 14260
rect -6439 14192 -6381 14226
rect -6439 14158 -6427 14192
rect -6393 14158 -6381 14192
rect -6439 14124 -6381 14158
rect -6439 14090 -6427 14124
rect -6393 14090 -6381 14124
rect -6439 14056 -6381 14090
rect -6439 14022 -6427 14056
rect -6393 14022 -6381 14056
rect -6439 13988 -6381 14022
rect -6439 13954 -6427 13988
rect -6393 13954 -6381 13988
rect -6439 13920 -6381 13954
rect -6439 13886 -6427 13920
rect -6393 13886 -6381 13920
rect -6439 13852 -6381 13886
rect -6439 13818 -6427 13852
rect -6393 13818 -6381 13852
rect -6439 13784 -6381 13818
rect -6439 13750 -6427 13784
rect -6393 13750 -6381 13784
rect -6439 13716 -6381 13750
rect -6439 13682 -6427 13716
rect -6393 13682 -6381 13716
rect -6439 13648 -6381 13682
rect -6439 13614 -6427 13648
rect -6393 13614 -6381 13648
rect -6439 13580 -6381 13614
rect -6439 13546 -6427 13580
rect -6393 13546 -6381 13580
rect -6439 13512 -6381 13546
rect -6439 13478 -6427 13512
rect -6393 13478 -6381 13512
rect -6439 13444 -6381 13478
rect -6439 13410 -6427 13444
rect -6393 13410 -6381 13444
rect -6439 13376 -6381 13410
rect -6439 13342 -6427 13376
rect -6393 13342 -6381 13376
rect -6439 13308 -6381 13342
rect -6439 13274 -6427 13308
rect -6393 13274 -6381 13308
rect -6439 13240 -6381 13274
rect -6439 13206 -6427 13240
rect -6393 13206 -6381 13240
rect -6439 13172 -6381 13206
rect -6439 13138 -6427 13172
rect -6393 13138 -6381 13172
rect -6439 13104 -6381 13138
rect -6439 13070 -6427 13104
rect -6393 13070 -6381 13104
rect -6439 13036 -6381 13070
rect -6439 13002 -6427 13036
rect -6393 13002 -6381 13036
rect -6439 12968 -6381 13002
rect -6439 12934 -6427 12968
rect -6393 12934 -6381 12968
rect -6439 12900 -6381 12934
rect -6439 12866 -6427 12900
rect -6393 12866 -6381 12900
rect -6439 12835 -6381 12866
rect -6181 14804 -6123 14835
rect -6181 14770 -6169 14804
rect -6135 14770 -6123 14804
rect -6181 14736 -6123 14770
rect -6181 14702 -6169 14736
rect -6135 14702 -6123 14736
rect -6181 14668 -6123 14702
rect -6181 14634 -6169 14668
rect -6135 14634 -6123 14668
rect -6181 14600 -6123 14634
rect -6181 14566 -6169 14600
rect -6135 14566 -6123 14600
rect -6181 14532 -6123 14566
rect -6181 14498 -6169 14532
rect -6135 14498 -6123 14532
rect -6181 14464 -6123 14498
rect -6181 14430 -6169 14464
rect -6135 14430 -6123 14464
rect -6181 14396 -6123 14430
rect -6181 14362 -6169 14396
rect -6135 14362 -6123 14396
rect -6181 14328 -6123 14362
rect -6181 14294 -6169 14328
rect -6135 14294 -6123 14328
rect -6181 14260 -6123 14294
rect -6181 14226 -6169 14260
rect -6135 14226 -6123 14260
rect -6181 14192 -6123 14226
rect -6181 14158 -6169 14192
rect -6135 14158 -6123 14192
rect -6181 14124 -6123 14158
rect -6181 14090 -6169 14124
rect -6135 14090 -6123 14124
rect -6181 14056 -6123 14090
rect -6181 14022 -6169 14056
rect -6135 14022 -6123 14056
rect -6181 13988 -6123 14022
rect -6181 13954 -6169 13988
rect -6135 13954 -6123 13988
rect -6181 13920 -6123 13954
rect -6181 13886 -6169 13920
rect -6135 13886 -6123 13920
rect -6181 13852 -6123 13886
rect -6181 13818 -6169 13852
rect -6135 13818 -6123 13852
rect -6181 13784 -6123 13818
rect -6181 13750 -6169 13784
rect -6135 13750 -6123 13784
rect -6181 13716 -6123 13750
rect -6181 13682 -6169 13716
rect -6135 13682 -6123 13716
rect -6181 13648 -6123 13682
rect -6181 13614 -6169 13648
rect -6135 13614 -6123 13648
rect -6181 13580 -6123 13614
rect -6181 13546 -6169 13580
rect -6135 13546 -6123 13580
rect -6181 13512 -6123 13546
rect -6181 13478 -6169 13512
rect -6135 13478 -6123 13512
rect -6181 13444 -6123 13478
rect -6181 13410 -6169 13444
rect -6135 13410 -6123 13444
rect -6181 13376 -6123 13410
rect -6181 13342 -6169 13376
rect -6135 13342 -6123 13376
rect -6181 13308 -6123 13342
rect -6181 13274 -6169 13308
rect -6135 13274 -6123 13308
rect -6181 13240 -6123 13274
rect -6181 13206 -6169 13240
rect -6135 13206 -6123 13240
rect -6181 13172 -6123 13206
rect -6181 13138 -6169 13172
rect -6135 13138 -6123 13172
rect -6181 13104 -6123 13138
rect -6181 13070 -6169 13104
rect -6135 13070 -6123 13104
rect -6181 13036 -6123 13070
rect -6181 13002 -6169 13036
rect -6135 13002 -6123 13036
rect -6181 12968 -6123 13002
rect -6181 12934 -6169 12968
rect -6135 12934 -6123 12968
rect -6181 12900 -6123 12934
rect -6181 12866 -6169 12900
rect -6135 12866 -6123 12900
rect -6181 12835 -6123 12866
rect -5923 14804 -5865 14835
rect -5923 14770 -5911 14804
rect -5877 14770 -5865 14804
rect -5923 14736 -5865 14770
rect -5923 14702 -5911 14736
rect -5877 14702 -5865 14736
rect -5923 14668 -5865 14702
rect -5923 14634 -5911 14668
rect -5877 14634 -5865 14668
rect -5923 14600 -5865 14634
rect -5923 14566 -5911 14600
rect -5877 14566 -5865 14600
rect -5923 14532 -5865 14566
rect -5923 14498 -5911 14532
rect -5877 14498 -5865 14532
rect -5923 14464 -5865 14498
rect -5923 14430 -5911 14464
rect -5877 14430 -5865 14464
rect -5923 14396 -5865 14430
rect -5923 14362 -5911 14396
rect -5877 14362 -5865 14396
rect -5923 14328 -5865 14362
rect -5923 14294 -5911 14328
rect -5877 14294 -5865 14328
rect -5923 14260 -5865 14294
rect -5923 14226 -5911 14260
rect -5877 14226 -5865 14260
rect -5923 14192 -5865 14226
rect -5923 14158 -5911 14192
rect -5877 14158 -5865 14192
rect -5923 14124 -5865 14158
rect -5923 14090 -5911 14124
rect -5877 14090 -5865 14124
rect -5923 14056 -5865 14090
rect -5923 14022 -5911 14056
rect -5877 14022 -5865 14056
rect -5923 13988 -5865 14022
rect -5923 13954 -5911 13988
rect -5877 13954 -5865 13988
rect -5923 13920 -5865 13954
rect -5923 13886 -5911 13920
rect -5877 13886 -5865 13920
rect -5923 13852 -5865 13886
rect -5923 13818 -5911 13852
rect -5877 13818 -5865 13852
rect -5923 13784 -5865 13818
rect -5923 13750 -5911 13784
rect -5877 13750 -5865 13784
rect -5923 13716 -5865 13750
rect -5923 13682 -5911 13716
rect -5877 13682 -5865 13716
rect -5923 13648 -5865 13682
rect -5923 13614 -5911 13648
rect -5877 13614 -5865 13648
rect -5923 13580 -5865 13614
rect -5923 13546 -5911 13580
rect -5877 13546 -5865 13580
rect -5923 13512 -5865 13546
rect -5923 13478 -5911 13512
rect -5877 13478 -5865 13512
rect -5923 13444 -5865 13478
rect -5923 13410 -5911 13444
rect -5877 13410 -5865 13444
rect -5923 13376 -5865 13410
rect -5923 13342 -5911 13376
rect -5877 13342 -5865 13376
rect -5923 13308 -5865 13342
rect -5923 13274 -5911 13308
rect -5877 13274 -5865 13308
rect -5923 13240 -5865 13274
rect -5923 13206 -5911 13240
rect -5877 13206 -5865 13240
rect -5923 13172 -5865 13206
rect -5923 13138 -5911 13172
rect -5877 13138 -5865 13172
rect -5923 13104 -5865 13138
rect -5923 13070 -5911 13104
rect -5877 13070 -5865 13104
rect -5923 13036 -5865 13070
rect -5923 13002 -5911 13036
rect -5877 13002 -5865 13036
rect -5923 12968 -5865 13002
rect -5923 12934 -5911 12968
rect -5877 12934 -5865 12968
rect -5923 12900 -5865 12934
rect -5923 12866 -5911 12900
rect -5877 12866 -5865 12900
rect -5923 12835 -5865 12866
rect -5665 14804 -5607 14835
rect -5665 14770 -5653 14804
rect -5619 14770 -5607 14804
rect -5665 14736 -5607 14770
rect -5665 14702 -5653 14736
rect -5619 14702 -5607 14736
rect -5665 14668 -5607 14702
rect -5665 14634 -5653 14668
rect -5619 14634 -5607 14668
rect -5665 14600 -5607 14634
rect -5665 14566 -5653 14600
rect -5619 14566 -5607 14600
rect -5665 14532 -5607 14566
rect -5665 14498 -5653 14532
rect -5619 14498 -5607 14532
rect -5665 14464 -5607 14498
rect -5665 14430 -5653 14464
rect -5619 14430 -5607 14464
rect -5665 14396 -5607 14430
rect -5665 14362 -5653 14396
rect -5619 14362 -5607 14396
rect -5665 14328 -5607 14362
rect -5665 14294 -5653 14328
rect -5619 14294 -5607 14328
rect -5665 14260 -5607 14294
rect -5665 14226 -5653 14260
rect -5619 14226 -5607 14260
rect -5665 14192 -5607 14226
rect -5665 14158 -5653 14192
rect -5619 14158 -5607 14192
rect -5665 14124 -5607 14158
rect -5665 14090 -5653 14124
rect -5619 14090 -5607 14124
rect -5665 14056 -5607 14090
rect -5665 14022 -5653 14056
rect -5619 14022 -5607 14056
rect -5665 13988 -5607 14022
rect -5665 13954 -5653 13988
rect -5619 13954 -5607 13988
rect -5665 13920 -5607 13954
rect -5665 13886 -5653 13920
rect -5619 13886 -5607 13920
rect -5665 13852 -5607 13886
rect -5665 13818 -5653 13852
rect -5619 13818 -5607 13852
rect -5665 13784 -5607 13818
rect -5665 13750 -5653 13784
rect -5619 13750 -5607 13784
rect -5665 13716 -5607 13750
rect -5665 13682 -5653 13716
rect -5619 13682 -5607 13716
rect -5665 13648 -5607 13682
rect -5665 13614 -5653 13648
rect -5619 13614 -5607 13648
rect -5665 13580 -5607 13614
rect -5665 13546 -5653 13580
rect -5619 13546 -5607 13580
rect -5665 13512 -5607 13546
rect -5665 13478 -5653 13512
rect -5619 13478 -5607 13512
rect -5665 13444 -5607 13478
rect -5665 13410 -5653 13444
rect -5619 13410 -5607 13444
rect -5665 13376 -5607 13410
rect -5665 13342 -5653 13376
rect -5619 13342 -5607 13376
rect -5665 13308 -5607 13342
rect -5665 13274 -5653 13308
rect -5619 13274 -5607 13308
rect -5665 13240 -5607 13274
rect -5665 13206 -5653 13240
rect -5619 13206 -5607 13240
rect -5665 13172 -5607 13206
rect -5665 13138 -5653 13172
rect -5619 13138 -5607 13172
rect -5665 13104 -5607 13138
rect -5665 13070 -5653 13104
rect -5619 13070 -5607 13104
rect -5665 13036 -5607 13070
rect -5665 13002 -5653 13036
rect -5619 13002 -5607 13036
rect -5665 12968 -5607 13002
rect -5665 12934 -5653 12968
rect -5619 12934 -5607 12968
rect -5665 12900 -5607 12934
rect -5665 12866 -5653 12900
rect -5619 12866 -5607 12900
rect -5665 12835 -5607 12866
rect -5407 14804 -5349 14835
rect -5407 14770 -5395 14804
rect -5361 14770 -5349 14804
rect -5407 14736 -5349 14770
rect -5407 14702 -5395 14736
rect -5361 14702 -5349 14736
rect -5407 14668 -5349 14702
rect -5407 14634 -5395 14668
rect -5361 14634 -5349 14668
rect -5407 14600 -5349 14634
rect -5407 14566 -5395 14600
rect -5361 14566 -5349 14600
rect -5407 14532 -5349 14566
rect -5407 14498 -5395 14532
rect -5361 14498 -5349 14532
rect -5407 14464 -5349 14498
rect -5407 14430 -5395 14464
rect -5361 14430 -5349 14464
rect -5407 14396 -5349 14430
rect -5407 14362 -5395 14396
rect -5361 14362 -5349 14396
rect -5407 14328 -5349 14362
rect -5407 14294 -5395 14328
rect -5361 14294 -5349 14328
rect -5407 14260 -5349 14294
rect -5407 14226 -5395 14260
rect -5361 14226 -5349 14260
rect -5407 14192 -5349 14226
rect -5407 14158 -5395 14192
rect -5361 14158 -5349 14192
rect -5407 14124 -5349 14158
rect -5407 14090 -5395 14124
rect -5361 14090 -5349 14124
rect -5407 14056 -5349 14090
rect -5407 14022 -5395 14056
rect -5361 14022 -5349 14056
rect -5407 13988 -5349 14022
rect -5407 13954 -5395 13988
rect -5361 13954 -5349 13988
rect -5407 13920 -5349 13954
rect -5407 13886 -5395 13920
rect -5361 13886 -5349 13920
rect -5407 13852 -5349 13886
rect -5407 13818 -5395 13852
rect -5361 13818 -5349 13852
rect -5407 13784 -5349 13818
rect -5407 13750 -5395 13784
rect -5361 13750 -5349 13784
rect -5407 13716 -5349 13750
rect -5407 13682 -5395 13716
rect -5361 13682 -5349 13716
rect -5407 13648 -5349 13682
rect -5407 13614 -5395 13648
rect -5361 13614 -5349 13648
rect -5407 13580 -5349 13614
rect -5407 13546 -5395 13580
rect -5361 13546 -5349 13580
rect -5407 13512 -5349 13546
rect -5407 13478 -5395 13512
rect -5361 13478 -5349 13512
rect -5407 13444 -5349 13478
rect -5407 13410 -5395 13444
rect -5361 13410 -5349 13444
rect -5407 13376 -5349 13410
rect -5407 13342 -5395 13376
rect -5361 13342 -5349 13376
rect -5407 13308 -5349 13342
rect -5407 13274 -5395 13308
rect -5361 13274 -5349 13308
rect -5407 13240 -5349 13274
rect -5407 13206 -5395 13240
rect -5361 13206 -5349 13240
rect -5407 13172 -5349 13206
rect -5407 13138 -5395 13172
rect -5361 13138 -5349 13172
rect -5407 13104 -5349 13138
rect -5407 13070 -5395 13104
rect -5361 13070 -5349 13104
rect -5407 13036 -5349 13070
rect -5407 13002 -5395 13036
rect -5361 13002 -5349 13036
rect -5407 12968 -5349 13002
rect -5407 12934 -5395 12968
rect -5361 12934 -5349 12968
rect -5407 12900 -5349 12934
rect -5407 12866 -5395 12900
rect -5361 12866 -5349 12900
rect -5407 12835 -5349 12866
rect -5149 14804 -5091 14835
rect -5149 14770 -5137 14804
rect -5103 14770 -5091 14804
rect -5149 14736 -5091 14770
rect -5149 14702 -5137 14736
rect -5103 14702 -5091 14736
rect -5149 14668 -5091 14702
rect -5149 14634 -5137 14668
rect -5103 14634 -5091 14668
rect -5149 14600 -5091 14634
rect -5149 14566 -5137 14600
rect -5103 14566 -5091 14600
rect -5149 14532 -5091 14566
rect -5149 14498 -5137 14532
rect -5103 14498 -5091 14532
rect -5149 14464 -5091 14498
rect -5149 14430 -5137 14464
rect -5103 14430 -5091 14464
rect -5149 14396 -5091 14430
rect -5149 14362 -5137 14396
rect -5103 14362 -5091 14396
rect -5149 14328 -5091 14362
rect -5149 14294 -5137 14328
rect -5103 14294 -5091 14328
rect -5149 14260 -5091 14294
rect -5149 14226 -5137 14260
rect -5103 14226 -5091 14260
rect -5149 14192 -5091 14226
rect -5149 14158 -5137 14192
rect -5103 14158 -5091 14192
rect -5149 14124 -5091 14158
rect -5149 14090 -5137 14124
rect -5103 14090 -5091 14124
rect -5149 14056 -5091 14090
rect -5149 14022 -5137 14056
rect -5103 14022 -5091 14056
rect -5149 13988 -5091 14022
rect -5149 13954 -5137 13988
rect -5103 13954 -5091 13988
rect -5149 13920 -5091 13954
rect -5149 13886 -5137 13920
rect -5103 13886 -5091 13920
rect -5149 13852 -5091 13886
rect -5149 13818 -5137 13852
rect -5103 13818 -5091 13852
rect -5149 13784 -5091 13818
rect -5149 13750 -5137 13784
rect -5103 13750 -5091 13784
rect -5149 13716 -5091 13750
rect -5149 13682 -5137 13716
rect -5103 13682 -5091 13716
rect -5149 13648 -5091 13682
rect -5149 13614 -5137 13648
rect -5103 13614 -5091 13648
rect -5149 13580 -5091 13614
rect -5149 13546 -5137 13580
rect -5103 13546 -5091 13580
rect -5149 13512 -5091 13546
rect -5149 13478 -5137 13512
rect -5103 13478 -5091 13512
rect -5149 13444 -5091 13478
rect -5149 13410 -5137 13444
rect -5103 13410 -5091 13444
rect -5149 13376 -5091 13410
rect -5149 13342 -5137 13376
rect -5103 13342 -5091 13376
rect -5149 13308 -5091 13342
rect -5149 13274 -5137 13308
rect -5103 13274 -5091 13308
rect -5149 13240 -5091 13274
rect -5149 13206 -5137 13240
rect -5103 13206 -5091 13240
rect -5149 13172 -5091 13206
rect -5149 13138 -5137 13172
rect -5103 13138 -5091 13172
rect -5149 13104 -5091 13138
rect -5149 13070 -5137 13104
rect -5103 13070 -5091 13104
rect -5149 13036 -5091 13070
rect -5149 13002 -5137 13036
rect -5103 13002 -5091 13036
rect -5149 12968 -5091 13002
rect -5149 12934 -5137 12968
rect -5103 12934 -5091 12968
rect -5149 12900 -5091 12934
rect -5149 12866 -5137 12900
rect -5103 12866 -5091 12900
rect -5149 12835 -5091 12866
rect -4891 14804 -4833 14835
rect -4891 14770 -4879 14804
rect -4845 14770 -4833 14804
rect -4891 14736 -4833 14770
rect -4891 14702 -4879 14736
rect -4845 14702 -4833 14736
rect -4891 14668 -4833 14702
rect -4891 14634 -4879 14668
rect -4845 14634 -4833 14668
rect -4891 14600 -4833 14634
rect -4891 14566 -4879 14600
rect -4845 14566 -4833 14600
rect -4891 14532 -4833 14566
rect -4891 14498 -4879 14532
rect -4845 14498 -4833 14532
rect -4891 14464 -4833 14498
rect -4891 14430 -4879 14464
rect -4845 14430 -4833 14464
rect -4891 14396 -4833 14430
rect -4891 14362 -4879 14396
rect -4845 14362 -4833 14396
rect -4891 14328 -4833 14362
rect -4891 14294 -4879 14328
rect -4845 14294 -4833 14328
rect -4891 14260 -4833 14294
rect -4891 14226 -4879 14260
rect -4845 14226 -4833 14260
rect -4891 14192 -4833 14226
rect -4891 14158 -4879 14192
rect -4845 14158 -4833 14192
rect -4891 14124 -4833 14158
rect -4891 14090 -4879 14124
rect -4845 14090 -4833 14124
rect -4891 14056 -4833 14090
rect -4891 14022 -4879 14056
rect -4845 14022 -4833 14056
rect -4891 13988 -4833 14022
rect -4891 13954 -4879 13988
rect -4845 13954 -4833 13988
rect -4891 13920 -4833 13954
rect -4891 13886 -4879 13920
rect -4845 13886 -4833 13920
rect -4891 13852 -4833 13886
rect -4891 13818 -4879 13852
rect -4845 13818 -4833 13852
rect -4891 13784 -4833 13818
rect -4891 13750 -4879 13784
rect -4845 13750 -4833 13784
rect -4891 13716 -4833 13750
rect -4891 13682 -4879 13716
rect -4845 13682 -4833 13716
rect -4891 13648 -4833 13682
rect -4891 13614 -4879 13648
rect -4845 13614 -4833 13648
rect -4891 13580 -4833 13614
rect -4891 13546 -4879 13580
rect -4845 13546 -4833 13580
rect -4891 13512 -4833 13546
rect -4891 13478 -4879 13512
rect -4845 13478 -4833 13512
rect -4891 13444 -4833 13478
rect -4891 13410 -4879 13444
rect -4845 13410 -4833 13444
rect -4891 13376 -4833 13410
rect -4891 13342 -4879 13376
rect -4845 13342 -4833 13376
rect -4891 13308 -4833 13342
rect -4891 13274 -4879 13308
rect -4845 13274 -4833 13308
rect -4891 13240 -4833 13274
rect -4891 13206 -4879 13240
rect -4845 13206 -4833 13240
rect -4891 13172 -4833 13206
rect -4891 13138 -4879 13172
rect -4845 13138 -4833 13172
rect -4891 13104 -4833 13138
rect -4891 13070 -4879 13104
rect -4845 13070 -4833 13104
rect -4891 13036 -4833 13070
rect -4891 13002 -4879 13036
rect -4845 13002 -4833 13036
rect -4891 12968 -4833 13002
rect -4891 12934 -4879 12968
rect -4845 12934 -4833 12968
rect -4891 12900 -4833 12934
rect -4891 12866 -4879 12900
rect -4845 12866 -4833 12900
rect -4891 12835 -4833 12866
rect -8827 11123 -8769 11164
rect -8827 11089 -8815 11123
rect -8781 11089 -8769 11123
rect -8827 11055 -8769 11089
rect -8827 11021 -8815 11055
rect -8781 11021 -8769 11055
rect -8827 10987 -8769 11021
rect -8827 10953 -8815 10987
rect -8781 10953 -8769 10987
rect -8827 10919 -8769 10953
rect -8827 10885 -8815 10919
rect -8781 10885 -8769 10919
rect -8827 10851 -8769 10885
rect -8827 10817 -8815 10851
rect -8781 10817 -8769 10851
rect -8827 10783 -8769 10817
rect -8827 10749 -8815 10783
rect -8781 10749 -8769 10783
rect -8827 10715 -8769 10749
rect -8827 10681 -8815 10715
rect -8781 10681 -8769 10715
rect -8827 10647 -8769 10681
rect -8827 10613 -8815 10647
rect -8781 10613 -8769 10647
rect -8827 10579 -8769 10613
rect -8827 10545 -8815 10579
rect -8781 10545 -8769 10579
rect -8827 10511 -8769 10545
rect -8827 10477 -8815 10511
rect -8781 10477 -8769 10511
rect -8827 10443 -8769 10477
rect -8827 10409 -8815 10443
rect -8781 10409 -8769 10443
rect -8827 10375 -8769 10409
rect -8827 10341 -8815 10375
rect -8781 10341 -8769 10375
rect -8827 10307 -8769 10341
rect -8827 10273 -8815 10307
rect -8781 10273 -8769 10307
rect -8827 10239 -8769 10273
rect -8827 10205 -8815 10239
rect -8781 10205 -8769 10239
rect -8827 10164 -8769 10205
rect -8569 11123 -8511 11164
rect -8569 11089 -8557 11123
rect -8523 11089 -8511 11123
rect -8569 11055 -8511 11089
rect -8569 11021 -8557 11055
rect -8523 11021 -8511 11055
rect -8569 10987 -8511 11021
rect -8569 10953 -8557 10987
rect -8523 10953 -8511 10987
rect -8569 10919 -8511 10953
rect -8569 10885 -8557 10919
rect -8523 10885 -8511 10919
rect -8569 10851 -8511 10885
rect -8569 10817 -8557 10851
rect -8523 10817 -8511 10851
rect -8569 10783 -8511 10817
rect -8569 10749 -8557 10783
rect -8523 10749 -8511 10783
rect -8569 10715 -8511 10749
rect -8569 10681 -8557 10715
rect -8523 10681 -8511 10715
rect -8569 10647 -8511 10681
rect -8569 10613 -8557 10647
rect -8523 10613 -8511 10647
rect -8569 10579 -8511 10613
rect -8569 10545 -8557 10579
rect -8523 10545 -8511 10579
rect -8569 10511 -8511 10545
rect -8569 10477 -8557 10511
rect -8523 10477 -8511 10511
rect -8569 10443 -8511 10477
rect -8569 10409 -8557 10443
rect -8523 10409 -8511 10443
rect -8569 10375 -8511 10409
rect -8569 10341 -8557 10375
rect -8523 10341 -8511 10375
rect -8569 10307 -8511 10341
rect -8569 10273 -8557 10307
rect -8523 10273 -8511 10307
rect -8569 10239 -8511 10273
rect -8569 10205 -8557 10239
rect -8523 10205 -8511 10239
rect -8569 10164 -8511 10205
rect -8311 11123 -8253 11164
rect -8311 11089 -8299 11123
rect -8265 11089 -8253 11123
rect -8311 11055 -8253 11089
rect -8311 11021 -8299 11055
rect -8265 11021 -8253 11055
rect -8311 10987 -8253 11021
rect -8311 10953 -8299 10987
rect -8265 10953 -8253 10987
rect -8311 10919 -8253 10953
rect -8311 10885 -8299 10919
rect -8265 10885 -8253 10919
rect -8311 10851 -8253 10885
rect -8311 10817 -8299 10851
rect -8265 10817 -8253 10851
rect -8311 10783 -8253 10817
rect -8311 10749 -8299 10783
rect -8265 10749 -8253 10783
rect -8311 10715 -8253 10749
rect -8311 10681 -8299 10715
rect -8265 10681 -8253 10715
rect -8311 10647 -8253 10681
rect -8311 10613 -8299 10647
rect -8265 10613 -8253 10647
rect -8311 10579 -8253 10613
rect -8311 10545 -8299 10579
rect -8265 10545 -8253 10579
rect -8311 10511 -8253 10545
rect -8311 10477 -8299 10511
rect -8265 10477 -8253 10511
rect -8311 10443 -8253 10477
rect -8311 10409 -8299 10443
rect -8265 10409 -8253 10443
rect -8311 10375 -8253 10409
rect -8311 10341 -8299 10375
rect -8265 10341 -8253 10375
rect -8311 10307 -8253 10341
rect -8311 10273 -8299 10307
rect -8265 10273 -8253 10307
rect -8311 10239 -8253 10273
rect -8311 10205 -8299 10239
rect -8265 10205 -8253 10239
rect -8311 10164 -8253 10205
rect -8053 11123 -7995 11164
rect -8053 11089 -8041 11123
rect -8007 11089 -7995 11123
rect -8053 11055 -7995 11089
rect -8053 11021 -8041 11055
rect -8007 11021 -7995 11055
rect -8053 10987 -7995 11021
rect -8053 10953 -8041 10987
rect -8007 10953 -7995 10987
rect -8053 10919 -7995 10953
rect -8053 10885 -8041 10919
rect -8007 10885 -7995 10919
rect -8053 10851 -7995 10885
rect -8053 10817 -8041 10851
rect -8007 10817 -7995 10851
rect -8053 10783 -7995 10817
rect -8053 10749 -8041 10783
rect -8007 10749 -7995 10783
rect -8053 10715 -7995 10749
rect -8053 10681 -8041 10715
rect -8007 10681 -7995 10715
rect -8053 10647 -7995 10681
rect -8053 10613 -8041 10647
rect -8007 10613 -7995 10647
rect -8053 10579 -7995 10613
rect -8053 10545 -8041 10579
rect -8007 10545 -7995 10579
rect -8053 10511 -7995 10545
rect -8053 10477 -8041 10511
rect -8007 10477 -7995 10511
rect -8053 10443 -7995 10477
rect -8053 10409 -8041 10443
rect -8007 10409 -7995 10443
rect -8053 10375 -7995 10409
rect -8053 10341 -8041 10375
rect -8007 10341 -7995 10375
rect -8053 10307 -7995 10341
rect -8053 10273 -8041 10307
rect -8007 10273 -7995 10307
rect -8053 10239 -7995 10273
rect -8053 10205 -8041 10239
rect -8007 10205 -7995 10239
rect -8053 10164 -7995 10205
rect -7795 11123 -7737 11164
rect -7795 11089 -7783 11123
rect -7749 11089 -7737 11123
rect -7795 11055 -7737 11089
rect -7795 11021 -7783 11055
rect -7749 11021 -7737 11055
rect -7795 10987 -7737 11021
rect -7795 10953 -7783 10987
rect -7749 10953 -7737 10987
rect -7795 10919 -7737 10953
rect -7795 10885 -7783 10919
rect -7749 10885 -7737 10919
rect -7795 10851 -7737 10885
rect -7795 10817 -7783 10851
rect -7749 10817 -7737 10851
rect -7795 10783 -7737 10817
rect -7795 10749 -7783 10783
rect -7749 10749 -7737 10783
rect -7795 10715 -7737 10749
rect -7795 10681 -7783 10715
rect -7749 10681 -7737 10715
rect -7795 10647 -7737 10681
rect -7795 10613 -7783 10647
rect -7749 10613 -7737 10647
rect -7795 10579 -7737 10613
rect -7795 10545 -7783 10579
rect -7749 10545 -7737 10579
rect -7795 10511 -7737 10545
rect -7795 10477 -7783 10511
rect -7749 10477 -7737 10511
rect -7795 10443 -7737 10477
rect -7795 10409 -7783 10443
rect -7749 10409 -7737 10443
rect -7795 10375 -7737 10409
rect -7795 10341 -7783 10375
rect -7749 10341 -7737 10375
rect -7795 10307 -7737 10341
rect -7795 10273 -7783 10307
rect -7749 10273 -7737 10307
rect -7795 10239 -7737 10273
rect -7795 10205 -7783 10239
rect -7749 10205 -7737 10239
rect -7795 10164 -7737 10205
rect -7537 11123 -7479 11164
rect -7537 11089 -7525 11123
rect -7491 11089 -7479 11123
rect -7537 11055 -7479 11089
rect -7537 11021 -7525 11055
rect -7491 11021 -7479 11055
rect -7537 10987 -7479 11021
rect -7537 10953 -7525 10987
rect -7491 10953 -7479 10987
rect -7537 10919 -7479 10953
rect -7537 10885 -7525 10919
rect -7491 10885 -7479 10919
rect -7537 10851 -7479 10885
rect -7537 10817 -7525 10851
rect -7491 10817 -7479 10851
rect -7537 10783 -7479 10817
rect -7537 10749 -7525 10783
rect -7491 10749 -7479 10783
rect -7537 10715 -7479 10749
rect -7537 10681 -7525 10715
rect -7491 10681 -7479 10715
rect -7537 10647 -7479 10681
rect -7537 10613 -7525 10647
rect -7491 10613 -7479 10647
rect -7537 10579 -7479 10613
rect -7537 10545 -7525 10579
rect -7491 10545 -7479 10579
rect -7537 10511 -7479 10545
rect -7537 10477 -7525 10511
rect -7491 10477 -7479 10511
rect -7537 10443 -7479 10477
rect -7537 10409 -7525 10443
rect -7491 10409 -7479 10443
rect -7537 10375 -7479 10409
rect -7537 10341 -7525 10375
rect -7491 10341 -7479 10375
rect -7537 10307 -7479 10341
rect -7537 10273 -7525 10307
rect -7491 10273 -7479 10307
rect -7537 10239 -7479 10273
rect -7537 10205 -7525 10239
rect -7491 10205 -7479 10239
rect -7537 10164 -7479 10205
rect -7279 11123 -7221 11164
rect -7279 11089 -7267 11123
rect -7233 11089 -7221 11123
rect -7279 11055 -7221 11089
rect -7279 11021 -7267 11055
rect -7233 11021 -7221 11055
rect -7279 10987 -7221 11021
rect -7279 10953 -7267 10987
rect -7233 10953 -7221 10987
rect -7279 10919 -7221 10953
rect -7279 10885 -7267 10919
rect -7233 10885 -7221 10919
rect -7279 10851 -7221 10885
rect -7279 10817 -7267 10851
rect -7233 10817 -7221 10851
rect -7279 10783 -7221 10817
rect -7279 10749 -7267 10783
rect -7233 10749 -7221 10783
rect -7279 10715 -7221 10749
rect -7279 10681 -7267 10715
rect -7233 10681 -7221 10715
rect -7279 10647 -7221 10681
rect -7279 10613 -7267 10647
rect -7233 10613 -7221 10647
rect -7279 10579 -7221 10613
rect -7279 10545 -7267 10579
rect -7233 10545 -7221 10579
rect -7279 10511 -7221 10545
rect -7279 10477 -7267 10511
rect -7233 10477 -7221 10511
rect -7279 10443 -7221 10477
rect -7279 10409 -7267 10443
rect -7233 10409 -7221 10443
rect -7279 10375 -7221 10409
rect -7279 10341 -7267 10375
rect -7233 10341 -7221 10375
rect -7279 10307 -7221 10341
rect -7279 10273 -7267 10307
rect -7233 10273 -7221 10307
rect -7279 10239 -7221 10273
rect -7279 10205 -7267 10239
rect -7233 10205 -7221 10239
rect -7279 10164 -7221 10205
rect -7021 11123 -6963 11164
rect -7021 11089 -7009 11123
rect -6975 11089 -6963 11123
rect -7021 11055 -6963 11089
rect -7021 11021 -7009 11055
rect -6975 11021 -6963 11055
rect -7021 10987 -6963 11021
rect -7021 10953 -7009 10987
rect -6975 10953 -6963 10987
rect -7021 10919 -6963 10953
rect -7021 10885 -7009 10919
rect -6975 10885 -6963 10919
rect -7021 10851 -6963 10885
rect -7021 10817 -7009 10851
rect -6975 10817 -6963 10851
rect -7021 10783 -6963 10817
rect -7021 10749 -7009 10783
rect -6975 10749 -6963 10783
rect -7021 10715 -6963 10749
rect -7021 10681 -7009 10715
rect -6975 10681 -6963 10715
rect -7021 10647 -6963 10681
rect -7021 10613 -7009 10647
rect -6975 10613 -6963 10647
rect -7021 10579 -6963 10613
rect -7021 10545 -7009 10579
rect -6975 10545 -6963 10579
rect -7021 10511 -6963 10545
rect -7021 10477 -7009 10511
rect -6975 10477 -6963 10511
rect -7021 10443 -6963 10477
rect -7021 10409 -7009 10443
rect -6975 10409 -6963 10443
rect -7021 10375 -6963 10409
rect -7021 10341 -7009 10375
rect -6975 10341 -6963 10375
rect -7021 10307 -6963 10341
rect -7021 10273 -7009 10307
rect -6975 10273 -6963 10307
rect -7021 10239 -6963 10273
rect -7021 10205 -7009 10239
rect -6975 10205 -6963 10239
rect -7021 10164 -6963 10205
rect -6763 11123 -6705 11164
rect -6763 11089 -6751 11123
rect -6717 11089 -6705 11123
rect -6763 11055 -6705 11089
rect -6763 11021 -6751 11055
rect -6717 11021 -6705 11055
rect -6763 10987 -6705 11021
rect -6763 10953 -6751 10987
rect -6717 10953 -6705 10987
rect -6763 10919 -6705 10953
rect -6763 10885 -6751 10919
rect -6717 10885 -6705 10919
rect -6763 10851 -6705 10885
rect -6763 10817 -6751 10851
rect -6717 10817 -6705 10851
rect -6763 10783 -6705 10817
rect -6763 10749 -6751 10783
rect -6717 10749 -6705 10783
rect -6763 10715 -6705 10749
rect -6763 10681 -6751 10715
rect -6717 10681 -6705 10715
rect -6763 10647 -6705 10681
rect -6763 10613 -6751 10647
rect -6717 10613 -6705 10647
rect -6763 10579 -6705 10613
rect -6763 10545 -6751 10579
rect -6717 10545 -6705 10579
rect -6763 10511 -6705 10545
rect -6763 10477 -6751 10511
rect -6717 10477 -6705 10511
rect -6763 10443 -6705 10477
rect -6763 10409 -6751 10443
rect -6717 10409 -6705 10443
rect -6763 10375 -6705 10409
rect -6763 10341 -6751 10375
rect -6717 10341 -6705 10375
rect -6763 10307 -6705 10341
rect -6763 10273 -6751 10307
rect -6717 10273 -6705 10307
rect -6763 10239 -6705 10273
rect -6763 10205 -6751 10239
rect -6717 10205 -6705 10239
rect -6763 10164 -6705 10205
rect -6505 11123 -6447 11164
rect -6505 11089 -6493 11123
rect -6459 11089 -6447 11123
rect -6505 11055 -6447 11089
rect -6505 11021 -6493 11055
rect -6459 11021 -6447 11055
rect -6505 10987 -6447 11021
rect -6505 10953 -6493 10987
rect -6459 10953 -6447 10987
rect -6505 10919 -6447 10953
rect -6505 10885 -6493 10919
rect -6459 10885 -6447 10919
rect -6505 10851 -6447 10885
rect -6505 10817 -6493 10851
rect -6459 10817 -6447 10851
rect -6505 10783 -6447 10817
rect -6505 10749 -6493 10783
rect -6459 10749 -6447 10783
rect -6505 10715 -6447 10749
rect -6505 10681 -6493 10715
rect -6459 10681 -6447 10715
rect -6505 10647 -6447 10681
rect -6505 10613 -6493 10647
rect -6459 10613 -6447 10647
rect -6505 10579 -6447 10613
rect -6505 10545 -6493 10579
rect -6459 10545 -6447 10579
rect -6505 10511 -6447 10545
rect -6505 10477 -6493 10511
rect -6459 10477 -6447 10511
rect -6505 10443 -6447 10477
rect -6505 10409 -6493 10443
rect -6459 10409 -6447 10443
rect -6505 10375 -6447 10409
rect -6505 10341 -6493 10375
rect -6459 10341 -6447 10375
rect -6505 10307 -6447 10341
rect -6505 10273 -6493 10307
rect -6459 10273 -6447 10307
rect -6505 10239 -6447 10273
rect -6505 10205 -6493 10239
rect -6459 10205 -6447 10239
rect -6505 10164 -6447 10205
rect -6247 11123 -6189 11164
rect -6247 11089 -6235 11123
rect -6201 11089 -6189 11123
rect -6247 11055 -6189 11089
rect -6247 11021 -6235 11055
rect -6201 11021 -6189 11055
rect -6247 10987 -6189 11021
rect -6247 10953 -6235 10987
rect -6201 10953 -6189 10987
rect -6247 10919 -6189 10953
rect -6247 10885 -6235 10919
rect -6201 10885 -6189 10919
rect -6247 10851 -6189 10885
rect -6247 10817 -6235 10851
rect -6201 10817 -6189 10851
rect -6247 10783 -6189 10817
rect -6247 10749 -6235 10783
rect -6201 10749 -6189 10783
rect -6247 10715 -6189 10749
rect -6247 10681 -6235 10715
rect -6201 10681 -6189 10715
rect -6247 10647 -6189 10681
rect -6247 10613 -6235 10647
rect -6201 10613 -6189 10647
rect -6247 10579 -6189 10613
rect -6247 10545 -6235 10579
rect -6201 10545 -6189 10579
rect -6247 10511 -6189 10545
rect -6247 10477 -6235 10511
rect -6201 10477 -6189 10511
rect -6247 10443 -6189 10477
rect -6247 10409 -6235 10443
rect -6201 10409 -6189 10443
rect -6247 10375 -6189 10409
rect -6247 10341 -6235 10375
rect -6201 10341 -6189 10375
rect -6247 10307 -6189 10341
rect -6247 10273 -6235 10307
rect -6201 10273 -6189 10307
rect -6247 10239 -6189 10273
rect -6247 10205 -6235 10239
rect -6201 10205 -6189 10239
rect -6247 10164 -6189 10205
rect -5989 11123 -5931 11164
rect -5989 11089 -5977 11123
rect -5943 11089 -5931 11123
rect -5989 11055 -5931 11089
rect -5989 11021 -5977 11055
rect -5943 11021 -5931 11055
rect -5989 10987 -5931 11021
rect -5989 10953 -5977 10987
rect -5943 10953 -5931 10987
rect -5989 10919 -5931 10953
rect -5989 10885 -5977 10919
rect -5943 10885 -5931 10919
rect -5989 10851 -5931 10885
rect -5989 10817 -5977 10851
rect -5943 10817 -5931 10851
rect -5989 10783 -5931 10817
rect -5989 10749 -5977 10783
rect -5943 10749 -5931 10783
rect -5989 10715 -5931 10749
rect -5989 10681 -5977 10715
rect -5943 10681 -5931 10715
rect -5989 10647 -5931 10681
rect -5989 10613 -5977 10647
rect -5943 10613 -5931 10647
rect -5989 10579 -5931 10613
rect -5989 10545 -5977 10579
rect -5943 10545 -5931 10579
rect -5989 10511 -5931 10545
rect -5989 10477 -5977 10511
rect -5943 10477 -5931 10511
rect -5989 10443 -5931 10477
rect -5989 10409 -5977 10443
rect -5943 10409 -5931 10443
rect -5989 10375 -5931 10409
rect -5989 10341 -5977 10375
rect -5943 10341 -5931 10375
rect -5989 10307 -5931 10341
rect -5989 10273 -5977 10307
rect -5943 10273 -5931 10307
rect -5989 10239 -5931 10273
rect -5989 10205 -5977 10239
rect -5943 10205 -5931 10239
rect -5989 10164 -5931 10205
rect -5731 11123 -5673 11164
rect -5731 11089 -5719 11123
rect -5685 11089 -5673 11123
rect -5731 11055 -5673 11089
rect -5731 11021 -5719 11055
rect -5685 11021 -5673 11055
rect -5731 10987 -5673 11021
rect -5731 10953 -5719 10987
rect -5685 10953 -5673 10987
rect -5731 10919 -5673 10953
rect -5731 10885 -5719 10919
rect -5685 10885 -5673 10919
rect -5731 10851 -5673 10885
rect -5731 10817 -5719 10851
rect -5685 10817 -5673 10851
rect -5731 10783 -5673 10817
rect -5731 10749 -5719 10783
rect -5685 10749 -5673 10783
rect -5731 10715 -5673 10749
rect -5731 10681 -5719 10715
rect -5685 10681 -5673 10715
rect -5731 10647 -5673 10681
rect -5731 10613 -5719 10647
rect -5685 10613 -5673 10647
rect -5731 10579 -5673 10613
rect -5731 10545 -5719 10579
rect -5685 10545 -5673 10579
rect -5731 10511 -5673 10545
rect -5731 10477 -5719 10511
rect -5685 10477 -5673 10511
rect -5731 10443 -5673 10477
rect -5731 10409 -5719 10443
rect -5685 10409 -5673 10443
rect -5731 10375 -5673 10409
rect -5731 10341 -5719 10375
rect -5685 10341 -5673 10375
rect -5731 10307 -5673 10341
rect -5731 10273 -5719 10307
rect -5685 10273 -5673 10307
rect -5731 10239 -5673 10273
rect -5731 10205 -5719 10239
rect -5685 10205 -5673 10239
rect -5731 10164 -5673 10205
rect -5473 11123 -5415 11164
rect -5473 11089 -5461 11123
rect -5427 11089 -5415 11123
rect -5473 11055 -5415 11089
rect -5473 11021 -5461 11055
rect -5427 11021 -5415 11055
rect -5473 10987 -5415 11021
rect -5473 10953 -5461 10987
rect -5427 10953 -5415 10987
rect -5473 10919 -5415 10953
rect -5473 10885 -5461 10919
rect -5427 10885 -5415 10919
rect -5473 10851 -5415 10885
rect -5473 10817 -5461 10851
rect -5427 10817 -5415 10851
rect -5473 10783 -5415 10817
rect -5473 10749 -5461 10783
rect -5427 10749 -5415 10783
rect -5473 10715 -5415 10749
rect -5473 10681 -5461 10715
rect -5427 10681 -5415 10715
rect -5473 10647 -5415 10681
rect -5473 10613 -5461 10647
rect -5427 10613 -5415 10647
rect -5473 10579 -5415 10613
rect -5473 10545 -5461 10579
rect -5427 10545 -5415 10579
rect -5473 10511 -5415 10545
rect -5473 10477 -5461 10511
rect -5427 10477 -5415 10511
rect -5473 10443 -5415 10477
rect -5473 10409 -5461 10443
rect -5427 10409 -5415 10443
rect -5473 10375 -5415 10409
rect -5473 10341 -5461 10375
rect -5427 10341 -5415 10375
rect -5473 10307 -5415 10341
rect -5473 10273 -5461 10307
rect -5427 10273 -5415 10307
rect -5473 10239 -5415 10273
rect -5473 10205 -5461 10239
rect -5427 10205 -5415 10239
rect -5473 10164 -5415 10205
rect -5215 11123 -5157 11164
rect -5215 11089 -5203 11123
rect -5169 11089 -5157 11123
rect -5215 11055 -5157 11089
rect -5215 11021 -5203 11055
rect -5169 11021 -5157 11055
rect -5215 10987 -5157 11021
rect -5215 10953 -5203 10987
rect -5169 10953 -5157 10987
rect -5215 10919 -5157 10953
rect -5215 10885 -5203 10919
rect -5169 10885 -5157 10919
rect -5215 10851 -5157 10885
rect -5215 10817 -5203 10851
rect -5169 10817 -5157 10851
rect -5215 10783 -5157 10817
rect -5215 10749 -5203 10783
rect -5169 10749 -5157 10783
rect -5215 10715 -5157 10749
rect -5215 10681 -5203 10715
rect -5169 10681 -5157 10715
rect -5215 10647 -5157 10681
rect -5215 10613 -5203 10647
rect -5169 10613 -5157 10647
rect -5215 10579 -5157 10613
rect -5215 10545 -5203 10579
rect -5169 10545 -5157 10579
rect -5215 10511 -5157 10545
rect -5215 10477 -5203 10511
rect -5169 10477 -5157 10511
rect -5215 10443 -5157 10477
rect -5215 10409 -5203 10443
rect -5169 10409 -5157 10443
rect -5215 10375 -5157 10409
rect -5215 10341 -5203 10375
rect -5169 10341 -5157 10375
rect -5215 10307 -5157 10341
rect -5215 10273 -5203 10307
rect -5169 10273 -5157 10307
rect -5215 10239 -5157 10273
rect -5215 10205 -5203 10239
rect -5169 10205 -5157 10239
rect -5215 10164 -5157 10205
rect -4957 11123 -4899 11164
rect -4957 11089 -4945 11123
rect -4911 11089 -4899 11123
rect -4957 11055 -4899 11089
rect -4957 11021 -4945 11055
rect -4911 11021 -4899 11055
rect -4957 10987 -4899 11021
rect -4957 10953 -4945 10987
rect -4911 10953 -4899 10987
rect -4957 10919 -4899 10953
rect -4957 10885 -4945 10919
rect -4911 10885 -4899 10919
rect -4957 10851 -4899 10885
rect -4957 10817 -4945 10851
rect -4911 10817 -4899 10851
rect -4957 10783 -4899 10817
rect -4957 10749 -4945 10783
rect -4911 10749 -4899 10783
rect -4957 10715 -4899 10749
rect -4957 10681 -4945 10715
rect -4911 10681 -4899 10715
rect -4957 10647 -4899 10681
rect -4957 10613 -4945 10647
rect -4911 10613 -4899 10647
rect -4957 10579 -4899 10613
rect -4957 10545 -4945 10579
rect -4911 10545 -4899 10579
rect -4957 10511 -4899 10545
rect -4957 10477 -4945 10511
rect -4911 10477 -4899 10511
rect -4957 10443 -4899 10477
rect -4957 10409 -4945 10443
rect -4911 10409 -4899 10443
rect -4957 10375 -4899 10409
rect -4957 10341 -4945 10375
rect -4911 10341 -4899 10375
rect -4957 10307 -4899 10341
rect -4957 10273 -4945 10307
rect -4911 10273 -4899 10307
rect -4957 10239 -4899 10273
rect -4957 10205 -4945 10239
rect -4911 10205 -4899 10239
rect -4957 10164 -4899 10205
rect -4699 11123 -4641 11164
rect -4699 11089 -4687 11123
rect -4653 11089 -4641 11123
rect -4699 11055 -4641 11089
rect -4699 11021 -4687 11055
rect -4653 11021 -4641 11055
rect -4699 10987 -4641 11021
rect -4699 10953 -4687 10987
rect -4653 10953 -4641 10987
rect -4699 10919 -4641 10953
rect -4699 10885 -4687 10919
rect -4653 10885 -4641 10919
rect -4699 10851 -4641 10885
rect -4699 10817 -4687 10851
rect -4653 10817 -4641 10851
rect -4699 10783 -4641 10817
rect -4699 10749 -4687 10783
rect -4653 10749 -4641 10783
rect -4699 10715 -4641 10749
rect -4699 10681 -4687 10715
rect -4653 10681 -4641 10715
rect -4699 10647 -4641 10681
rect -4699 10613 -4687 10647
rect -4653 10613 -4641 10647
rect -4699 10579 -4641 10613
rect -4699 10545 -4687 10579
rect -4653 10545 -4641 10579
rect -4699 10511 -4641 10545
rect -4699 10477 -4687 10511
rect -4653 10477 -4641 10511
rect -4699 10443 -4641 10477
rect -4699 10409 -4687 10443
rect -4653 10409 -4641 10443
rect -4699 10375 -4641 10409
rect -4699 10341 -4687 10375
rect -4653 10341 -4641 10375
rect -4699 10307 -4641 10341
rect -4699 10273 -4687 10307
rect -4653 10273 -4641 10307
rect -4699 10239 -4641 10273
rect -4699 10205 -4687 10239
rect -4653 10205 -4641 10239
rect -4699 10164 -4641 10205
rect -4441 11123 -4383 11164
rect -4441 11089 -4429 11123
rect -4395 11089 -4383 11123
rect -4441 11055 -4383 11089
rect -4441 11021 -4429 11055
rect -4395 11021 -4383 11055
rect -4441 10987 -4383 11021
rect -4441 10953 -4429 10987
rect -4395 10953 -4383 10987
rect -4441 10919 -4383 10953
rect -4441 10885 -4429 10919
rect -4395 10885 -4383 10919
rect -4441 10851 -4383 10885
rect -4441 10817 -4429 10851
rect -4395 10817 -4383 10851
rect -4441 10783 -4383 10817
rect -4441 10749 -4429 10783
rect -4395 10749 -4383 10783
rect -4441 10715 -4383 10749
rect -4441 10681 -4429 10715
rect -4395 10681 -4383 10715
rect -4441 10647 -4383 10681
rect -4441 10613 -4429 10647
rect -4395 10613 -4383 10647
rect -4441 10579 -4383 10613
rect -4441 10545 -4429 10579
rect -4395 10545 -4383 10579
rect -4441 10511 -4383 10545
rect -4441 10477 -4429 10511
rect -4395 10477 -4383 10511
rect -4441 10443 -4383 10477
rect -4441 10409 -4429 10443
rect -4395 10409 -4383 10443
rect -4441 10375 -4383 10409
rect -4441 10341 -4429 10375
rect -4395 10341 -4383 10375
rect -4441 10307 -4383 10341
rect -4441 10273 -4429 10307
rect -4395 10273 -4383 10307
rect -4441 10239 -4383 10273
rect -4441 10205 -4429 10239
rect -4395 10205 -4383 10239
rect -4441 10164 -4383 10205
rect -4183 11123 -4125 11164
rect -4183 11089 -4171 11123
rect -4137 11089 -4125 11123
rect -4183 11055 -4125 11089
rect -4183 11021 -4171 11055
rect -4137 11021 -4125 11055
rect -4183 10987 -4125 11021
rect -4183 10953 -4171 10987
rect -4137 10953 -4125 10987
rect -4183 10919 -4125 10953
rect -4183 10885 -4171 10919
rect -4137 10885 -4125 10919
rect -4183 10851 -4125 10885
rect -4183 10817 -4171 10851
rect -4137 10817 -4125 10851
rect -4183 10783 -4125 10817
rect -4183 10749 -4171 10783
rect -4137 10749 -4125 10783
rect -4183 10715 -4125 10749
rect -4183 10681 -4171 10715
rect -4137 10681 -4125 10715
rect -4183 10647 -4125 10681
rect -4183 10613 -4171 10647
rect -4137 10613 -4125 10647
rect -4183 10579 -4125 10613
rect -4183 10545 -4171 10579
rect -4137 10545 -4125 10579
rect -4183 10511 -4125 10545
rect -4183 10477 -4171 10511
rect -4137 10477 -4125 10511
rect -4183 10443 -4125 10477
rect -4183 10409 -4171 10443
rect -4137 10409 -4125 10443
rect -4183 10375 -4125 10409
rect -4183 10341 -4171 10375
rect -4137 10341 -4125 10375
rect -4183 10307 -4125 10341
rect -4183 10273 -4171 10307
rect -4137 10273 -4125 10307
rect -4183 10239 -4125 10273
rect -4183 10205 -4171 10239
rect -4137 10205 -4125 10239
rect -4183 10164 -4125 10205
rect -3925 11123 -3867 11164
rect -3925 11089 -3913 11123
rect -3879 11089 -3867 11123
rect -3925 11055 -3867 11089
rect -3925 11021 -3913 11055
rect -3879 11021 -3867 11055
rect -3925 10987 -3867 11021
rect -3925 10953 -3913 10987
rect -3879 10953 -3867 10987
rect -3925 10919 -3867 10953
rect -3925 10885 -3913 10919
rect -3879 10885 -3867 10919
rect -3925 10851 -3867 10885
rect -3925 10817 -3913 10851
rect -3879 10817 -3867 10851
rect -3925 10783 -3867 10817
rect -3925 10749 -3913 10783
rect -3879 10749 -3867 10783
rect -3925 10715 -3867 10749
rect -3925 10681 -3913 10715
rect -3879 10681 -3867 10715
rect -3925 10647 -3867 10681
rect -3925 10613 -3913 10647
rect -3879 10613 -3867 10647
rect -3925 10579 -3867 10613
rect -3925 10545 -3913 10579
rect -3879 10545 -3867 10579
rect -3925 10511 -3867 10545
rect -3925 10477 -3913 10511
rect -3879 10477 -3867 10511
rect -3925 10443 -3867 10477
rect -3925 10409 -3913 10443
rect -3879 10409 -3867 10443
rect -3925 10375 -3867 10409
rect -3925 10341 -3913 10375
rect -3879 10341 -3867 10375
rect -3925 10307 -3867 10341
rect -3925 10273 -3913 10307
rect -3879 10273 -3867 10307
rect -3925 10239 -3867 10273
rect -3925 10205 -3913 10239
rect -3879 10205 -3867 10239
rect -3925 10164 -3867 10205
rect -3667 11123 -3609 11164
rect -3667 11089 -3655 11123
rect -3621 11089 -3609 11123
rect -3667 11055 -3609 11089
rect -3667 11021 -3655 11055
rect -3621 11021 -3609 11055
rect -3667 10987 -3609 11021
rect -3667 10953 -3655 10987
rect -3621 10953 -3609 10987
rect -3667 10919 -3609 10953
rect -3667 10885 -3655 10919
rect -3621 10885 -3609 10919
rect -3667 10851 -3609 10885
rect -3667 10817 -3655 10851
rect -3621 10817 -3609 10851
rect -3667 10783 -3609 10817
rect -3667 10749 -3655 10783
rect -3621 10749 -3609 10783
rect -3667 10715 -3609 10749
rect -3667 10681 -3655 10715
rect -3621 10681 -3609 10715
rect -3667 10647 -3609 10681
rect -3667 10613 -3655 10647
rect -3621 10613 -3609 10647
rect -3667 10579 -3609 10613
rect -3667 10545 -3655 10579
rect -3621 10545 -3609 10579
rect -3667 10511 -3609 10545
rect -3667 10477 -3655 10511
rect -3621 10477 -3609 10511
rect -3667 10443 -3609 10477
rect -3667 10409 -3655 10443
rect -3621 10409 -3609 10443
rect -3667 10375 -3609 10409
rect -3667 10341 -3655 10375
rect -3621 10341 -3609 10375
rect -3667 10307 -3609 10341
rect -3667 10273 -3655 10307
rect -3621 10273 -3609 10307
rect -3667 10239 -3609 10273
rect -3667 10205 -3655 10239
rect -3621 10205 -3609 10239
rect -3667 10164 -3609 10205
rect -7792 9758 -7734 9799
rect -7792 9724 -7780 9758
rect -7746 9724 -7734 9758
rect -7792 9690 -7734 9724
rect -7792 9656 -7780 9690
rect -7746 9656 -7734 9690
rect -7792 9622 -7734 9656
rect -7792 9588 -7780 9622
rect -7746 9588 -7734 9622
rect -7792 9554 -7734 9588
rect -7792 9520 -7780 9554
rect -7746 9520 -7734 9554
rect -7792 9486 -7734 9520
rect -7792 9452 -7780 9486
rect -7746 9452 -7734 9486
rect -7792 9418 -7734 9452
rect -7792 9384 -7780 9418
rect -7746 9384 -7734 9418
rect -7792 9350 -7734 9384
rect -7792 9316 -7780 9350
rect -7746 9316 -7734 9350
rect -7792 9282 -7734 9316
rect -7792 9248 -7780 9282
rect -7746 9248 -7734 9282
rect -7792 9214 -7734 9248
rect -7792 9180 -7780 9214
rect -7746 9180 -7734 9214
rect -7792 9146 -7734 9180
rect -7792 9112 -7780 9146
rect -7746 9112 -7734 9146
rect -7792 9078 -7734 9112
rect -7792 9044 -7780 9078
rect -7746 9044 -7734 9078
rect -7792 9010 -7734 9044
rect -7792 8976 -7780 9010
rect -7746 8976 -7734 9010
rect -7792 8942 -7734 8976
rect -7792 8908 -7780 8942
rect -7746 8908 -7734 8942
rect -7792 8874 -7734 8908
rect -7792 8840 -7780 8874
rect -7746 8840 -7734 8874
rect -7792 8799 -7734 8840
rect -7534 9758 -7476 9799
rect -7534 9724 -7522 9758
rect -7488 9724 -7476 9758
rect -7534 9690 -7476 9724
rect -7534 9656 -7522 9690
rect -7488 9656 -7476 9690
rect -7534 9622 -7476 9656
rect -7534 9588 -7522 9622
rect -7488 9588 -7476 9622
rect -7534 9554 -7476 9588
rect -7534 9520 -7522 9554
rect -7488 9520 -7476 9554
rect -7534 9486 -7476 9520
rect -7534 9452 -7522 9486
rect -7488 9452 -7476 9486
rect -7534 9418 -7476 9452
rect -7534 9384 -7522 9418
rect -7488 9384 -7476 9418
rect -7534 9350 -7476 9384
rect -7534 9316 -7522 9350
rect -7488 9316 -7476 9350
rect -7534 9282 -7476 9316
rect -7534 9248 -7522 9282
rect -7488 9248 -7476 9282
rect -7534 9214 -7476 9248
rect -7534 9180 -7522 9214
rect -7488 9180 -7476 9214
rect -7534 9146 -7476 9180
rect -7534 9112 -7522 9146
rect -7488 9112 -7476 9146
rect -7534 9078 -7476 9112
rect -7534 9044 -7522 9078
rect -7488 9044 -7476 9078
rect -7534 9010 -7476 9044
rect -7534 8976 -7522 9010
rect -7488 8976 -7476 9010
rect -7534 8942 -7476 8976
rect -7534 8908 -7522 8942
rect -7488 8908 -7476 8942
rect -7534 8874 -7476 8908
rect -7534 8840 -7522 8874
rect -7488 8840 -7476 8874
rect -7534 8799 -7476 8840
rect -7326 9758 -7268 9799
rect -7326 9724 -7314 9758
rect -7280 9724 -7268 9758
rect -7326 9690 -7268 9724
rect -7326 9656 -7314 9690
rect -7280 9656 -7268 9690
rect -7326 9622 -7268 9656
rect -7326 9588 -7314 9622
rect -7280 9588 -7268 9622
rect -7326 9554 -7268 9588
rect -7326 9520 -7314 9554
rect -7280 9520 -7268 9554
rect -7326 9486 -7268 9520
rect -7326 9452 -7314 9486
rect -7280 9452 -7268 9486
rect -7326 9418 -7268 9452
rect -7326 9384 -7314 9418
rect -7280 9384 -7268 9418
rect -7326 9350 -7268 9384
rect -7326 9316 -7314 9350
rect -7280 9316 -7268 9350
rect -7326 9282 -7268 9316
rect -7326 9248 -7314 9282
rect -7280 9248 -7268 9282
rect -7326 9214 -7268 9248
rect -7326 9180 -7314 9214
rect -7280 9180 -7268 9214
rect -7326 9146 -7268 9180
rect -7326 9112 -7314 9146
rect -7280 9112 -7268 9146
rect -7326 9078 -7268 9112
rect -7326 9044 -7314 9078
rect -7280 9044 -7268 9078
rect -7326 9010 -7268 9044
rect -7326 8976 -7314 9010
rect -7280 8976 -7268 9010
rect -7326 8942 -7268 8976
rect -7326 8908 -7314 8942
rect -7280 8908 -7268 8942
rect -7326 8874 -7268 8908
rect -7326 8840 -7314 8874
rect -7280 8840 -7268 8874
rect -7326 8799 -7268 8840
rect -7068 9758 -7010 9799
rect -7068 9724 -7056 9758
rect -7022 9724 -7010 9758
rect -7068 9690 -7010 9724
rect -7068 9656 -7056 9690
rect -7022 9656 -7010 9690
rect -7068 9622 -7010 9656
rect -7068 9588 -7056 9622
rect -7022 9588 -7010 9622
rect -7068 9554 -7010 9588
rect -7068 9520 -7056 9554
rect -7022 9520 -7010 9554
rect -7068 9486 -7010 9520
rect -7068 9452 -7056 9486
rect -7022 9452 -7010 9486
rect -7068 9418 -7010 9452
rect -7068 9384 -7056 9418
rect -7022 9384 -7010 9418
rect -7068 9350 -7010 9384
rect -7068 9316 -7056 9350
rect -7022 9316 -7010 9350
rect -7068 9282 -7010 9316
rect -7068 9248 -7056 9282
rect -7022 9248 -7010 9282
rect -7068 9214 -7010 9248
rect -7068 9180 -7056 9214
rect -7022 9180 -7010 9214
rect -7068 9146 -7010 9180
rect -7068 9112 -7056 9146
rect -7022 9112 -7010 9146
rect -7068 9078 -7010 9112
rect -7068 9044 -7056 9078
rect -7022 9044 -7010 9078
rect -7068 9010 -7010 9044
rect -7068 8976 -7056 9010
rect -7022 8976 -7010 9010
rect -7068 8942 -7010 8976
rect -7068 8908 -7056 8942
rect -7022 8908 -7010 8942
rect -7068 8874 -7010 8908
rect -7068 8840 -7056 8874
rect -7022 8840 -7010 8874
rect -7068 8799 -7010 8840
rect -6810 9758 -6752 9799
rect -6810 9724 -6798 9758
rect -6764 9724 -6752 9758
rect -6810 9690 -6752 9724
rect -6810 9656 -6798 9690
rect -6764 9656 -6752 9690
rect -6810 9622 -6752 9656
rect -6810 9588 -6798 9622
rect -6764 9588 -6752 9622
rect -6810 9554 -6752 9588
rect -6810 9520 -6798 9554
rect -6764 9520 -6752 9554
rect -6810 9486 -6752 9520
rect -6810 9452 -6798 9486
rect -6764 9452 -6752 9486
rect -6810 9418 -6752 9452
rect -6810 9384 -6798 9418
rect -6764 9384 -6752 9418
rect -6810 9350 -6752 9384
rect -6810 9316 -6798 9350
rect -6764 9316 -6752 9350
rect -6810 9282 -6752 9316
rect -6810 9248 -6798 9282
rect -6764 9248 -6752 9282
rect -6810 9214 -6752 9248
rect -6810 9180 -6798 9214
rect -6764 9180 -6752 9214
rect -6810 9146 -6752 9180
rect -6810 9112 -6798 9146
rect -6764 9112 -6752 9146
rect -6810 9078 -6752 9112
rect -6810 9044 -6798 9078
rect -6764 9044 -6752 9078
rect -6810 9010 -6752 9044
rect -6810 8976 -6798 9010
rect -6764 8976 -6752 9010
rect -6810 8942 -6752 8976
rect -6810 8908 -6798 8942
rect -6764 8908 -6752 8942
rect -6810 8874 -6752 8908
rect -6810 8840 -6798 8874
rect -6764 8840 -6752 8874
rect -6810 8799 -6752 8840
rect -6552 9758 -6494 9799
rect -6552 9724 -6540 9758
rect -6506 9724 -6494 9758
rect -6552 9690 -6494 9724
rect -6552 9656 -6540 9690
rect -6506 9656 -6494 9690
rect -6552 9622 -6494 9656
rect -6552 9588 -6540 9622
rect -6506 9588 -6494 9622
rect -6552 9554 -6494 9588
rect -6552 9520 -6540 9554
rect -6506 9520 -6494 9554
rect -6552 9486 -6494 9520
rect -6552 9452 -6540 9486
rect -6506 9452 -6494 9486
rect -6552 9418 -6494 9452
rect -6552 9384 -6540 9418
rect -6506 9384 -6494 9418
rect -6552 9350 -6494 9384
rect -6552 9316 -6540 9350
rect -6506 9316 -6494 9350
rect -6552 9282 -6494 9316
rect -6552 9248 -6540 9282
rect -6506 9248 -6494 9282
rect -6552 9214 -6494 9248
rect -6552 9180 -6540 9214
rect -6506 9180 -6494 9214
rect -6552 9146 -6494 9180
rect -6552 9112 -6540 9146
rect -6506 9112 -6494 9146
rect -6552 9078 -6494 9112
rect -6552 9044 -6540 9078
rect -6506 9044 -6494 9078
rect -6552 9010 -6494 9044
rect -6552 8976 -6540 9010
rect -6506 8976 -6494 9010
rect -6552 8942 -6494 8976
rect -6552 8908 -6540 8942
rect -6506 8908 -6494 8942
rect -6552 8874 -6494 8908
rect -6552 8840 -6540 8874
rect -6506 8840 -6494 8874
rect -6552 8799 -6494 8840
rect -6294 9758 -6236 9799
rect -6294 9724 -6282 9758
rect -6248 9724 -6236 9758
rect -6294 9690 -6236 9724
rect -6294 9656 -6282 9690
rect -6248 9656 -6236 9690
rect -6294 9622 -6236 9656
rect -6294 9588 -6282 9622
rect -6248 9588 -6236 9622
rect -6294 9554 -6236 9588
rect -6294 9520 -6282 9554
rect -6248 9520 -6236 9554
rect -6294 9486 -6236 9520
rect -6294 9452 -6282 9486
rect -6248 9452 -6236 9486
rect -6294 9418 -6236 9452
rect -6294 9384 -6282 9418
rect -6248 9384 -6236 9418
rect -6294 9350 -6236 9384
rect -6294 9316 -6282 9350
rect -6248 9316 -6236 9350
rect -6294 9282 -6236 9316
rect -6294 9248 -6282 9282
rect -6248 9248 -6236 9282
rect -6294 9214 -6236 9248
rect -6294 9180 -6282 9214
rect -6248 9180 -6236 9214
rect -6294 9146 -6236 9180
rect -6294 9112 -6282 9146
rect -6248 9112 -6236 9146
rect -6294 9078 -6236 9112
rect -6294 9044 -6282 9078
rect -6248 9044 -6236 9078
rect -6294 9010 -6236 9044
rect -6294 8976 -6282 9010
rect -6248 8976 -6236 9010
rect -6294 8942 -6236 8976
rect -6294 8908 -6282 8942
rect -6248 8908 -6236 8942
rect -6294 8874 -6236 8908
rect -6294 8840 -6282 8874
rect -6248 8840 -6236 8874
rect -6294 8799 -6236 8840
rect -6036 9758 -5978 9799
rect -6036 9724 -6024 9758
rect -5990 9724 -5978 9758
rect -6036 9690 -5978 9724
rect -6036 9656 -6024 9690
rect -5990 9656 -5978 9690
rect -6036 9622 -5978 9656
rect -6036 9588 -6024 9622
rect -5990 9588 -5978 9622
rect -6036 9554 -5978 9588
rect -6036 9520 -6024 9554
rect -5990 9520 -5978 9554
rect -6036 9486 -5978 9520
rect -6036 9452 -6024 9486
rect -5990 9452 -5978 9486
rect -6036 9418 -5978 9452
rect -6036 9384 -6024 9418
rect -5990 9384 -5978 9418
rect -6036 9350 -5978 9384
rect -6036 9316 -6024 9350
rect -5990 9316 -5978 9350
rect -6036 9282 -5978 9316
rect -6036 9248 -6024 9282
rect -5990 9248 -5978 9282
rect -6036 9214 -5978 9248
rect -6036 9180 -6024 9214
rect -5990 9180 -5978 9214
rect -6036 9146 -5978 9180
rect -6036 9112 -6024 9146
rect -5990 9112 -5978 9146
rect -6036 9078 -5978 9112
rect -6036 9044 -6024 9078
rect -5990 9044 -5978 9078
rect -6036 9010 -5978 9044
rect -6036 8976 -6024 9010
rect -5990 8976 -5978 9010
rect -6036 8942 -5978 8976
rect -6036 8908 -6024 8942
rect -5990 8908 -5978 8942
rect -6036 8874 -5978 8908
rect -6036 8840 -6024 8874
rect -5990 8840 -5978 8874
rect -6036 8799 -5978 8840
rect -5778 9758 -5720 9799
rect -5778 9724 -5766 9758
rect -5732 9724 -5720 9758
rect -5778 9690 -5720 9724
rect -5778 9656 -5766 9690
rect -5732 9656 -5720 9690
rect -5778 9622 -5720 9656
rect -5778 9588 -5766 9622
rect -5732 9588 -5720 9622
rect -5778 9554 -5720 9588
rect -5778 9520 -5766 9554
rect -5732 9520 -5720 9554
rect -5778 9486 -5720 9520
rect -5778 9452 -5766 9486
rect -5732 9452 -5720 9486
rect -5778 9418 -5720 9452
rect -5778 9384 -5766 9418
rect -5732 9384 -5720 9418
rect -5778 9350 -5720 9384
rect -5778 9316 -5766 9350
rect -5732 9316 -5720 9350
rect -5778 9282 -5720 9316
rect -5778 9248 -5766 9282
rect -5732 9248 -5720 9282
rect -5778 9214 -5720 9248
rect -5778 9180 -5766 9214
rect -5732 9180 -5720 9214
rect -5778 9146 -5720 9180
rect -5778 9112 -5766 9146
rect -5732 9112 -5720 9146
rect -5778 9078 -5720 9112
rect -5778 9044 -5766 9078
rect -5732 9044 -5720 9078
rect -5778 9010 -5720 9044
rect -5778 8976 -5766 9010
rect -5732 8976 -5720 9010
rect -5778 8942 -5720 8976
rect -5778 8908 -5766 8942
rect -5732 8908 -5720 8942
rect -5778 8874 -5720 8908
rect -5778 8840 -5766 8874
rect -5732 8840 -5720 8874
rect -5778 8799 -5720 8840
rect -5520 9758 -5462 9799
rect -5520 9724 -5508 9758
rect -5474 9724 -5462 9758
rect -5520 9690 -5462 9724
rect -5520 9656 -5508 9690
rect -5474 9656 -5462 9690
rect -5520 9622 -5462 9656
rect -5520 9588 -5508 9622
rect -5474 9588 -5462 9622
rect -5520 9554 -5462 9588
rect -5520 9520 -5508 9554
rect -5474 9520 -5462 9554
rect -5520 9486 -5462 9520
rect -5520 9452 -5508 9486
rect -5474 9452 -5462 9486
rect -5520 9418 -5462 9452
rect -5520 9384 -5508 9418
rect -5474 9384 -5462 9418
rect -5520 9350 -5462 9384
rect -5520 9316 -5508 9350
rect -5474 9316 -5462 9350
rect -5520 9282 -5462 9316
rect -5520 9248 -5508 9282
rect -5474 9248 -5462 9282
rect -5520 9214 -5462 9248
rect -5520 9180 -5508 9214
rect -5474 9180 -5462 9214
rect -5520 9146 -5462 9180
rect -5520 9112 -5508 9146
rect -5474 9112 -5462 9146
rect -5520 9078 -5462 9112
rect -5520 9044 -5508 9078
rect -5474 9044 -5462 9078
rect -5520 9010 -5462 9044
rect -5520 8976 -5508 9010
rect -5474 8976 -5462 9010
rect -5520 8942 -5462 8976
rect -5520 8908 -5508 8942
rect -5474 8908 -5462 8942
rect -5520 8874 -5462 8908
rect -5520 8840 -5508 8874
rect -5474 8840 -5462 8874
rect -5520 8799 -5462 8840
rect -5262 9758 -5204 9799
rect -5262 9724 -5250 9758
rect -5216 9724 -5204 9758
rect -5262 9690 -5204 9724
rect -5262 9656 -5250 9690
rect -5216 9656 -5204 9690
rect -5262 9622 -5204 9656
rect -5262 9588 -5250 9622
rect -5216 9588 -5204 9622
rect -5262 9554 -5204 9588
rect -5262 9520 -5250 9554
rect -5216 9520 -5204 9554
rect -5262 9486 -5204 9520
rect -5262 9452 -5250 9486
rect -5216 9452 -5204 9486
rect -5262 9418 -5204 9452
rect -5262 9384 -5250 9418
rect -5216 9384 -5204 9418
rect -5262 9350 -5204 9384
rect -5262 9316 -5250 9350
rect -5216 9316 -5204 9350
rect -5262 9282 -5204 9316
rect -5262 9248 -5250 9282
rect -5216 9248 -5204 9282
rect -5262 9214 -5204 9248
rect -5262 9180 -5250 9214
rect -5216 9180 -5204 9214
rect -5262 9146 -5204 9180
rect -5262 9112 -5250 9146
rect -5216 9112 -5204 9146
rect -5262 9078 -5204 9112
rect -5262 9044 -5250 9078
rect -5216 9044 -5204 9078
rect -5262 9010 -5204 9044
rect -5262 8976 -5250 9010
rect -5216 8976 -5204 9010
rect -5262 8942 -5204 8976
rect -5262 8908 -5250 8942
rect -5216 8908 -5204 8942
rect -5262 8874 -5204 8908
rect -5262 8840 -5250 8874
rect -5216 8840 -5204 8874
rect -5262 8799 -5204 8840
rect -5004 9758 -4946 9799
rect -5004 9724 -4992 9758
rect -4958 9724 -4946 9758
rect -5004 9690 -4946 9724
rect -5004 9656 -4992 9690
rect -4958 9656 -4946 9690
rect -5004 9622 -4946 9656
rect -5004 9588 -4992 9622
rect -4958 9588 -4946 9622
rect -5004 9554 -4946 9588
rect -5004 9520 -4992 9554
rect -4958 9520 -4946 9554
rect -5004 9486 -4946 9520
rect -5004 9452 -4992 9486
rect -4958 9452 -4946 9486
rect -5004 9418 -4946 9452
rect -5004 9384 -4992 9418
rect -4958 9384 -4946 9418
rect -5004 9350 -4946 9384
rect -5004 9316 -4992 9350
rect -4958 9316 -4946 9350
rect -5004 9282 -4946 9316
rect -5004 9248 -4992 9282
rect -4958 9248 -4946 9282
rect -5004 9214 -4946 9248
rect -5004 9180 -4992 9214
rect -4958 9180 -4946 9214
rect -5004 9146 -4946 9180
rect -5004 9112 -4992 9146
rect -4958 9112 -4946 9146
rect -5004 9078 -4946 9112
rect -5004 9044 -4992 9078
rect -4958 9044 -4946 9078
rect -5004 9010 -4946 9044
rect -5004 8976 -4992 9010
rect -4958 8976 -4946 9010
rect -5004 8942 -4946 8976
rect -5004 8908 -4992 8942
rect -4958 8908 -4946 8942
rect -5004 8874 -4946 8908
rect -5004 8840 -4992 8874
rect -4958 8840 -4946 8874
rect -5004 8799 -4946 8840
rect -4746 9758 -4688 9799
rect -4746 9724 -4734 9758
rect -4700 9724 -4688 9758
rect -4746 9690 -4688 9724
rect -4746 9656 -4734 9690
rect -4700 9656 -4688 9690
rect -4746 9622 -4688 9656
rect -4746 9588 -4734 9622
rect -4700 9588 -4688 9622
rect -4746 9554 -4688 9588
rect -4746 9520 -4734 9554
rect -4700 9520 -4688 9554
rect -4746 9486 -4688 9520
rect -4746 9452 -4734 9486
rect -4700 9452 -4688 9486
rect -4746 9418 -4688 9452
rect -4746 9384 -4734 9418
rect -4700 9384 -4688 9418
rect -4746 9350 -4688 9384
rect -4746 9316 -4734 9350
rect -4700 9316 -4688 9350
rect -4746 9282 -4688 9316
rect -4746 9248 -4734 9282
rect -4700 9248 -4688 9282
rect -4746 9214 -4688 9248
rect -4746 9180 -4734 9214
rect -4700 9180 -4688 9214
rect -4746 9146 -4688 9180
rect -4746 9112 -4734 9146
rect -4700 9112 -4688 9146
rect -4746 9078 -4688 9112
rect -4746 9044 -4734 9078
rect -4700 9044 -4688 9078
rect -4746 9010 -4688 9044
rect -4746 8976 -4734 9010
rect -4700 8976 -4688 9010
rect -4746 8942 -4688 8976
rect -4746 8908 -4734 8942
rect -4700 8908 -4688 8942
rect -4746 8874 -4688 8908
rect -4746 8840 -4734 8874
rect -4700 8840 -4688 8874
rect -4746 8799 -4688 8840
rect -7792 7507 -7734 7538
rect -7792 7473 -7780 7507
rect -7746 7473 -7734 7507
rect -7792 7439 -7734 7473
rect -7792 7405 -7780 7439
rect -7746 7405 -7734 7439
rect -7792 7371 -7734 7405
rect -7792 7337 -7780 7371
rect -7746 7337 -7734 7371
rect -7792 7303 -7734 7337
rect -7792 7269 -7780 7303
rect -7746 7269 -7734 7303
rect -7792 7235 -7734 7269
rect -7792 7201 -7780 7235
rect -7746 7201 -7734 7235
rect -7792 7167 -7734 7201
rect -7792 7133 -7780 7167
rect -7746 7133 -7734 7167
rect -7792 7099 -7734 7133
rect -7792 7065 -7780 7099
rect -7746 7065 -7734 7099
rect -7792 7031 -7734 7065
rect -7792 6997 -7780 7031
rect -7746 6997 -7734 7031
rect -7792 6963 -7734 6997
rect -7792 6929 -7780 6963
rect -7746 6929 -7734 6963
rect -7792 6895 -7734 6929
rect -7792 6861 -7780 6895
rect -7746 6861 -7734 6895
rect -7792 6827 -7734 6861
rect -7792 6793 -7780 6827
rect -7746 6793 -7734 6827
rect -7792 6759 -7734 6793
rect -7792 6725 -7780 6759
rect -7746 6725 -7734 6759
rect -7792 6691 -7734 6725
rect -7792 6657 -7780 6691
rect -7746 6657 -7734 6691
rect -7792 6623 -7734 6657
rect -7792 6589 -7780 6623
rect -7746 6589 -7734 6623
rect -7792 6555 -7734 6589
rect -7792 6521 -7780 6555
rect -7746 6521 -7734 6555
rect -7792 6487 -7734 6521
rect -7792 6453 -7780 6487
rect -7746 6453 -7734 6487
rect -7792 6419 -7734 6453
rect -7792 6385 -7780 6419
rect -7746 6385 -7734 6419
rect -7792 6351 -7734 6385
rect -7792 6317 -7780 6351
rect -7746 6317 -7734 6351
rect -7792 6283 -7734 6317
rect -7792 6249 -7780 6283
rect -7746 6249 -7734 6283
rect -7792 6215 -7734 6249
rect -7792 6181 -7780 6215
rect -7746 6181 -7734 6215
rect -7792 6147 -7734 6181
rect -7792 6113 -7780 6147
rect -7746 6113 -7734 6147
rect -7792 6079 -7734 6113
rect -7792 6045 -7780 6079
rect -7746 6045 -7734 6079
rect -7792 6011 -7734 6045
rect -7792 5977 -7780 6011
rect -7746 5977 -7734 6011
rect -7792 5943 -7734 5977
rect -7792 5909 -7780 5943
rect -7746 5909 -7734 5943
rect -7792 5875 -7734 5909
rect -7792 5841 -7780 5875
rect -7746 5841 -7734 5875
rect -7792 5807 -7734 5841
rect -7792 5773 -7780 5807
rect -7746 5773 -7734 5807
rect -7792 5739 -7734 5773
rect -7792 5705 -7780 5739
rect -7746 5705 -7734 5739
rect -7792 5671 -7734 5705
rect -7792 5637 -7780 5671
rect -7746 5637 -7734 5671
rect -7792 5603 -7734 5637
rect -7792 5569 -7780 5603
rect -7746 5569 -7734 5603
rect -7792 5538 -7734 5569
rect -7534 7507 -7476 7538
rect -7534 7473 -7522 7507
rect -7488 7473 -7476 7507
rect -7534 7439 -7476 7473
rect -7534 7405 -7522 7439
rect -7488 7405 -7476 7439
rect -7534 7371 -7476 7405
rect -7534 7337 -7522 7371
rect -7488 7337 -7476 7371
rect -7534 7303 -7476 7337
rect -7534 7269 -7522 7303
rect -7488 7269 -7476 7303
rect -7534 7235 -7476 7269
rect -7534 7201 -7522 7235
rect -7488 7201 -7476 7235
rect -7534 7167 -7476 7201
rect -7534 7133 -7522 7167
rect -7488 7133 -7476 7167
rect -7534 7099 -7476 7133
rect -7534 7065 -7522 7099
rect -7488 7065 -7476 7099
rect -7534 7031 -7476 7065
rect -7534 6997 -7522 7031
rect -7488 6997 -7476 7031
rect -7534 6963 -7476 6997
rect -7534 6929 -7522 6963
rect -7488 6929 -7476 6963
rect -7534 6895 -7476 6929
rect -7534 6861 -7522 6895
rect -7488 6861 -7476 6895
rect -7534 6827 -7476 6861
rect -7534 6793 -7522 6827
rect -7488 6793 -7476 6827
rect -7534 6759 -7476 6793
rect -7534 6725 -7522 6759
rect -7488 6725 -7476 6759
rect -7534 6691 -7476 6725
rect -7534 6657 -7522 6691
rect -7488 6657 -7476 6691
rect -7534 6623 -7476 6657
rect -7534 6589 -7522 6623
rect -7488 6589 -7476 6623
rect -7534 6555 -7476 6589
rect -7534 6521 -7522 6555
rect -7488 6521 -7476 6555
rect -7534 6487 -7476 6521
rect -7534 6453 -7522 6487
rect -7488 6453 -7476 6487
rect -7534 6419 -7476 6453
rect -7534 6385 -7522 6419
rect -7488 6385 -7476 6419
rect -7534 6351 -7476 6385
rect -7534 6317 -7522 6351
rect -7488 6317 -7476 6351
rect -7534 6283 -7476 6317
rect -7534 6249 -7522 6283
rect -7488 6249 -7476 6283
rect -7534 6215 -7476 6249
rect -7534 6181 -7522 6215
rect -7488 6181 -7476 6215
rect -7534 6147 -7476 6181
rect -7534 6113 -7522 6147
rect -7488 6113 -7476 6147
rect -7534 6079 -7476 6113
rect -7534 6045 -7522 6079
rect -7488 6045 -7476 6079
rect -7534 6011 -7476 6045
rect -7534 5977 -7522 6011
rect -7488 5977 -7476 6011
rect -7534 5943 -7476 5977
rect -7534 5909 -7522 5943
rect -7488 5909 -7476 5943
rect -7534 5875 -7476 5909
rect -7534 5841 -7522 5875
rect -7488 5841 -7476 5875
rect -7534 5807 -7476 5841
rect -7534 5773 -7522 5807
rect -7488 5773 -7476 5807
rect -7534 5739 -7476 5773
rect -7534 5705 -7522 5739
rect -7488 5705 -7476 5739
rect -7534 5671 -7476 5705
rect -7534 5637 -7522 5671
rect -7488 5637 -7476 5671
rect -7534 5603 -7476 5637
rect -7534 5569 -7522 5603
rect -7488 5569 -7476 5603
rect -7534 5538 -7476 5569
rect -7276 7507 -7218 7538
rect -7276 7473 -7264 7507
rect -7230 7473 -7218 7507
rect -7276 7439 -7218 7473
rect -7276 7405 -7264 7439
rect -7230 7405 -7218 7439
rect -7276 7371 -7218 7405
rect -7276 7337 -7264 7371
rect -7230 7337 -7218 7371
rect -7276 7303 -7218 7337
rect -7276 7269 -7264 7303
rect -7230 7269 -7218 7303
rect -7276 7235 -7218 7269
rect -7276 7201 -7264 7235
rect -7230 7201 -7218 7235
rect -7276 7167 -7218 7201
rect -7276 7133 -7264 7167
rect -7230 7133 -7218 7167
rect -7276 7099 -7218 7133
rect -7276 7065 -7264 7099
rect -7230 7065 -7218 7099
rect -7276 7031 -7218 7065
rect -7276 6997 -7264 7031
rect -7230 6997 -7218 7031
rect -7276 6963 -7218 6997
rect -7276 6929 -7264 6963
rect -7230 6929 -7218 6963
rect -7276 6895 -7218 6929
rect -7276 6861 -7264 6895
rect -7230 6861 -7218 6895
rect -7276 6827 -7218 6861
rect -7276 6793 -7264 6827
rect -7230 6793 -7218 6827
rect -7276 6759 -7218 6793
rect -7276 6725 -7264 6759
rect -7230 6725 -7218 6759
rect -7276 6691 -7218 6725
rect -7276 6657 -7264 6691
rect -7230 6657 -7218 6691
rect -7276 6623 -7218 6657
rect -7276 6589 -7264 6623
rect -7230 6589 -7218 6623
rect -7276 6555 -7218 6589
rect -7276 6521 -7264 6555
rect -7230 6521 -7218 6555
rect -7276 6487 -7218 6521
rect -7276 6453 -7264 6487
rect -7230 6453 -7218 6487
rect -7276 6419 -7218 6453
rect -7276 6385 -7264 6419
rect -7230 6385 -7218 6419
rect -7276 6351 -7218 6385
rect -7276 6317 -7264 6351
rect -7230 6317 -7218 6351
rect -7276 6283 -7218 6317
rect -7276 6249 -7264 6283
rect -7230 6249 -7218 6283
rect -7276 6215 -7218 6249
rect -7276 6181 -7264 6215
rect -7230 6181 -7218 6215
rect -7276 6147 -7218 6181
rect -7276 6113 -7264 6147
rect -7230 6113 -7218 6147
rect -7276 6079 -7218 6113
rect -7276 6045 -7264 6079
rect -7230 6045 -7218 6079
rect -7276 6011 -7218 6045
rect -7276 5977 -7264 6011
rect -7230 5977 -7218 6011
rect -7276 5943 -7218 5977
rect -7276 5909 -7264 5943
rect -7230 5909 -7218 5943
rect -7276 5875 -7218 5909
rect -7276 5841 -7264 5875
rect -7230 5841 -7218 5875
rect -7276 5807 -7218 5841
rect -7276 5773 -7264 5807
rect -7230 5773 -7218 5807
rect -7276 5739 -7218 5773
rect -7276 5705 -7264 5739
rect -7230 5705 -7218 5739
rect -7276 5671 -7218 5705
rect -7276 5637 -7264 5671
rect -7230 5637 -7218 5671
rect -7276 5603 -7218 5637
rect -7276 5569 -7264 5603
rect -7230 5569 -7218 5603
rect -7276 5538 -7218 5569
rect -7018 7507 -6960 7538
rect -7018 7473 -7006 7507
rect -6972 7473 -6960 7507
rect -7018 7439 -6960 7473
rect -7018 7405 -7006 7439
rect -6972 7405 -6960 7439
rect -7018 7371 -6960 7405
rect -7018 7337 -7006 7371
rect -6972 7337 -6960 7371
rect -7018 7303 -6960 7337
rect -7018 7269 -7006 7303
rect -6972 7269 -6960 7303
rect -7018 7235 -6960 7269
rect -7018 7201 -7006 7235
rect -6972 7201 -6960 7235
rect -7018 7167 -6960 7201
rect -7018 7133 -7006 7167
rect -6972 7133 -6960 7167
rect -7018 7099 -6960 7133
rect -7018 7065 -7006 7099
rect -6972 7065 -6960 7099
rect -7018 7031 -6960 7065
rect -7018 6997 -7006 7031
rect -6972 6997 -6960 7031
rect -7018 6963 -6960 6997
rect -7018 6929 -7006 6963
rect -6972 6929 -6960 6963
rect -7018 6895 -6960 6929
rect -7018 6861 -7006 6895
rect -6972 6861 -6960 6895
rect -7018 6827 -6960 6861
rect -7018 6793 -7006 6827
rect -6972 6793 -6960 6827
rect -7018 6759 -6960 6793
rect -7018 6725 -7006 6759
rect -6972 6725 -6960 6759
rect -7018 6691 -6960 6725
rect -7018 6657 -7006 6691
rect -6972 6657 -6960 6691
rect -7018 6623 -6960 6657
rect -7018 6589 -7006 6623
rect -6972 6589 -6960 6623
rect -7018 6555 -6960 6589
rect -7018 6521 -7006 6555
rect -6972 6521 -6960 6555
rect -7018 6487 -6960 6521
rect -7018 6453 -7006 6487
rect -6972 6453 -6960 6487
rect -7018 6419 -6960 6453
rect -7018 6385 -7006 6419
rect -6972 6385 -6960 6419
rect -7018 6351 -6960 6385
rect -7018 6317 -7006 6351
rect -6972 6317 -6960 6351
rect -7018 6283 -6960 6317
rect -7018 6249 -7006 6283
rect -6972 6249 -6960 6283
rect -7018 6215 -6960 6249
rect -7018 6181 -7006 6215
rect -6972 6181 -6960 6215
rect -7018 6147 -6960 6181
rect -7018 6113 -7006 6147
rect -6972 6113 -6960 6147
rect -7018 6079 -6960 6113
rect -7018 6045 -7006 6079
rect -6972 6045 -6960 6079
rect -7018 6011 -6960 6045
rect -7018 5977 -7006 6011
rect -6972 5977 -6960 6011
rect -7018 5943 -6960 5977
rect -7018 5909 -7006 5943
rect -6972 5909 -6960 5943
rect -7018 5875 -6960 5909
rect -7018 5841 -7006 5875
rect -6972 5841 -6960 5875
rect -7018 5807 -6960 5841
rect -7018 5773 -7006 5807
rect -6972 5773 -6960 5807
rect -7018 5739 -6960 5773
rect -7018 5705 -7006 5739
rect -6972 5705 -6960 5739
rect -7018 5671 -6960 5705
rect -7018 5637 -7006 5671
rect -6972 5637 -6960 5671
rect -7018 5603 -6960 5637
rect -7018 5569 -7006 5603
rect -6972 5569 -6960 5603
rect -7018 5538 -6960 5569
rect -6760 7507 -6702 7538
rect -6760 7473 -6748 7507
rect -6714 7473 -6702 7507
rect -6760 7439 -6702 7473
rect -6760 7405 -6748 7439
rect -6714 7405 -6702 7439
rect -6760 7371 -6702 7405
rect -6760 7337 -6748 7371
rect -6714 7337 -6702 7371
rect -6760 7303 -6702 7337
rect -6760 7269 -6748 7303
rect -6714 7269 -6702 7303
rect -6760 7235 -6702 7269
rect -6760 7201 -6748 7235
rect -6714 7201 -6702 7235
rect -6760 7167 -6702 7201
rect -6760 7133 -6748 7167
rect -6714 7133 -6702 7167
rect -6760 7099 -6702 7133
rect -6760 7065 -6748 7099
rect -6714 7065 -6702 7099
rect -6760 7031 -6702 7065
rect -6760 6997 -6748 7031
rect -6714 6997 -6702 7031
rect -6760 6963 -6702 6997
rect -6760 6929 -6748 6963
rect -6714 6929 -6702 6963
rect -6760 6895 -6702 6929
rect -6760 6861 -6748 6895
rect -6714 6861 -6702 6895
rect -6760 6827 -6702 6861
rect -6760 6793 -6748 6827
rect -6714 6793 -6702 6827
rect -6760 6759 -6702 6793
rect -6760 6725 -6748 6759
rect -6714 6725 -6702 6759
rect -6760 6691 -6702 6725
rect -6760 6657 -6748 6691
rect -6714 6657 -6702 6691
rect -6760 6623 -6702 6657
rect -6760 6589 -6748 6623
rect -6714 6589 -6702 6623
rect -6760 6555 -6702 6589
rect -6760 6521 -6748 6555
rect -6714 6521 -6702 6555
rect -6760 6487 -6702 6521
rect -6760 6453 -6748 6487
rect -6714 6453 -6702 6487
rect -6760 6419 -6702 6453
rect -6760 6385 -6748 6419
rect -6714 6385 -6702 6419
rect -6760 6351 -6702 6385
rect -6760 6317 -6748 6351
rect -6714 6317 -6702 6351
rect -6760 6283 -6702 6317
rect -6760 6249 -6748 6283
rect -6714 6249 -6702 6283
rect -6760 6215 -6702 6249
rect -6760 6181 -6748 6215
rect -6714 6181 -6702 6215
rect -6760 6147 -6702 6181
rect -6760 6113 -6748 6147
rect -6714 6113 -6702 6147
rect -6760 6079 -6702 6113
rect -6760 6045 -6748 6079
rect -6714 6045 -6702 6079
rect -6760 6011 -6702 6045
rect -6760 5977 -6748 6011
rect -6714 5977 -6702 6011
rect -6760 5943 -6702 5977
rect -6760 5909 -6748 5943
rect -6714 5909 -6702 5943
rect -6760 5875 -6702 5909
rect -6760 5841 -6748 5875
rect -6714 5841 -6702 5875
rect -6760 5807 -6702 5841
rect -6760 5773 -6748 5807
rect -6714 5773 -6702 5807
rect -6760 5739 -6702 5773
rect -6760 5705 -6748 5739
rect -6714 5705 -6702 5739
rect -6760 5671 -6702 5705
rect -6760 5637 -6748 5671
rect -6714 5637 -6702 5671
rect -6760 5603 -6702 5637
rect -6760 5569 -6748 5603
rect -6714 5569 -6702 5603
rect -6760 5538 -6702 5569
rect -6502 7507 -6444 7538
rect -6502 7473 -6490 7507
rect -6456 7473 -6444 7507
rect -6502 7439 -6444 7473
rect -6502 7405 -6490 7439
rect -6456 7405 -6444 7439
rect -6502 7371 -6444 7405
rect -6502 7337 -6490 7371
rect -6456 7337 -6444 7371
rect -6502 7303 -6444 7337
rect -6502 7269 -6490 7303
rect -6456 7269 -6444 7303
rect -6502 7235 -6444 7269
rect -6502 7201 -6490 7235
rect -6456 7201 -6444 7235
rect -6502 7167 -6444 7201
rect -6502 7133 -6490 7167
rect -6456 7133 -6444 7167
rect -6502 7099 -6444 7133
rect -6502 7065 -6490 7099
rect -6456 7065 -6444 7099
rect -6502 7031 -6444 7065
rect -6502 6997 -6490 7031
rect -6456 6997 -6444 7031
rect -6502 6963 -6444 6997
rect -6502 6929 -6490 6963
rect -6456 6929 -6444 6963
rect -6502 6895 -6444 6929
rect -6502 6861 -6490 6895
rect -6456 6861 -6444 6895
rect -6502 6827 -6444 6861
rect -6502 6793 -6490 6827
rect -6456 6793 -6444 6827
rect -6502 6759 -6444 6793
rect -6502 6725 -6490 6759
rect -6456 6725 -6444 6759
rect -6502 6691 -6444 6725
rect -6502 6657 -6490 6691
rect -6456 6657 -6444 6691
rect -6502 6623 -6444 6657
rect -6502 6589 -6490 6623
rect -6456 6589 -6444 6623
rect -6502 6555 -6444 6589
rect -6502 6521 -6490 6555
rect -6456 6521 -6444 6555
rect -6502 6487 -6444 6521
rect -6502 6453 -6490 6487
rect -6456 6453 -6444 6487
rect -6502 6419 -6444 6453
rect -6502 6385 -6490 6419
rect -6456 6385 -6444 6419
rect -6502 6351 -6444 6385
rect -6502 6317 -6490 6351
rect -6456 6317 -6444 6351
rect -6502 6283 -6444 6317
rect -6502 6249 -6490 6283
rect -6456 6249 -6444 6283
rect -6502 6215 -6444 6249
rect -6502 6181 -6490 6215
rect -6456 6181 -6444 6215
rect -6502 6147 -6444 6181
rect -6502 6113 -6490 6147
rect -6456 6113 -6444 6147
rect -6502 6079 -6444 6113
rect -6502 6045 -6490 6079
rect -6456 6045 -6444 6079
rect -6502 6011 -6444 6045
rect -6502 5977 -6490 6011
rect -6456 5977 -6444 6011
rect -6502 5943 -6444 5977
rect -6502 5909 -6490 5943
rect -6456 5909 -6444 5943
rect -6502 5875 -6444 5909
rect -6502 5841 -6490 5875
rect -6456 5841 -6444 5875
rect -6502 5807 -6444 5841
rect -6502 5773 -6490 5807
rect -6456 5773 -6444 5807
rect -6502 5739 -6444 5773
rect -6502 5705 -6490 5739
rect -6456 5705 -6444 5739
rect -6502 5671 -6444 5705
rect -6502 5637 -6490 5671
rect -6456 5637 -6444 5671
rect -6502 5603 -6444 5637
rect -6502 5569 -6490 5603
rect -6456 5569 -6444 5603
rect -6502 5538 -6444 5569
rect -6244 7507 -6186 7538
rect -6244 7473 -6232 7507
rect -6198 7473 -6186 7507
rect -6244 7439 -6186 7473
rect -6244 7405 -6232 7439
rect -6198 7405 -6186 7439
rect -6244 7371 -6186 7405
rect -6244 7337 -6232 7371
rect -6198 7337 -6186 7371
rect -6244 7303 -6186 7337
rect -6244 7269 -6232 7303
rect -6198 7269 -6186 7303
rect -6244 7235 -6186 7269
rect -6244 7201 -6232 7235
rect -6198 7201 -6186 7235
rect -6244 7167 -6186 7201
rect -6244 7133 -6232 7167
rect -6198 7133 -6186 7167
rect -6244 7099 -6186 7133
rect -6244 7065 -6232 7099
rect -6198 7065 -6186 7099
rect -6244 7031 -6186 7065
rect -6244 6997 -6232 7031
rect -6198 6997 -6186 7031
rect -6244 6963 -6186 6997
rect -6244 6929 -6232 6963
rect -6198 6929 -6186 6963
rect -6244 6895 -6186 6929
rect -6244 6861 -6232 6895
rect -6198 6861 -6186 6895
rect -6244 6827 -6186 6861
rect -6244 6793 -6232 6827
rect -6198 6793 -6186 6827
rect -6244 6759 -6186 6793
rect -6244 6725 -6232 6759
rect -6198 6725 -6186 6759
rect -6244 6691 -6186 6725
rect -6244 6657 -6232 6691
rect -6198 6657 -6186 6691
rect -6244 6623 -6186 6657
rect -6244 6589 -6232 6623
rect -6198 6589 -6186 6623
rect -6244 6555 -6186 6589
rect -6244 6521 -6232 6555
rect -6198 6521 -6186 6555
rect -6244 6487 -6186 6521
rect -6244 6453 -6232 6487
rect -6198 6453 -6186 6487
rect -6244 6419 -6186 6453
rect -6244 6385 -6232 6419
rect -6198 6385 -6186 6419
rect -6244 6351 -6186 6385
rect -6244 6317 -6232 6351
rect -6198 6317 -6186 6351
rect -6244 6283 -6186 6317
rect -6244 6249 -6232 6283
rect -6198 6249 -6186 6283
rect -6244 6215 -6186 6249
rect -6244 6181 -6232 6215
rect -6198 6181 -6186 6215
rect -6244 6147 -6186 6181
rect -6244 6113 -6232 6147
rect -6198 6113 -6186 6147
rect -6244 6079 -6186 6113
rect -6244 6045 -6232 6079
rect -6198 6045 -6186 6079
rect -6244 6011 -6186 6045
rect -6244 5977 -6232 6011
rect -6198 5977 -6186 6011
rect -6244 5943 -6186 5977
rect -6244 5909 -6232 5943
rect -6198 5909 -6186 5943
rect -6244 5875 -6186 5909
rect -6244 5841 -6232 5875
rect -6198 5841 -6186 5875
rect -6244 5807 -6186 5841
rect -6244 5773 -6232 5807
rect -6198 5773 -6186 5807
rect -6244 5739 -6186 5773
rect -6244 5705 -6232 5739
rect -6198 5705 -6186 5739
rect -6244 5671 -6186 5705
rect -6244 5637 -6232 5671
rect -6198 5637 -6186 5671
rect -6244 5603 -6186 5637
rect -6244 5569 -6232 5603
rect -6198 5569 -6186 5603
rect -6244 5538 -6186 5569
rect -5986 7507 -5928 7538
rect -5986 7473 -5974 7507
rect -5940 7473 -5928 7507
rect -5986 7439 -5928 7473
rect -5986 7405 -5974 7439
rect -5940 7405 -5928 7439
rect -5986 7371 -5928 7405
rect -5986 7337 -5974 7371
rect -5940 7337 -5928 7371
rect -5986 7303 -5928 7337
rect -5986 7269 -5974 7303
rect -5940 7269 -5928 7303
rect -5986 7235 -5928 7269
rect -5986 7201 -5974 7235
rect -5940 7201 -5928 7235
rect -5986 7167 -5928 7201
rect -5986 7133 -5974 7167
rect -5940 7133 -5928 7167
rect -5986 7099 -5928 7133
rect -5986 7065 -5974 7099
rect -5940 7065 -5928 7099
rect -5986 7031 -5928 7065
rect -5986 6997 -5974 7031
rect -5940 6997 -5928 7031
rect -5986 6963 -5928 6997
rect -5986 6929 -5974 6963
rect -5940 6929 -5928 6963
rect -5986 6895 -5928 6929
rect -5986 6861 -5974 6895
rect -5940 6861 -5928 6895
rect -5986 6827 -5928 6861
rect -5986 6793 -5974 6827
rect -5940 6793 -5928 6827
rect -5986 6759 -5928 6793
rect -5986 6725 -5974 6759
rect -5940 6725 -5928 6759
rect -5986 6691 -5928 6725
rect -5986 6657 -5974 6691
rect -5940 6657 -5928 6691
rect -5986 6623 -5928 6657
rect -5986 6589 -5974 6623
rect -5940 6589 -5928 6623
rect -5986 6555 -5928 6589
rect -5986 6521 -5974 6555
rect -5940 6521 -5928 6555
rect -5986 6487 -5928 6521
rect -5986 6453 -5974 6487
rect -5940 6453 -5928 6487
rect -5986 6419 -5928 6453
rect -5986 6385 -5974 6419
rect -5940 6385 -5928 6419
rect -5986 6351 -5928 6385
rect -5986 6317 -5974 6351
rect -5940 6317 -5928 6351
rect -5986 6283 -5928 6317
rect -5986 6249 -5974 6283
rect -5940 6249 -5928 6283
rect -5986 6215 -5928 6249
rect -5986 6181 -5974 6215
rect -5940 6181 -5928 6215
rect -5986 6147 -5928 6181
rect -5986 6113 -5974 6147
rect -5940 6113 -5928 6147
rect -5986 6079 -5928 6113
rect -5986 6045 -5974 6079
rect -5940 6045 -5928 6079
rect -5986 6011 -5928 6045
rect -5986 5977 -5974 6011
rect -5940 5977 -5928 6011
rect -5986 5943 -5928 5977
rect -5986 5909 -5974 5943
rect -5940 5909 -5928 5943
rect -5986 5875 -5928 5909
rect -5986 5841 -5974 5875
rect -5940 5841 -5928 5875
rect -5986 5807 -5928 5841
rect -5986 5773 -5974 5807
rect -5940 5773 -5928 5807
rect -5986 5739 -5928 5773
rect -5986 5705 -5974 5739
rect -5940 5705 -5928 5739
rect -5986 5671 -5928 5705
rect -5986 5637 -5974 5671
rect -5940 5637 -5928 5671
rect -5986 5603 -5928 5637
rect -5986 5569 -5974 5603
rect -5940 5569 -5928 5603
rect -5986 5538 -5928 5569
rect -5728 7507 -5670 7538
rect -5728 7473 -5716 7507
rect -5682 7473 -5670 7507
rect -5728 7439 -5670 7473
rect -5728 7405 -5716 7439
rect -5682 7405 -5670 7439
rect -5728 7371 -5670 7405
rect -5728 7337 -5716 7371
rect -5682 7337 -5670 7371
rect -5728 7303 -5670 7337
rect -5728 7269 -5716 7303
rect -5682 7269 -5670 7303
rect -5728 7235 -5670 7269
rect -5728 7201 -5716 7235
rect -5682 7201 -5670 7235
rect -5728 7167 -5670 7201
rect -5728 7133 -5716 7167
rect -5682 7133 -5670 7167
rect -5728 7099 -5670 7133
rect -5728 7065 -5716 7099
rect -5682 7065 -5670 7099
rect -5728 7031 -5670 7065
rect -5728 6997 -5716 7031
rect -5682 6997 -5670 7031
rect -5728 6963 -5670 6997
rect -5728 6929 -5716 6963
rect -5682 6929 -5670 6963
rect -5728 6895 -5670 6929
rect -5728 6861 -5716 6895
rect -5682 6861 -5670 6895
rect -5728 6827 -5670 6861
rect -5728 6793 -5716 6827
rect -5682 6793 -5670 6827
rect -5728 6759 -5670 6793
rect -5728 6725 -5716 6759
rect -5682 6725 -5670 6759
rect -5728 6691 -5670 6725
rect -5728 6657 -5716 6691
rect -5682 6657 -5670 6691
rect -5728 6623 -5670 6657
rect -5728 6589 -5716 6623
rect -5682 6589 -5670 6623
rect -5728 6555 -5670 6589
rect -5728 6521 -5716 6555
rect -5682 6521 -5670 6555
rect -5728 6487 -5670 6521
rect -5728 6453 -5716 6487
rect -5682 6453 -5670 6487
rect -5728 6419 -5670 6453
rect -5728 6385 -5716 6419
rect -5682 6385 -5670 6419
rect -5728 6351 -5670 6385
rect -5728 6317 -5716 6351
rect -5682 6317 -5670 6351
rect -5728 6283 -5670 6317
rect -5728 6249 -5716 6283
rect -5682 6249 -5670 6283
rect -5728 6215 -5670 6249
rect -5728 6181 -5716 6215
rect -5682 6181 -5670 6215
rect -5728 6147 -5670 6181
rect -5728 6113 -5716 6147
rect -5682 6113 -5670 6147
rect -5728 6079 -5670 6113
rect -5728 6045 -5716 6079
rect -5682 6045 -5670 6079
rect -5728 6011 -5670 6045
rect -5728 5977 -5716 6011
rect -5682 5977 -5670 6011
rect -5728 5943 -5670 5977
rect -5728 5909 -5716 5943
rect -5682 5909 -5670 5943
rect -5728 5875 -5670 5909
rect -5728 5841 -5716 5875
rect -5682 5841 -5670 5875
rect -5728 5807 -5670 5841
rect -5728 5773 -5716 5807
rect -5682 5773 -5670 5807
rect -5728 5739 -5670 5773
rect -5728 5705 -5716 5739
rect -5682 5705 -5670 5739
rect -5728 5671 -5670 5705
rect -5728 5637 -5716 5671
rect -5682 5637 -5670 5671
rect -5728 5603 -5670 5637
rect -5728 5569 -5716 5603
rect -5682 5569 -5670 5603
rect -5728 5538 -5670 5569
rect -5470 7507 -5412 7538
rect -5470 7473 -5458 7507
rect -5424 7473 -5412 7507
rect -5470 7439 -5412 7473
rect -5470 7405 -5458 7439
rect -5424 7405 -5412 7439
rect -5470 7371 -5412 7405
rect -5470 7337 -5458 7371
rect -5424 7337 -5412 7371
rect -5470 7303 -5412 7337
rect -5470 7269 -5458 7303
rect -5424 7269 -5412 7303
rect -5470 7235 -5412 7269
rect -5470 7201 -5458 7235
rect -5424 7201 -5412 7235
rect -5470 7167 -5412 7201
rect -5470 7133 -5458 7167
rect -5424 7133 -5412 7167
rect -5470 7099 -5412 7133
rect -5470 7065 -5458 7099
rect -5424 7065 -5412 7099
rect -5470 7031 -5412 7065
rect -5470 6997 -5458 7031
rect -5424 6997 -5412 7031
rect -5470 6963 -5412 6997
rect -5470 6929 -5458 6963
rect -5424 6929 -5412 6963
rect -5470 6895 -5412 6929
rect -5470 6861 -5458 6895
rect -5424 6861 -5412 6895
rect -5470 6827 -5412 6861
rect -5470 6793 -5458 6827
rect -5424 6793 -5412 6827
rect -5470 6759 -5412 6793
rect -5470 6725 -5458 6759
rect -5424 6725 -5412 6759
rect -5470 6691 -5412 6725
rect -5470 6657 -5458 6691
rect -5424 6657 -5412 6691
rect -5470 6623 -5412 6657
rect -5470 6589 -5458 6623
rect -5424 6589 -5412 6623
rect -5470 6555 -5412 6589
rect -5470 6521 -5458 6555
rect -5424 6521 -5412 6555
rect -5470 6487 -5412 6521
rect -5470 6453 -5458 6487
rect -5424 6453 -5412 6487
rect -5470 6419 -5412 6453
rect -5470 6385 -5458 6419
rect -5424 6385 -5412 6419
rect -5470 6351 -5412 6385
rect -5470 6317 -5458 6351
rect -5424 6317 -5412 6351
rect -5470 6283 -5412 6317
rect -5470 6249 -5458 6283
rect -5424 6249 -5412 6283
rect -5470 6215 -5412 6249
rect -5470 6181 -5458 6215
rect -5424 6181 -5412 6215
rect -5470 6147 -5412 6181
rect -5470 6113 -5458 6147
rect -5424 6113 -5412 6147
rect -5470 6079 -5412 6113
rect -5470 6045 -5458 6079
rect -5424 6045 -5412 6079
rect -5470 6011 -5412 6045
rect -5470 5977 -5458 6011
rect -5424 5977 -5412 6011
rect -5470 5943 -5412 5977
rect -5470 5909 -5458 5943
rect -5424 5909 -5412 5943
rect -5470 5875 -5412 5909
rect -5470 5841 -5458 5875
rect -5424 5841 -5412 5875
rect -5470 5807 -5412 5841
rect -5470 5773 -5458 5807
rect -5424 5773 -5412 5807
rect -5470 5739 -5412 5773
rect -5470 5705 -5458 5739
rect -5424 5705 -5412 5739
rect -5470 5671 -5412 5705
rect -5470 5637 -5458 5671
rect -5424 5637 -5412 5671
rect -5470 5603 -5412 5637
rect -5470 5569 -5458 5603
rect -5424 5569 -5412 5603
rect -5470 5538 -5412 5569
rect -5212 7507 -5154 7538
rect -5212 7473 -5200 7507
rect -5166 7473 -5154 7507
rect -5212 7439 -5154 7473
rect -5212 7405 -5200 7439
rect -5166 7405 -5154 7439
rect -5212 7371 -5154 7405
rect -5212 7337 -5200 7371
rect -5166 7337 -5154 7371
rect -5212 7303 -5154 7337
rect -5212 7269 -5200 7303
rect -5166 7269 -5154 7303
rect -5212 7235 -5154 7269
rect -5212 7201 -5200 7235
rect -5166 7201 -5154 7235
rect -5212 7167 -5154 7201
rect -5212 7133 -5200 7167
rect -5166 7133 -5154 7167
rect -5212 7099 -5154 7133
rect -5212 7065 -5200 7099
rect -5166 7065 -5154 7099
rect -5212 7031 -5154 7065
rect -5212 6997 -5200 7031
rect -5166 6997 -5154 7031
rect -5212 6963 -5154 6997
rect -5212 6929 -5200 6963
rect -5166 6929 -5154 6963
rect -5212 6895 -5154 6929
rect -5212 6861 -5200 6895
rect -5166 6861 -5154 6895
rect -5212 6827 -5154 6861
rect -5212 6793 -5200 6827
rect -5166 6793 -5154 6827
rect -5212 6759 -5154 6793
rect -5212 6725 -5200 6759
rect -5166 6725 -5154 6759
rect -5212 6691 -5154 6725
rect -5212 6657 -5200 6691
rect -5166 6657 -5154 6691
rect -5212 6623 -5154 6657
rect -5212 6589 -5200 6623
rect -5166 6589 -5154 6623
rect -5212 6555 -5154 6589
rect -5212 6521 -5200 6555
rect -5166 6521 -5154 6555
rect -5212 6487 -5154 6521
rect -5212 6453 -5200 6487
rect -5166 6453 -5154 6487
rect -5212 6419 -5154 6453
rect -5212 6385 -5200 6419
rect -5166 6385 -5154 6419
rect -5212 6351 -5154 6385
rect -5212 6317 -5200 6351
rect -5166 6317 -5154 6351
rect -5212 6283 -5154 6317
rect -5212 6249 -5200 6283
rect -5166 6249 -5154 6283
rect -5212 6215 -5154 6249
rect -5212 6181 -5200 6215
rect -5166 6181 -5154 6215
rect -5212 6147 -5154 6181
rect -5212 6113 -5200 6147
rect -5166 6113 -5154 6147
rect -5212 6079 -5154 6113
rect -5212 6045 -5200 6079
rect -5166 6045 -5154 6079
rect -5212 6011 -5154 6045
rect -5212 5977 -5200 6011
rect -5166 5977 -5154 6011
rect -5212 5943 -5154 5977
rect -5212 5909 -5200 5943
rect -5166 5909 -5154 5943
rect -5212 5875 -5154 5909
rect -5212 5841 -5200 5875
rect -5166 5841 -5154 5875
rect -5212 5807 -5154 5841
rect -5212 5773 -5200 5807
rect -5166 5773 -5154 5807
rect -5212 5739 -5154 5773
rect -5212 5705 -5200 5739
rect -5166 5705 -5154 5739
rect -5212 5671 -5154 5705
rect -5212 5637 -5200 5671
rect -5166 5637 -5154 5671
rect -5212 5603 -5154 5637
rect -5212 5569 -5200 5603
rect -5166 5569 -5154 5603
rect -5212 5538 -5154 5569
rect -4954 7507 -4896 7538
rect -4954 7473 -4942 7507
rect -4908 7473 -4896 7507
rect -4954 7439 -4896 7473
rect -4954 7405 -4942 7439
rect -4908 7405 -4896 7439
rect -4954 7371 -4896 7405
rect -4954 7337 -4942 7371
rect -4908 7337 -4896 7371
rect -4954 7303 -4896 7337
rect -4954 7269 -4942 7303
rect -4908 7269 -4896 7303
rect -4954 7235 -4896 7269
rect -4954 7201 -4942 7235
rect -4908 7201 -4896 7235
rect -4954 7167 -4896 7201
rect -4954 7133 -4942 7167
rect -4908 7133 -4896 7167
rect -4954 7099 -4896 7133
rect -4954 7065 -4942 7099
rect -4908 7065 -4896 7099
rect -4954 7031 -4896 7065
rect -4954 6997 -4942 7031
rect -4908 6997 -4896 7031
rect -4954 6963 -4896 6997
rect -4954 6929 -4942 6963
rect -4908 6929 -4896 6963
rect -4954 6895 -4896 6929
rect -4954 6861 -4942 6895
rect -4908 6861 -4896 6895
rect -4954 6827 -4896 6861
rect -4954 6793 -4942 6827
rect -4908 6793 -4896 6827
rect -4954 6759 -4896 6793
rect -4954 6725 -4942 6759
rect -4908 6725 -4896 6759
rect -4954 6691 -4896 6725
rect -4954 6657 -4942 6691
rect -4908 6657 -4896 6691
rect -4954 6623 -4896 6657
rect -4954 6589 -4942 6623
rect -4908 6589 -4896 6623
rect -4954 6555 -4896 6589
rect -4954 6521 -4942 6555
rect -4908 6521 -4896 6555
rect -4954 6487 -4896 6521
rect -4954 6453 -4942 6487
rect -4908 6453 -4896 6487
rect -4954 6419 -4896 6453
rect -4954 6385 -4942 6419
rect -4908 6385 -4896 6419
rect -4954 6351 -4896 6385
rect -4954 6317 -4942 6351
rect -4908 6317 -4896 6351
rect -4954 6283 -4896 6317
rect -4954 6249 -4942 6283
rect -4908 6249 -4896 6283
rect -4954 6215 -4896 6249
rect -4954 6181 -4942 6215
rect -4908 6181 -4896 6215
rect -4954 6147 -4896 6181
rect -4954 6113 -4942 6147
rect -4908 6113 -4896 6147
rect -4954 6079 -4896 6113
rect -4954 6045 -4942 6079
rect -4908 6045 -4896 6079
rect -4954 6011 -4896 6045
rect -4954 5977 -4942 6011
rect -4908 5977 -4896 6011
rect -4954 5943 -4896 5977
rect -4954 5909 -4942 5943
rect -4908 5909 -4896 5943
rect -4954 5875 -4896 5909
rect -4954 5841 -4942 5875
rect -4908 5841 -4896 5875
rect -4954 5807 -4896 5841
rect -4954 5773 -4942 5807
rect -4908 5773 -4896 5807
rect -4954 5739 -4896 5773
rect -4954 5705 -4942 5739
rect -4908 5705 -4896 5739
rect -4954 5671 -4896 5705
rect -4954 5637 -4942 5671
rect -4908 5637 -4896 5671
rect -4954 5603 -4896 5637
rect -4954 5569 -4942 5603
rect -4908 5569 -4896 5603
rect -4954 5538 -4896 5569
rect -4696 7507 -4638 7538
rect -4696 7473 -4684 7507
rect -4650 7473 -4638 7507
rect -4696 7439 -4638 7473
rect -4696 7405 -4684 7439
rect -4650 7405 -4638 7439
rect -4696 7371 -4638 7405
rect -4696 7337 -4684 7371
rect -4650 7337 -4638 7371
rect -4696 7303 -4638 7337
rect -4696 7269 -4684 7303
rect -4650 7269 -4638 7303
rect -4696 7235 -4638 7269
rect -4696 7201 -4684 7235
rect -4650 7201 -4638 7235
rect -4696 7167 -4638 7201
rect -4696 7133 -4684 7167
rect -4650 7133 -4638 7167
rect -4696 7099 -4638 7133
rect -4696 7065 -4684 7099
rect -4650 7065 -4638 7099
rect -4696 7031 -4638 7065
rect -4696 6997 -4684 7031
rect -4650 6997 -4638 7031
rect -4696 6963 -4638 6997
rect -4696 6929 -4684 6963
rect -4650 6929 -4638 6963
rect -4696 6895 -4638 6929
rect -4696 6861 -4684 6895
rect -4650 6861 -4638 6895
rect -4696 6827 -4638 6861
rect -4696 6793 -4684 6827
rect -4650 6793 -4638 6827
rect -4696 6759 -4638 6793
rect -4696 6725 -4684 6759
rect -4650 6725 -4638 6759
rect -4696 6691 -4638 6725
rect -4696 6657 -4684 6691
rect -4650 6657 -4638 6691
rect -4696 6623 -4638 6657
rect -4696 6589 -4684 6623
rect -4650 6589 -4638 6623
rect -4696 6555 -4638 6589
rect -4696 6521 -4684 6555
rect -4650 6521 -4638 6555
rect -4696 6487 -4638 6521
rect -4696 6453 -4684 6487
rect -4650 6453 -4638 6487
rect -4696 6419 -4638 6453
rect -4696 6385 -4684 6419
rect -4650 6385 -4638 6419
rect -4696 6351 -4638 6385
rect -4696 6317 -4684 6351
rect -4650 6317 -4638 6351
rect -4696 6283 -4638 6317
rect -4696 6249 -4684 6283
rect -4650 6249 -4638 6283
rect -4696 6215 -4638 6249
rect -4696 6181 -4684 6215
rect -4650 6181 -4638 6215
rect -4696 6147 -4638 6181
rect -4696 6113 -4684 6147
rect -4650 6113 -4638 6147
rect -4696 6079 -4638 6113
rect -4696 6045 -4684 6079
rect -4650 6045 -4638 6079
rect -4696 6011 -4638 6045
rect -4696 5977 -4684 6011
rect -4650 5977 -4638 6011
rect -4696 5943 -4638 5977
rect -4696 5909 -4684 5943
rect -4650 5909 -4638 5943
rect -4696 5875 -4638 5909
rect -4696 5841 -4684 5875
rect -4650 5841 -4638 5875
rect -4696 5807 -4638 5841
rect -4696 5773 -4684 5807
rect -4650 5773 -4638 5807
rect -4696 5739 -4638 5773
rect -4696 5705 -4684 5739
rect -4650 5705 -4638 5739
rect -4696 5671 -4638 5705
rect -4696 5637 -4684 5671
rect -4650 5637 -4638 5671
rect -4696 5603 -4638 5637
rect -4696 5569 -4684 5603
rect -4650 5569 -4638 5603
rect -4696 5538 -4638 5569
rect -4438 7507 -4380 7538
rect -4438 7473 -4426 7507
rect -4392 7473 -4380 7507
rect -4438 7439 -4380 7473
rect -4438 7405 -4426 7439
rect -4392 7405 -4380 7439
rect -4438 7371 -4380 7405
rect -4438 7337 -4426 7371
rect -4392 7337 -4380 7371
rect -4438 7303 -4380 7337
rect -4438 7269 -4426 7303
rect -4392 7269 -4380 7303
rect -4438 7235 -4380 7269
rect -4438 7201 -4426 7235
rect -4392 7201 -4380 7235
rect -4438 7167 -4380 7201
rect -4438 7133 -4426 7167
rect -4392 7133 -4380 7167
rect -4438 7099 -4380 7133
rect -4438 7065 -4426 7099
rect -4392 7065 -4380 7099
rect -4438 7031 -4380 7065
rect -4438 6997 -4426 7031
rect -4392 6997 -4380 7031
rect -4438 6963 -4380 6997
rect -4438 6929 -4426 6963
rect -4392 6929 -4380 6963
rect -4438 6895 -4380 6929
rect -4438 6861 -4426 6895
rect -4392 6861 -4380 6895
rect -4438 6827 -4380 6861
rect -4438 6793 -4426 6827
rect -4392 6793 -4380 6827
rect -4438 6759 -4380 6793
rect -4438 6725 -4426 6759
rect -4392 6725 -4380 6759
rect -4438 6691 -4380 6725
rect -4438 6657 -4426 6691
rect -4392 6657 -4380 6691
rect -4438 6623 -4380 6657
rect -4438 6589 -4426 6623
rect -4392 6589 -4380 6623
rect -4438 6555 -4380 6589
rect -4438 6521 -4426 6555
rect -4392 6521 -4380 6555
rect -4438 6487 -4380 6521
rect -4438 6453 -4426 6487
rect -4392 6453 -4380 6487
rect -4438 6419 -4380 6453
rect -4438 6385 -4426 6419
rect -4392 6385 -4380 6419
rect -4438 6351 -4380 6385
rect -4438 6317 -4426 6351
rect -4392 6317 -4380 6351
rect -4438 6283 -4380 6317
rect -4438 6249 -4426 6283
rect -4392 6249 -4380 6283
rect -4438 6215 -4380 6249
rect -4438 6181 -4426 6215
rect -4392 6181 -4380 6215
rect -4438 6147 -4380 6181
rect -4438 6113 -4426 6147
rect -4392 6113 -4380 6147
rect -4438 6079 -4380 6113
rect -4438 6045 -4426 6079
rect -4392 6045 -4380 6079
rect -4438 6011 -4380 6045
rect -4438 5977 -4426 6011
rect -4392 5977 -4380 6011
rect -4438 5943 -4380 5977
rect -4438 5909 -4426 5943
rect -4392 5909 -4380 5943
rect -4438 5875 -4380 5909
rect -4438 5841 -4426 5875
rect -4392 5841 -4380 5875
rect -4438 5807 -4380 5841
rect -4438 5773 -4426 5807
rect -4392 5773 -4380 5807
rect -4438 5739 -4380 5773
rect -4438 5705 -4426 5739
rect -4392 5705 -4380 5739
rect -4438 5671 -4380 5705
rect -4438 5637 -4426 5671
rect -4392 5637 -4380 5671
rect -4438 5603 -4380 5637
rect -4438 5569 -4426 5603
rect -4392 5569 -4380 5603
rect -4438 5538 -4380 5569
rect -4180 7507 -4122 7538
rect -4180 7473 -4168 7507
rect -4134 7473 -4122 7507
rect -4180 7439 -4122 7473
rect -4180 7405 -4168 7439
rect -4134 7405 -4122 7439
rect -4180 7371 -4122 7405
rect -4180 7337 -4168 7371
rect -4134 7337 -4122 7371
rect -4180 7303 -4122 7337
rect -4180 7269 -4168 7303
rect -4134 7269 -4122 7303
rect -4180 7235 -4122 7269
rect -4180 7201 -4168 7235
rect -4134 7201 -4122 7235
rect -4180 7167 -4122 7201
rect -4180 7133 -4168 7167
rect -4134 7133 -4122 7167
rect -4180 7099 -4122 7133
rect -4180 7065 -4168 7099
rect -4134 7065 -4122 7099
rect -4180 7031 -4122 7065
rect -4180 6997 -4168 7031
rect -4134 6997 -4122 7031
rect -4180 6963 -4122 6997
rect -4180 6929 -4168 6963
rect -4134 6929 -4122 6963
rect -4180 6895 -4122 6929
rect -4180 6861 -4168 6895
rect -4134 6861 -4122 6895
rect -4180 6827 -4122 6861
rect -4180 6793 -4168 6827
rect -4134 6793 -4122 6827
rect -4180 6759 -4122 6793
rect -4180 6725 -4168 6759
rect -4134 6725 -4122 6759
rect -4180 6691 -4122 6725
rect -4180 6657 -4168 6691
rect -4134 6657 -4122 6691
rect -4180 6623 -4122 6657
rect -4180 6589 -4168 6623
rect -4134 6589 -4122 6623
rect -4180 6555 -4122 6589
rect -4180 6521 -4168 6555
rect -4134 6521 -4122 6555
rect -4180 6487 -4122 6521
rect -4180 6453 -4168 6487
rect -4134 6453 -4122 6487
rect -4180 6419 -4122 6453
rect -4180 6385 -4168 6419
rect -4134 6385 -4122 6419
rect -4180 6351 -4122 6385
rect -4180 6317 -4168 6351
rect -4134 6317 -4122 6351
rect -4180 6283 -4122 6317
rect -4180 6249 -4168 6283
rect -4134 6249 -4122 6283
rect -4180 6215 -4122 6249
rect -4180 6181 -4168 6215
rect -4134 6181 -4122 6215
rect -4180 6147 -4122 6181
rect -4180 6113 -4168 6147
rect -4134 6113 -4122 6147
rect -4180 6079 -4122 6113
rect -4180 6045 -4168 6079
rect -4134 6045 -4122 6079
rect -4180 6011 -4122 6045
rect -4180 5977 -4168 6011
rect -4134 5977 -4122 6011
rect -4180 5943 -4122 5977
rect -4180 5909 -4168 5943
rect -4134 5909 -4122 5943
rect -4180 5875 -4122 5909
rect -4180 5841 -4168 5875
rect -4134 5841 -4122 5875
rect -4180 5807 -4122 5841
rect -4180 5773 -4168 5807
rect -4134 5773 -4122 5807
rect -4180 5739 -4122 5773
rect -4180 5705 -4168 5739
rect -4134 5705 -4122 5739
rect -4180 5671 -4122 5705
rect -4180 5637 -4168 5671
rect -4134 5637 -4122 5671
rect -4180 5603 -4122 5637
rect -4180 5569 -4168 5603
rect -4134 5569 -4122 5603
rect -4180 5538 -4122 5569
rect -3922 7507 -3864 7538
rect -3922 7473 -3910 7507
rect -3876 7473 -3864 7507
rect -3922 7439 -3864 7473
rect -3922 7405 -3910 7439
rect -3876 7405 -3864 7439
rect -3922 7371 -3864 7405
rect -3922 7337 -3910 7371
rect -3876 7337 -3864 7371
rect -3922 7303 -3864 7337
rect -3922 7269 -3910 7303
rect -3876 7269 -3864 7303
rect -3922 7235 -3864 7269
rect -3922 7201 -3910 7235
rect -3876 7201 -3864 7235
rect -3922 7167 -3864 7201
rect -3922 7133 -3910 7167
rect -3876 7133 -3864 7167
rect -3922 7099 -3864 7133
rect -3922 7065 -3910 7099
rect -3876 7065 -3864 7099
rect -3922 7031 -3864 7065
rect -3922 6997 -3910 7031
rect -3876 6997 -3864 7031
rect -3922 6963 -3864 6997
rect -3922 6929 -3910 6963
rect -3876 6929 -3864 6963
rect -3922 6895 -3864 6929
rect -3922 6861 -3910 6895
rect -3876 6861 -3864 6895
rect -3922 6827 -3864 6861
rect -3922 6793 -3910 6827
rect -3876 6793 -3864 6827
rect -3922 6759 -3864 6793
rect -3922 6725 -3910 6759
rect -3876 6725 -3864 6759
rect -3922 6691 -3864 6725
rect -3922 6657 -3910 6691
rect -3876 6657 -3864 6691
rect -3922 6623 -3864 6657
rect -3922 6589 -3910 6623
rect -3876 6589 -3864 6623
rect -3922 6555 -3864 6589
rect -3922 6521 -3910 6555
rect -3876 6521 -3864 6555
rect -3922 6487 -3864 6521
rect -3922 6453 -3910 6487
rect -3876 6453 -3864 6487
rect -3922 6419 -3864 6453
rect -3922 6385 -3910 6419
rect -3876 6385 -3864 6419
rect -3922 6351 -3864 6385
rect -3922 6317 -3910 6351
rect -3876 6317 -3864 6351
rect -3922 6283 -3864 6317
rect -3922 6249 -3910 6283
rect -3876 6249 -3864 6283
rect -3922 6215 -3864 6249
rect -3922 6181 -3910 6215
rect -3876 6181 -3864 6215
rect -3922 6147 -3864 6181
rect -3922 6113 -3910 6147
rect -3876 6113 -3864 6147
rect -3922 6079 -3864 6113
rect -3922 6045 -3910 6079
rect -3876 6045 -3864 6079
rect -3922 6011 -3864 6045
rect -3922 5977 -3910 6011
rect -3876 5977 -3864 6011
rect -3922 5943 -3864 5977
rect -3922 5909 -3910 5943
rect -3876 5909 -3864 5943
rect -3922 5875 -3864 5909
rect -3922 5841 -3910 5875
rect -3876 5841 -3864 5875
rect -3922 5807 -3864 5841
rect -3922 5773 -3910 5807
rect -3876 5773 -3864 5807
rect -3922 5739 -3864 5773
rect -3922 5705 -3910 5739
rect -3876 5705 -3864 5739
rect -3922 5671 -3864 5705
rect -3922 5637 -3910 5671
rect -3876 5637 -3864 5671
rect -3922 5603 -3864 5637
rect -3922 5569 -3910 5603
rect -3876 5569 -3864 5603
rect -3922 5538 -3864 5569
rect -3664 7507 -3606 7538
rect -3664 7473 -3652 7507
rect -3618 7473 -3606 7507
rect -3664 7439 -3606 7473
rect -3664 7405 -3652 7439
rect -3618 7405 -3606 7439
rect -3664 7371 -3606 7405
rect -3664 7337 -3652 7371
rect -3618 7337 -3606 7371
rect -3664 7303 -3606 7337
rect -3664 7269 -3652 7303
rect -3618 7269 -3606 7303
rect -3664 7235 -3606 7269
rect -3664 7201 -3652 7235
rect -3618 7201 -3606 7235
rect -3664 7167 -3606 7201
rect -3664 7133 -3652 7167
rect -3618 7133 -3606 7167
rect -3664 7099 -3606 7133
rect -3664 7065 -3652 7099
rect -3618 7065 -3606 7099
rect -3664 7031 -3606 7065
rect -3664 6997 -3652 7031
rect -3618 6997 -3606 7031
rect -3664 6963 -3606 6997
rect -3664 6929 -3652 6963
rect -3618 6929 -3606 6963
rect -3664 6895 -3606 6929
rect -3664 6861 -3652 6895
rect -3618 6861 -3606 6895
rect -3664 6827 -3606 6861
rect -3664 6793 -3652 6827
rect -3618 6793 -3606 6827
rect -3664 6759 -3606 6793
rect -3664 6725 -3652 6759
rect -3618 6725 -3606 6759
rect -3664 6691 -3606 6725
rect -3664 6657 -3652 6691
rect -3618 6657 -3606 6691
rect -3664 6623 -3606 6657
rect -3664 6589 -3652 6623
rect -3618 6589 -3606 6623
rect -3664 6555 -3606 6589
rect -3664 6521 -3652 6555
rect -3618 6521 -3606 6555
rect -3664 6487 -3606 6521
rect -3664 6453 -3652 6487
rect -3618 6453 -3606 6487
rect -3664 6419 -3606 6453
rect -3664 6385 -3652 6419
rect -3618 6385 -3606 6419
rect -3664 6351 -3606 6385
rect -3664 6317 -3652 6351
rect -3618 6317 -3606 6351
rect -3664 6283 -3606 6317
rect -3664 6249 -3652 6283
rect -3618 6249 -3606 6283
rect -3664 6215 -3606 6249
rect -3664 6181 -3652 6215
rect -3618 6181 -3606 6215
rect -3664 6147 -3606 6181
rect -3664 6113 -3652 6147
rect -3618 6113 -3606 6147
rect -3664 6079 -3606 6113
rect -3664 6045 -3652 6079
rect -3618 6045 -3606 6079
rect -3664 6011 -3606 6045
rect -3664 5977 -3652 6011
rect -3618 5977 -3606 6011
rect -3664 5943 -3606 5977
rect -3664 5909 -3652 5943
rect -3618 5909 -3606 5943
rect -3664 5875 -3606 5909
rect -3664 5841 -3652 5875
rect -3618 5841 -3606 5875
rect -3664 5807 -3606 5841
rect -3664 5773 -3652 5807
rect -3618 5773 -3606 5807
rect -3664 5739 -3606 5773
rect -3664 5705 -3652 5739
rect -3618 5705 -3606 5739
rect -3664 5671 -3606 5705
rect -3664 5637 -3652 5671
rect -3618 5637 -3606 5671
rect -3664 5603 -3606 5637
rect -3664 5569 -3652 5603
rect -3618 5569 -3606 5603
rect -3664 5538 -3606 5569
rect 17422 7527 17480 7548
rect 17422 7493 17434 7527
rect 17468 7493 17480 7527
rect 17422 7459 17480 7493
rect 17422 7425 17434 7459
rect 17468 7425 17480 7459
rect 17422 7391 17480 7425
rect 17422 7357 17434 7391
rect 17468 7357 17480 7391
rect 17422 7323 17480 7357
rect 17422 7289 17434 7323
rect 17468 7289 17480 7323
rect 17422 7255 17480 7289
rect 17422 7221 17434 7255
rect 17468 7221 17480 7255
rect 17422 7187 17480 7221
rect 17422 7153 17434 7187
rect 17468 7153 17480 7187
rect 17422 7119 17480 7153
rect 17422 7085 17434 7119
rect 17468 7085 17480 7119
rect 17422 7051 17480 7085
rect 17422 7017 17434 7051
rect 17468 7017 17480 7051
rect 17422 6983 17480 7017
rect 17422 6949 17434 6983
rect 17468 6949 17480 6983
rect 17422 6915 17480 6949
rect 17422 6881 17434 6915
rect 17468 6881 17480 6915
rect 17422 6847 17480 6881
rect 17422 6813 17434 6847
rect 17468 6813 17480 6847
rect 17422 6779 17480 6813
rect 17422 6745 17434 6779
rect 17468 6745 17480 6779
rect 17422 6711 17480 6745
rect 17422 6677 17434 6711
rect 17468 6677 17480 6711
rect 17422 6643 17480 6677
rect 17422 6609 17434 6643
rect 17468 6609 17480 6643
rect 17422 6575 17480 6609
rect 17422 6541 17434 6575
rect 17468 6541 17480 6575
rect 17422 6507 17480 6541
rect 17422 6473 17434 6507
rect 17468 6473 17480 6507
rect 17422 6439 17480 6473
rect 17422 6405 17434 6439
rect 17468 6405 17480 6439
rect 17422 6371 17480 6405
rect 17422 6337 17434 6371
rect 17468 6337 17480 6371
rect 17422 6303 17480 6337
rect 17422 6269 17434 6303
rect 17468 6269 17480 6303
rect 17422 6235 17480 6269
rect 17422 6201 17434 6235
rect 17468 6201 17480 6235
rect 17422 6167 17480 6201
rect 17422 6133 17434 6167
rect 17468 6133 17480 6167
rect 17422 6099 17480 6133
rect 17422 6065 17434 6099
rect 17468 6065 17480 6099
rect 17422 6031 17480 6065
rect 17422 5997 17434 6031
rect 17468 5997 17480 6031
rect 17422 5963 17480 5997
rect 17422 5929 17434 5963
rect 17468 5929 17480 5963
rect 17422 5895 17480 5929
rect 17422 5861 17434 5895
rect 17468 5861 17480 5895
rect 17422 5827 17480 5861
rect 17422 5793 17434 5827
rect 17468 5793 17480 5827
rect 17422 5759 17480 5793
rect 17422 5725 17434 5759
rect 17468 5725 17480 5759
rect 17422 5691 17480 5725
rect 17422 5657 17434 5691
rect 17468 5657 17480 5691
rect 17422 5623 17480 5657
rect 17422 5589 17434 5623
rect 17468 5589 17480 5623
rect 17422 5555 17480 5589
rect 17422 5521 17434 5555
rect 17468 5521 17480 5555
rect 17422 5487 17480 5521
rect 17422 5453 17434 5487
rect 17468 5453 17480 5487
rect 17422 5419 17480 5453
rect 17422 5385 17434 5419
rect 17468 5385 17480 5419
rect 17422 5351 17480 5385
rect 17422 5317 17434 5351
rect 17468 5317 17480 5351
rect 17422 5283 17480 5317
rect 17422 5249 17434 5283
rect 17468 5249 17480 5283
rect 17422 5215 17480 5249
rect 17422 5181 17434 5215
rect 17468 5181 17480 5215
rect 17422 5147 17480 5181
rect 17422 5113 17434 5147
rect 17468 5113 17480 5147
rect 17422 5079 17480 5113
rect 17422 5045 17434 5079
rect 17468 5045 17480 5079
rect 17422 5011 17480 5045
rect 17422 4977 17434 5011
rect 17468 4977 17480 5011
rect 17422 4943 17480 4977
rect 17422 4909 17434 4943
rect 17468 4909 17480 4943
rect 17422 4875 17480 4909
rect 17422 4841 17434 4875
rect 17468 4841 17480 4875
rect 17422 4807 17480 4841
rect 17422 4773 17434 4807
rect 17468 4773 17480 4807
rect 17422 4739 17480 4773
rect 17422 4705 17434 4739
rect 17468 4705 17480 4739
rect 17422 4671 17480 4705
rect 17422 4637 17434 4671
rect 17468 4637 17480 4671
rect 17422 4603 17480 4637
rect 17422 4569 17434 4603
rect 17468 4569 17480 4603
rect 17422 4548 17480 4569
rect 18480 7527 18538 7548
rect 18480 7493 18492 7527
rect 18526 7493 18538 7527
rect 18480 7459 18538 7493
rect 18480 7425 18492 7459
rect 18526 7425 18538 7459
rect 18480 7391 18538 7425
rect 18480 7357 18492 7391
rect 18526 7357 18538 7391
rect 18480 7323 18538 7357
rect 18480 7289 18492 7323
rect 18526 7289 18538 7323
rect 18480 7255 18538 7289
rect 18480 7221 18492 7255
rect 18526 7221 18538 7255
rect 18480 7187 18538 7221
rect 18480 7153 18492 7187
rect 18526 7153 18538 7187
rect 18480 7119 18538 7153
rect 18480 7085 18492 7119
rect 18526 7085 18538 7119
rect 18480 7051 18538 7085
rect 18480 7017 18492 7051
rect 18526 7017 18538 7051
rect 18480 6983 18538 7017
rect 18480 6949 18492 6983
rect 18526 6949 18538 6983
rect 18480 6915 18538 6949
rect 18480 6881 18492 6915
rect 18526 6881 18538 6915
rect 18480 6847 18538 6881
rect 18480 6813 18492 6847
rect 18526 6813 18538 6847
rect 18480 6779 18538 6813
rect 18480 6745 18492 6779
rect 18526 6745 18538 6779
rect 18480 6711 18538 6745
rect 18480 6677 18492 6711
rect 18526 6677 18538 6711
rect 18480 6643 18538 6677
rect 18480 6609 18492 6643
rect 18526 6609 18538 6643
rect 18480 6575 18538 6609
rect 18480 6541 18492 6575
rect 18526 6541 18538 6575
rect 18480 6507 18538 6541
rect 18480 6473 18492 6507
rect 18526 6473 18538 6507
rect 18480 6439 18538 6473
rect 18480 6405 18492 6439
rect 18526 6405 18538 6439
rect 18480 6371 18538 6405
rect 18480 6337 18492 6371
rect 18526 6337 18538 6371
rect 18480 6303 18538 6337
rect 18480 6269 18492 6303
rect 18526 6269 18538 6303
rect 18480 6235 18538 6269
rect 18480 6201 18492 6235
rect 18526 6201 18538 6235
rect 18480 6167 18538 6201
rect 18480 6133 18492 6167
rect 18526 6133 18538 6167
rect 18480 6099 18538 6133
rect 18480 6065 18492 6099
rect 18526 6065 18538 6099
rect 18480 6031 18538 6065
rect 18480 5997 18492 6031
rect 18526 5997 18538 6031
rect 18480 5963 18538 5997
rect 18480 5929 18492 5963
rect 18526 5929 18538 5963
rect 18480 5895 18538 5929
rect 18480 5861 18492 5895
rect 18526 5861 18538 5895
rect 18480 5827 18538 5861
rect 18480 5793 18492 5827
rect 18526 5793 18538 5827
rect 18480 5759 18538 5793
rect 18480 5725 18492 5759
rect 18526 5725 18538 5759
rect 18480 5691 18538 5725
rect 18480 5657 18492 5691
rect 18526 5657 18538 5691
rect 18480 5623 18538 5657
rect 18480 5589 18492 5623
rect 18526 5589 18538 5623
rect 18480 5555 18538 5589
rect 18480 5521 18492 5555
rect 18526 5521 18538 5555
rect 18480 5487 18538 5521
rect 18480 5453 18492 5487
rect 18526 5453 18538 5487
rect 18480 5419 18538 5453
rect 18480 5385 18492 5419
rect 18526 5385 18538 5419
rect 18480 5351 18538 5385
rect 18480 5317 18492 5351
rect 18526 5317 18538 5351
rect 18480 5283 18538 5317
rect 18480 5249 18492 5283
rect 18526 5249 18538 5283
rect 18480 5215 18538 5249
rect 18480 5181 18492 5215
rect 18526 5181 18538 5215
rect 18480 5147 18538 5181
rect 18480 5113 18492 5147
rect 18526 5113 18538 5147
rect 18480 5079 18538 5113
rect 18480 5045 18492 5079
rect 18526 5045 18538 5079
rect 18480 5011 18538 5045
rect 18480 4977 18492 5011
rect 18526 4977 18538 5011
rect 18480 4943 18538 4977
rect 18480 4909 18492 4943
rect 18526 4909 18538 4943
rect 18480 4875 18538 4909
rect 18480 4841 18492 4875
rect 18526 4841 18538 4875
rect 18480 4807 18538 4841
rect 18480 4773 18492 4807
rect 18526 4773 18538 4807
rect 18480 4739 18538 4773
rect 18480 4705 18492 4739
rect 18526 4705 18538 4739
rect 18480 4671 18538 4705
rect 18480 4637 18492 4671
rect 18526 4637 18538 4671
rect 18480 4603 18538 4637
rect 18480 4569 18492 4603
rect 18526 4569 18538 4603
rect 18480 4548 18538 4569
rect 18872 7527 18930 7548
rect 18872 7493 18884 7527
rect 18918 7493 18930 7527
rect 18872 7459 18930 7493
rect 18872 7425 18884 7459
rect 18918 7425 18930 7459
rect 18872 7391 18930 7425
rect 18872 7357 18884 7391
rect 18918 7357 18930 7391
rect 18872 7323 18930 7357
rect 18872 7289 18884 7323
rect 18918 7289 18930 7323
rect 18872 7255 18930 7289
rect 18872 7221 18884 7255
rect 18918 7221 18930 7255
rect 18872 7187 18930 7221
rect 18872 7153 18884 7187
rect 18918 7153 18930 7187
rect 18872 7119 18930 7153
rect 18872 7085 18884 7119
rect 18918 7085 18930 7119
rect 18872 7051 18930 7085
rect 18872 7017 18884 7051
rect 18918 7017 18930 7051
rect 18872 6983 18930 7017
rect 18872 6949 18884 6983
rect 18918 6949 18930 6983
rect 18872 6915 18930 6949
rect 18872 6881 18884 6915
rect 18918 6881 18930 6915
rect 18872 6847 18930 6881
rect 18872 6813 18884 6847
rect 18918 6813 18930 6847
rect 18872 6779 18930 6813
rect 18872 6745 18884 6779
rect 18918 6745 18930 6779
rect 18872 6711 18930 6745
rect 18872 6677 18884 6711
rect 18918 6677 18930 6711
rect 18872 6643 18930 6677
rect 18872 6609 18884 6643
rect 18918 6609 18930 6643
rect 18872 6575 18930 6609
rect 18872 6541 18884 6575
rect 18918 6541 18930 6575
rect 18872 6507 18930 6541
rect 18872 6473 18884 6507
rect 18918 6473 18930 6507
rect 18872 6439 18930 6473
rect 18872 6405 18884 6439
rect 18918 6405 18930 6439
rect 18872 6371 18930 6405
rect 18872 6337 18884 6371
rect 18918 6337 18930 6371
rect 18872 6303 18930 6337
rect 18872 6269 18884 6303
rect 18918 6269 18930 6303
rect 18872 6235 18930 6269
rect 18872 6201 18884 6235
rect 18918 6201 18930 6235
rect 18872 6167 18930 6201
rect 18872 6133 18884 6167
rect 18918 6133 18930 6167
rect 18872 6099 18930 6133
rect 18872 6065 18884 6099
rect 18918 6065 18930 6099
rect 18872 6031 18930 6065
rect 18872 5997 18884 6031
rect 18918 5997 18930 6031
rect 18872 5963 18930 5997
rect 18872 5929 18884 5963
rect 18918 5929 18930 5963
rect 18872 5895 18930 5929
rect 18872 5861 18884 5895
rect 18918 5861 18930 5895
rect 18872 5827 18930 5861
rect 18872 5793 18884 5827
rect 18918 5793 18930 5827
rect 18872 5759 18930 5793
rect 18872 5725 18884 5759
rect 18918 5725 18930 5759
rect 18872 5691 18930 5725
rect 18872 5657 18884 5691
rect 18918 5657 18930 5691
rect 18872 5623 18930 5657
rect 18872 5589 18884 5623
rect 18918 5589 18930 5623
rect 18872 5555 18930 5589
rect 18872 5521 18884 5555
rect 18918 5521 18930 5555
rect 18872 5487 18930 5521
rect 18872 5453 18884 5487
rect 18918 5453 18930 5487
rect 18872 5419 18930 5453
rect 18872 5385 18884 5419
rect 18918 5385 18930 5419
rect 18872 5351 18930 5385
rect 18872 5317 18884 5351
rect 18918 5317 18930 5351
rect 18872 5283 18930 5317
rect 18872 5249 18884 5283
rect 18918 5249 18930 5283
rect 18872 5215 18930 5249
rect 18872 5181 18884 5215
rect 18918 5181 18930 5215
rect 18872 5147 18930 5181
rect 18872 5113 18884 5147
rect 18918 5113 18930 5147
rect 18872 5079 18930 5113
rect 18872 5045 18884 5079
rect 18918 5045 18930 5079
rect 18872 5011 18930 5045
rect 18872 4977 18884 5011
rect 18918 4977 18930 5011
rect 18872 4943 18930 4977
rect 18872 4909 18884 4943
rect 18918 4909 18930 4943
rect 18872 4875 18930 4909
rect 18872 4841 18884 4875
rect 18918 4841 18930 4875
rect 18872 4807 18930 4841
rect 18872 4773 18884 4807
rect 18918 4773 18930 4807
rect 18872 4739 18930 4773
rect 18872 4705 18884 4739
rect 18918 4705 18930 4739
rect 18872 4671 18930 4705
rect 18872 4637 18884 4671
rect 18918 4637 18930 4671
rect 18872 4603 18930 4637
rect 18872 4569 18884 4603
rect 18918 4569 18930 4603
rect 18872 4548 18930 4569
rect 19930 7527 19988 7548
rect 19930 7493 19942 7527
rect 19976 7493 19988 7527
rect 19930 7459 19988 7493
rect 19930 7425 19942 7459
rect 19976 7425 19988 7459
rect 19930 7391 19988 7425
rect 19930 7357 19942 7391
rect 19976 7357 19988 7391
rect 19930 7323 19988 7357
rect 19930 7289 19942 7323
rect 19976 7289 19988 7323
rect 19930 7255 19988 7289
rect 19930 7221 19942 7255
rect 19976 7221 19988 7255
rect 19930 7187 19988 7221
rect 19930 7153 19942 7187
rect 19976 7153 19988 7187
rect 19930 7119 19988 7153
rect 19930 7085 19942 7119
rect 19976 7085 19988 7119
rect 19930 7051 19988 7085
rect 19930 7017 19942 7051
rect 19976 7017 19988 7051
rect 19930 6983 19988 7017
rect 19930 6949 19942 6983
rect 19976 6949 19988 6983
rect 19930 6915 19988 6949
rect 19930 6881 19942 6915
rect 19976 6881 19988 6915
rect 19930 6847 19988 6881
rect 19930 6813 19942 6847
rect 19976 6813 19988 6847
rect 19930 6779 19988 6813
rect 19930 6745 19942 6779
rect 19976 6745 19988 6779
rect 19930 6711 19988 6745
rect 19930 6677 19942 6711
rect 19976 6677 19988 6711
rect 19930 6643 19988 6677
rect 19930 6609 19942 6643
rect 19976 6609 19988 6643
rect 19930 6575 19988 6609
rect 19930 6541 19942 6575
rect 19976 6541 19988 6575
rect 19930 6507 19988 6541
rect 19930 6473 19942 6507
rect 19976 6473 19988 6507
rect 19930 6439 19988 6473
rect 19930 6405 19942 6439
rect 19976 6405 19988 6439
rect 19930 6371 19988 6405
rect 19930 6337 19942 6371
rect 19976 6337 19988 6371
rect 19930 6303 19988 6337
rect 19930 6269 19942 6303
rect 19976 6269 19988 6303
rect 19930 6235 19988 6269
rect 19930 6201 19942 6235
rect 19976 6201 19988 6235
rect 19930 6167 19988 6201
rect 19930 6133 19942 6167
rect 19976 6133 19988 6167
rect 19930 6099 19988 6133
rect 19930 6065 19942 6099
rect 19976 6065 19988 6099
rect 19930 6031 19988 6065
rect 19930 5997 19942 6031
rect 19976 5997 19988 6031
rect 19930 5963 19988 5997
rect 19930 5929 19942 5963
rect 19976 5929 19988 5963
rect 19930 5895 19988 5929
rect 19930 5861 19942 5895
rect 19976 5861 19988 5895
rect 19930 5827 19988 5861
rect 19930 5793 19942 5827
rect 19976 5793 19988 5827
rect 19930 5759 19988 5793
rect 19930 5725 19942 5759
rect 19976 5725 19988 5759
rect 19930 5691 19988 5725
rect 19930 5657 19942 5691
rect 19976 5657 19988 5691
rect 19930 5623 19988 5657
rect 19930 5589 19942 5623
rect 19976 5589 19988 5623
rect 19930 5555 19988 5589
rect 19930 5521 19942 5555
rect 19976 5521 19988 5555
rect 19930 5487 19988 5521
rect 19930 5453 19942 5487
rect 19976 5453 19988 5487
rect 19930 5419 19988 5453
rect 19930 5385 19942 5419
rect 19976 5385 19988 5419
rect 19930 5351 19988 5385
rect 19930 5317 19942 5351
rect 19976 5317 19988 5351
rect 19930 5283 19988 5317
rect 19930 5249 19942 5283
rect 19976 5249 19988 5283
rect 19930 5215 19988 5249
rect 19930 5181 19942 5215
rect 19976 5181 19988 5215
rect 19930 5147 19988 5181
rect 19930 5113 19942 5147
rect 19976 5113 19988 5147
rect 19930 5079 19988 5113
rect 19930 5045 19942 5079
rect 19976 5045 19988 5079
rect 19930 5011 19988 5045
rect 19930 4977 19942 5011
rect 19976 4977 19988 5011
rect 19930 4943 19988 4977
rect 19930 4909 19942 4943
rect 19976 4909 19988 4943
rect 19930 4875 19988 4909
rect 19930 4841 19942 4875
rect 19976 4841 19988 4875
rect 19930 4807 19988 4841
rect 19930 4773 19942 4807
rect 19976 4773 19988 4807
rect 19930 4739 19988 4773
rect 19930 4705 19942 4739
rect 19976 4705 19988 4739
rect 19930 4671 19988 4705
rect 19930 4637 19942 4671
rect 19976 4637 19988 4671
rect 19930 4603 19988 4637
rect 19930 4569 19942 4603
rect 19976 4569 19988 4603
rect 19930 4548 19988 4569
rect 38121 15554 38179 15585
rect 38121 15520 38133 15554
rect 38167 15520 38179 15554
rect 38121 15486 38179 15520
rect 38121 15452 38133 15486
rect 38167 15452 38179 15486
rect 38121 15418 38179 15452
rect 38121 15384 38133 15418
rect 38167 15384 38179 15418
rect 38121 15350 38179 15384
rect 38121 15316 38133 15350
rect 38167 15316 38179 15350
rect 38121 15282 38179 15316
rect 38121 15248 38133 15282
rect 38167 15248 38179 15282
rect 38121 15214 38179 15248
rect 38121 15180 38133 15214
rect 38167 15180 38179 15214
rect 38121 15146 38179 15180
rect 38121 15112 38133 15146
rect 38167 15112 38179 15146
rect 38121 15078 38179 15112
rect 38121 15044 38133 15078
rect 38167 15044 38179 15078
rect 38121 15010 38179 15044
rect 38121 14976 38133 15010
rect 38167 14976 38179 15010
rect 38121 14942 38179 14976
rect 38121 14908 38133 14942
rect 38167 14908 38179 14942
rect 38121 14874 38179 14908
rect 38121 14840 38133 14874
rect 38167 14840 38179 14874
rect 38121 14806 38179 14840
rect 38121 14772 38133 14806
rect 38167 14772 38179 14806
rect 38121 14738 38179 14772
rect 38121 14704 38133 14738
rect 38167 14704 38179 14738
rect 38121 14670 38179 14704
rect 38121 14636 38133 14670
rect 38167 14636 38179 14670
rect 38121 14602 38179 14636
rect 38121 14568 38133 14602
rect 38167 14568 38179 14602
rect 38121 14534 38179 14568
rect 38121 14500 38133 14534
rect 38167 14500 38179 14534
rect 38121 14466 38179 14500
rect 38121 14432 38133 14466
rect 38167 14432 38179 14466
rect 38121 14398 38179 14432
rect 38121 14364 38133 14398
rect 38167 14364 38179 14398
rect 38121 14330 38179 14364
rect 38121 14296 38133 14330
rect 38167 14296 38179 14330
rect 38121 14262 38179 14296
rect 38121 14228 38133 14262
rect 38167 14228 38179 14262
rect 38121 14194 38179 14228
rect 38121 14160 38133 14194
rect 38167 14160 38179 14194
rect 38121 14126 38179 14160
rect 38121 14092 38133 14126
rect 38167 14092 38179 14126
rect 38121 14058 38179 14092
rect 38121 14024 38133 14058
rect 38167 14024 38179 14058
rect 38121 13990 38179 14024
rect 38121 13956 38133 13990
rect 38167 13956 38179 13990
rect 38121 13922 38179 13956
rect 38121 13888 38133 13922
rect 38167 13888 38179 13922
rect 38121 13854 38179 13888
rect 38121 13820 38133 13854
rect 38167 13820 38179 13854
rect 38121 13786 38179 13820
rect 38121 13752 38133 13786
rect 38167 13752 38179 13786
rect 38121 13718 38179 13752
rect 38121 13684 38133 13718
rect 38167 13684 38179 13718
rect 38121 13650 38179 13684
rect 38121 13616 38133 13650
rect 38167 13616 38179 13650
rect 38121 13585 38179 13616
rect 38379 15554 38437 15585
rect 38379 15520 38391 15554
rect 38425 15520 38437 15554
rect 38379 15486 38437 15520
rect 38379 15452 38391 15486
rect 38425 15452 38437 15486
rect 38379 15418 38437 15452
rect 38379 15384 38391 15418
rect 38425 15384 38437 15418
rect 38379 15350 38437 15384
rect 38379 15316 38391 15350
rect 38425 15316 38437 15350
rect 38379 15282 38437 15316
rect 38379 15248 38391 15282
rect 38425 15248 38437 15282
rect 38379 15214 38437 15248
rect 38379 15180 38391 15214
rect 38425 15180 38437 15214
rect 38379 15146 38437 15180
rect 38379 15112 38391 15146
rect 38425 15112 38437 15146
rect 38379 15078 38437 15112
rect 38379 15044 38391 15078
rect 38425 15044 38437 15078
rect 38379 15010 38437 15044
rect 38379 14976 38391 15010
rect 38425 14976 38437 15010
rect 38379 14942 38437 14976
rect 38379 14908 38391 14942
rect 38425 14908 38437 14942
rect 38379 14874 38437 14908
rect 38379 14840 38391 14874
rect 38425 14840 38437 14874
rect 38379 14806 38437 14840
rect 38379 14772 38391 14806
rect 38425 14772 38437 14806
rect 38379 14738 38437 14772
rect 38379 14704 38391 14738
rect 38425 14704 38437 14738
rect 38379 14670 38437 14704
rect 38379 14636 38391 14670
rect 38425 14636 38437 14670
rect 38379 14602 38437 14636
rect 38379 14568 38391 14602
rect 38425 14568 38437 14602
rect 38379 14534 38437 14568
rect 38379 14500 38391 14534
rect 38425 14500 38437 14534
rect 38379 14466 38437 14500
rect 38379 14432 38391 14466
rect 38425 14432 38437 14466
rect 38379 14398 38437 14432
rect 38379 14364 38391 14398
rect 38425 14364 38437 14398
rect 38379 14330 38437 14364
rect 38379 14296 38391 14330
rect 38425 14296 38437 14330
rect 38379 14262 38437 14296
rect 38379 14228 38391 14262
rect 38425 14228 38437 14262
rect 38379 14194 38437 14228
rect 38379 14160 38391 14194
rect 38425 14160 38437 14194
rect 38379 14126 38437 14160
rect 38379 14092 38391 14126
rect 38425 14092 38437 14126
rect 38379 14058 38437 14092
rect 38379 14024 38391 14058
rect 38425 14024 38437 14058
rect 38379 13990 38437 14024
rect 38379 13956 38391 13990
rect 38425 13956 38437 13990
rect 38379 13922 38437 13956
rect 38379 13888 38391 13922
rect 38425 13888 38437 13922
rect 38379 13854 38437 13888
rect 38379 13820 38391 13854
rect 38425 13820 38437 13854
rect 38379 13786 38437 13820
rect 38379 13752 38391 13786
rect 38425 13752 38437 13786
rect 38379 13718 38437 13752
rect 38379 13684 38391 13718
rect 38425 13684 38437 13718
rect 38379 13650 38437 13684
rect 38379 13616 38391 13650
rect 38425 13616 38437 13650
rect 38379 13585 38437 13616
rect 38637 15554 38695 15585
rect 38637 15520 38649 15554
rect 38683 15520 38695 15554
rect 38637 15486 38695 15520
rect 38637 15452 38649 15486
rect 38683 15452 38695 15486
rect 38637 15418 38695 15452
rect 38637 15384 38649 15418
rect 38683 15384 38695 15418
rect 38637 15350 38695 15384
rect 38637 15316 38649 15350
rect 38683 15316 38695 15350
rect 38637 15282 38695 15316
rect 38637 15248 38649 15282
rect 38683 15248 38695 15282
rect 38637 15214 38695 15248
rect 38637 15180 38649 15214
rect 38683 15180 38695 15214
rect 38637 15146 38695 15180
rect 38637 15112 38649 15146
rect 38683 15112 38695 15146
rect 38637 15078 38695 15112
rect 38637 15044 38649 15078
rect 38683 15044 38695 15078
rect 38637 15010 38695 15044
rect 38637 14976 38649 15010
rect 38683 14976 38695 15010
rect 38637 14942 38695 14976
rect 38637 14908 38649 14942
rect 38683 14908 38695 14942
rect 38637 14874 38695 14908
rect 38637 14840 38649 14874
rect 38683 14840 38695 14874
rect 38637 14806 38695 14840
rect 38637 14772 38649 14806
rect 38683 14772 38695 14806
rect 38637 14738 38695 14772
rect 38637 14704 38649 14738
rect 38683 14704 38695 14738
rect 38637 14670 38695 14704
rect 38637 14636 38649 14670
rect 38683 14636 38695 14670
rect 38637 14602 38695 14636
rect 38637 14568 38649 14602
rect 38683 14568 38695 14602
rect 38637 14534 38695 14568
rect 38637 14500 38649 14534
rect 38683 14500 38695 14534
rect 38637 14466 38695 14500
rect 38637 14432 38649 14466
rect 38683 14432 38695 14466
rect 38637 14398 38695 14432
rect 38637 14364 38649 14398
rect 38683 14364 38695 14398
rect 38637 14330 38695 14364
rect 38637 14296 38649 14330
rect 38683 14296 38695 14330
rect 38637 14262 38695 14296
rect 38637 14228 38649 14262
rect 38683 14228 38695 14262
rect 38637 14194 38695 14228
rect 38637 14160 38649 14194
rect 38683 14160 38695 14194
rect 38637 14126 38695 14160
rect 38637 14092 38649 14126
rect 38683 14092 38695 14126
rect 38637 14058 38695 14092
rect 38637 14024 38649 14058
rect 38683 14024 38695 14058
rect 38637 13990 38695 14024
rect 38637 13956 38649 13990
rect 38683 13956 38695 13990
rect 38637 13922 38695 13956
rect 38637 13888 38649 13922
rect 38683 13888 38695 13922
rect 38637 13854 38695 13888
rect 38637 13820 38649 13854
rect 38683 13820 38695 13854
rect 38637 13786 38695 13820
rect 38637 13752 38649 13786
rect 38683 13752 38695 13786
rect 38637 13718 38695 13752
rect 38637 13684 38649 13718
rect 38683 13684 38695 13718
rect 38637 13650 38695 13684
rect 38637 13616 38649 13650
rect 38683 13616 38695 13650
rect 38637 13585 38695 13616
rect 38895 15554 38953 15585
rect 38895 15520 38907 15554
rect 38941 15520 38953 15554
rect 38895 15486 38953 15520
rect 38895 15452 38907 15486
rect 38941 15452 38953 15486
rect 38895 15418 38953 15452
rect 38895 15384 38907 15418
rect 38941 15384 38953 15418
rect 38895 15350 38953 15384
rect 38895 15316 38907 15350
rect 38941 15316 38953 15350
rect 38895 15282 38953 15316
rect 38895 15248 38907 15282
rect 38941 15248 38953 15282
rect 38895 15214 38953 15248
rect 38895 15180 38907 15214
rect 38941 15180 38953 15214
rect 38895 15146 38953 15180
rect 38895 15112 38907 15146
rect 38941 15112 38953 15146
rect 38895 15078 38953 15112
rect 38895 15044 38907 15078
rect 38941 15044 38953 15078
rect 38895 15010 38953 15044
rect 38895 14976 38907 15010
rect 38941 14976 38953 15010
rect 38895 14942 38953 14976
rect 38895 14908 38907 14942
rect 38941 14908 38953 14942
rect 38895 14874 38953 14908
rect 38895 14840 38907 14874
rect 38941 14840 38953 14874
rect 38895 14806 38953 14840
rect 38895 14772 38907 14806
rect 38941 14772 38953 14806
rect 38895 14738 38953 14772
rect 38895 14704 38907 14738
rect 38941 14704 38953 14738
rect 38895 14670 38953 14704
rect 38895 14636 38907 14670
rect 38941 14636 38953 14670
rect 38895 14602 38953 14636
rect 38895 14568 38907 14602
rect 38941 14568 38953 14602
rect 38895 14534 38953 14568
rect 38895 14500 38907 14534
rect 38941 14500 38953 14534
rect 38895 14466 38953 14500
rect 38895 14432 38907 14466
rect 38941 14432 38953 14466
rect 38895 14398 38953 14432
rect 38895 14364 38907 14398
rect 38941 14364 38953 14398
rect 38895 14330 38953 14364
rect 38895 14296 38907 14330
rect 38941 14296 38953 14330
rect 38895 14262 38953 14296
rect 38895 14228 38907 14262
rect 38941 14228 38953 14262
rect 38895 14194 38953 14228
rect 38895 14160 38907 14194
rect 38941 14160 38953 14194
rect 38895 14126 38953 14160
rect 38895 14092 38907 14126
rect 38941 14092 38953 14126
rect 38895 14058 38953 14092
rect 38895 14024 38907 14058
rect 38941 14024 38953 14058
rect 38895 13990 38953 14024
rect 38895 13956 38907 13990
rect 38941 13956 38953 13990
rect 38895 13922 38953 13956
rect 38895 13888 38907 13922
rect 38941 13888 38953 13922
rect 38895 13854 38953 13888
rect 38895 13820 38907 13854
rect 38941 13820 38953 13854
rect 38895 13786 38953 13820
rect 38895 13752 38907 13786
rect 38941 13752 38953 13786
rect 38895 13718 38953 13752
rect 38895 13684 38907 13718
rect 38941 13684 38953 13718
rect 38895 13650 38953 13684
rect 38895 13616 38907 13650
rect 38941 13616 38953 13650
rect 38895 13585 38953 13616
rect 39153 15554 39211 15585
rect 39153 15520 39165 15554
rect 39199 15520 39211 15554
rect 39153 15486 39211 15520
rect 39153 15452 39165 15486
rect 39199 15452 39211 15486
rect 39153 15418 39211 15452
rect 39153 15384 39165 15418
rect 39199 15384 39211 15418
rect 39153 15350 39211 15384
rect 39153 15316 39165 15350
rect 39199 15316 39211 15350
rect 39153 15282 39211 15316
rect 39153 15248 39165 15282
rect 39199 15248 39211 15282
rect 39153 15214 39211 15248
rect 39153 15180 39165 15214
rect 39199 15180 39211 15214
rect 39153 15146 39211 15180
rect 39153 15112 39165 15146
rect 39199 15112 39211 15146
rect 39153 15078 39211 15112
rect 39153 15044 39165 15078
rect 39199 15044 39211 15078
rect 39153 15010 39211 15044
rect 39153 14976 39165 15010
rect 39199 14976 39211 15010
rect 39153 14942 39211 14976
rect 39153 14908 39165 14942
rect 39199 14908 39211 14942
rect 39153 14874 39211 14908
rect 39153 14840 39165 14874
rect 39199 14840 39211 14874
rect 39153 14806 39211 14840
rect 39153 14772 39165 14806
rect 39199 14772 39211 14806
rect 39153 14738 39211 14772
rect 39153 14704 39165 14738
rect 39199 14704 39211 14738
rect 39153 14670 39211 14704
rect 39153 14636 39165 14670
rect 39199 14636 39211 14670
rect 39153 14602 39211 14636
rect 39153 14568 39165 14602
rect 39199 14568 39211 14602
rect 39153 14534 39211 14568
rect 39153 14500 39165 14534
rect 39199 14500 39211 14534
rect 39153 14466 39211 14500
rect 39153 14432 39165 14466
rect 39199 14432 39211 14466
rect 39153 14398 39211 14432
rect 39153 14364 39165 14398
rect 39199 14364 39211 14398
rect 39153 14330 39211 14364
rect 39153 14296 39165 14330
rect 39199 14296 39211 14330
rect 39153 14262 39211 14296
rect 39153 14228 39165 14262
rect 39199 14228 39211 14262
rect 39153 14194 39211 14228
rect 39153 14160 39165 14194
rect 39199 14160 39211 14194
rect 39153 14126 39211 14160
rect 39153 14092 39165 14126
rect 39199 14092 39211 14126
rect 39153 14058 39211 14092
rect 39153 14024 39165 14058
rect 39199 14024 39211 14058
rect 39153 13990 39211 14024
rect 39153 13956 39165 13990
rect 39199 13956 39211 13990
rect 39153 13922 39211 13956
rect 39153 13888 39165 13922
rect 39199 13888 39211 13922
rect 39153 13854 39211 13888
rect 39153 13820 39165 13854
rect 39199 13820 39211 13854
rect 39153 13786 39211 13820
rect 39153 13752 39165 13786
rect 39199 13752 39211 13786
rect 39153 13718 39211 13752
rect 39153 13684 39165 13718
rect 39199 13684 39211 13718
rect 39153 13650 39211 13684
rect 39153 13616 39165 13650
rect 39199 13616 39211 13650
rect 39153 13585 39211 13616
rect 39411 15554 39469 15585
rect 39411 15520 39423 15554
rect 39457 15520 39469 15554
rect 39411 15486 39469 15520
rect 39411 15452 39423 15486
rect 39457 15452 39469 15486
rect 39411 15418 39469 15452
rect 39411 15384 39423 15418
rect 39457 15384 39469 15418
rect 39411 15350 39469 15384
rect 39411 15316 39423 15350
rect 39457 15316 39469 15350
rect 39411 15282 39469 15316
rect 39411 15248 39423 15282
rect 39457 15248 39469 15282
rect 39411 15214 39469 15248
rect 39411 15180 39423 15214
rect 39457 15180 39469 15214
rect 39411 15146 39469 15180
rect 39411 15112 39423 15146
rect 39457 15112 39469 15146
rect 39411 15078 39469 15112
rect 39411 15044 39423 15078
rect 39457 15044 39469 15078
rect 39411 15010 39469 15044
rect 39411 14976 39423 15010
rect 39457 14976 39469 15010
rect 39411 14942 39469 14976
rect 39411 14908 39423 14942
rect 39457 14908 39469 14942
rect 39411 14874 39469 14908
rect 39411 14840 39423 14874
rect 39457 14840 39469 14874
rect 39411 14806 39469 14840
rect 39411 14772 39423 14806
rect 39457 14772 39469 14806
rect 39411 14738 39469 14772
rect 39411 14704 39423 14738
rect 39457 14704 39469 14738
rect 39411 14670 39469 14704
rect 39411 14636 39423 14670
rect 39457 14636 39469 14670
rect 39411 14602 39469 14636
rect 39411 14568 39423 14602
rect 39457 14568 39469 14602
rect 39411 14534 39469 14568
rect 39411 14500 39423 14534
rect 39457 14500 39469 14534
rect 39411 14466 39469 14500
rect 39411 14432 39423 14466
rect 39457 14432 39469 14466
rect 39411 14398 39469 14432
rect 39411 14364 39423 14398
rect 39457 14364 39469 14398
rect 39411 14330 39469 14364
rect 39411 14296 39423 14330
rect 39457 14296 39469 14330
rect 39411 14262 39469 14296
rect 39411 14228 39423 14262
rect 39457 14228 39469 14262
rect 39411 14194 39469 14228
rect 39411 14160 39423 14194
rect 39457 14160 39469 14194
rect 39411 14126 39469 14160
rect 39411 14092 39423 14126
rect 39457 14092 39469 14126
rect 39411 14058 39469 14092
rect 39411 14024 39423 14058
rect 39457 14024 39469 14058
rect 39411 13990 39469 14024
rect 39411 13956 39423 13990
rect 39457 13956 39469 13990
rect 39411 13922 39469 13956
rect 39411 13888 39423 13922
rect 39457 13888 39469 13922
rect 39411 13854 39469 13888
rect 39411 13820 39423 13854
rect 39457 13820 39469 13854
rect 39411 13786 39469 13820
rect 39411 13752 39423 13786
rect 39457 13752 39469 13786
rect 39411 13718 39469 13752
rect 39411 13684 39423 13718
rect 39457 13684 39469 13718
rect 39411 13650 39469 13684
rect 39411 13616 39423 13650
rect 39457 13616 39469 13650
rect 39411 13585 39469 13616
rect 39669 15554 39727 15585
rect 39669 15520 39681 15554
rect 39715 15520 39727 15554
rect 39669 15486 39727 15520
rect 39669 15452 39681 15486
rect 39715 15452 39727 15486
rect 39669 15418 39727 15452
rect 39669 15384 39681 15418
rect 39715 15384 39727 15418
rect 39669 15350 39727 15384
rect 39669 15316 39681 15350
rect 39715 15316 39727 15350
rect 39669 15282 39727 15316
rect 39669 15248 39681 15282
rect 39715 15248 39727 15282
rect 39669 15214 39727 15248
rect 39669 15180 39681 15214
rect 39715 15180 39727 15214
rect 39669 15146 39727 15180
rect 39669 15112 39681 15146
rect 39715 15112 39727 15146
rect 39669 15078 39727 15112
rect 39669 15044 39681 15078
rect 39715 15044 39727 15078
rect 39669 15010 39727 15044
rect 39669 14976 39681 15010
rect 39715 14976 39727 15010
rect 39669 14942 39727 14976
rect 39669 14908 39681 14942
rect 39715 14908 39727 14942
rect 39669 14874 39727 14908
rect 39669 14840 39681 14874
rect 39715 14840 39727 14874
rect 39669 14806 39727 14840
rect 39669 14772 39681 14806
rect 39715 14772 39727 14806
rect 39669 14738 39727 14772
rect 39669 14704 39681 14738
rect 39715 14704 39727 14738
rect 39669 14670 39727 14704
rect 39669 14636 39681 14670
rect 39715 14636 39727 14670
rect 39669 14602 39727 14636
rect 39669 14568 39681 14602
rect 39715 14568 39727 14602
rect 39669 14534 39727 14568
rect 39669 14500 39681 14534
rect 39715 14500 39727 14534
rect 39669 14466 39727 14500
rect 39669 14432 39681 14466
rect 39715 14432 39727 14466
rect 39669 14398 39727 14432
rect 39669 14364 39681 14398
rect 39715 14364 39727 14398
rect 39669 14330 39727 14364
rect 39669 14296 39681 14330
rect 39715 14296 39727 14330
rect 39669 14262 39727 14296
rect 39669 14228 39681 14262
rect 39715 14228 39727 14262
rect 39669 14194 39727 14228
rect 39669 14160 39681 14194
rect 39715 14160 39727 14194
rect 39669 14126 39727 14160
rect 39669 14092 39681 14126
rect 39715 14092 39727 14126
rect 39669 14058 39727 14092
rect 39669 14024 39681 14058
rect 39715 14024 39727 14058
rect 39669 13990 39727 14024
rect 39669 13956 39681 13990
rect 39715 13956 39727 13990
rect 39669 13922 39727 13956
rect 39669 13888 39681 13922
rect 39715 13888 39727 13922
rect 39669 13854 39727 13888
rect 39669 13820 39681 13854
rect 39715 13820 39727 13854
rect 39669 13786 39727 13820
rect 39669 13752 39681 13786
rect 39715 13752 39727 13786
rect 39669 13718 39727 13752
rect 39669 13684 39681 13718
rect 39715 13684 39727 13718
rect 39669 13650 39727 13684
rect 39669 13616 39681 13650
rect 39715 13616 39727 13650
rect 39669 13585 39727 13616
rect 39927 15554 39985 15585
rect 39927 15520 39939 15554
rect 39973 15520 39985 15554
rect 39927 15486 39985 15520
rect 39927 15452 39939 15486
rect 39973 15452 39985 15486
rect 39927 15418 39985 15452
rect 39927 15384 39939 15418
rect 39973 15384 39985 15418
rect 39927 15350 39985 15384
rect 39927 15316 39939 15350
rect 39973 15316 39985 15350
rect 39927 15282 39985 15316
rect 39927 15248 39939 15282
rect 39973 15248 39985 15282
rect 39927 15214 39985 15248
rect 39927 15180 39939 15214
rect 39973 15180 39985 15214
rect 39927 15146 39985 15180
rect 39927 15112 39939 15146
rect 39973 15112 39985 15146
rect 39927 15078 39985 15112
rect 39927 15044 39939 15078
rect 39973 15044 39985 15078
rect 39927 15010 39985 15044
rect 39927 14976 39939 15010
rect 39973 14976 39985 15010
rect 39927 14942 39985 14976
rect 39927 14908 39939 14942
rect 39973 14908 39985 14942
rect 39927 14874 39985 14908
rect 39927 14840 39939 14874
rect 39973 14840 39985 14874
rect 39927 14806 39985 14840
rect 39927 14772 39939 14806
rect 39973 14772 39985 14806
rect 39927 14738 39985 14772
rect 39927 14704 39939 14738
rect 39973 14704 39985 14738
rect 39927 14670 39985 14704
rect 39927 14636 39939 14670
rect 39973 14636 39985 14670
rect 39927 14602 39985 14636
rect 39927 14568 39939 14602
rect 39973 14568 39985 14602
rect 39927 14534 39985 14568
rect 39927 14500 39939 14534
rect 39973 14500 39985 14534
rect 39927 14466 39985 14500
rect 39927 14432 39939 14466
rect 39973 14432 39985 14466
rect 39927 14398 39985 14432
rect 39927 14364 39939 14398
rect 39973 14364 39985 14398
rect 39927 14330 39985 14364
rect 39927 14296 39939 14330
rect 39973 14296 39985 14330
rect 39927 14262 39985 14296
rect 39927 14228 39939 14262
rect 39973 14228 39985 14262
rect 39927 14194 39985 14228
rect 39927 14160 39939 14194
rect 39973 14160 39985 14194
rect 39927 14126 39985 14160
rect 39927 14092 39939 14126
rect 39973 14092 39985 14126
rect 39927 14058 39985 14092
rect 39927 14024 39939 14058
rect 39973 14024 39985 14058
rect 39927 13990 39985 14024
rect 39927 13956 39939 13990
rect 39973 13956 39985 13990
rect 39927 13922 39985 13956
rect 39927 13888 39939 13922
rect 39973 13888 39985 13922
rect 39927 13854 39985 13888
rect 39927 13820 39939 13854
rect 39973 13820 39985 13854
rect 39927 13786 39985 13820
rect 39927 13752 39939 13786
rect 39973 13752 39985 13786
rect 39927 13718 39985 13752
rect 39927 13684 39939 13718
rect 39973 13684 39985 13718
rect 39927 13650 39985 13684
rect 39927 13616 39939 13650
rect 39973 13616 39985 13650
rect 39927 13585 39985 13616
rect 40185 15554 40243 15585
rect 40185 15520 40197 15554
rect 40231 15520 40243 15554
rect 40185 15486 40243 15520
rect 40185 15452 40197 15486
rect 40231 15452 40243 15486
rect 40185 15418 40243 15452
rect 40185 15384 40197 15418
rect 40231 15384 40243 15418
rect 40185 15350 40243 15384
rect 40185 15316 40197 15350
rect 40231 15316 40243 15350
rect 40185 15282 40243 15316
rect 40185 15248 40197 15282
rect 40231 15248 40243 15282
rect 40185 15214 40243 15248
rect 40185 15180 40197 15214
rect 40231 15180 40243 15214
rect 40185 15146 40243 15180
rect 40185 15112 40197 15146
rect 40231 15112 40243 15146
rect 40185 15078 40243 15112
rect 40185 15044 40197 15078
rect 40231 15044 40243 15078
rect 40185 15010 40243 15044
rect 40185 14976 40197 15010
rect 40231 14976 40243 15010
rect 40185 14942 40243 14976
rect 40185 14908 40197 14942
rect 40231 14908 40243 14942
rect 40185 14874 40243 14908
rect 40185 14840 40197 14874
rect 40231 14840 40243 14874
rect 40185 14806 40243 14840
rect 40185 14772 40197 14806
rect 40231 14772 40243 14806
rect 40185 14738 40243 14772
rect 40185 14704 40197 14738
rect 40231 14704 40243 14738
rect 40185 14670 40243 14704
rect 40185 14636 40197 14670
rect 40231 14636 40243 14670
rect 40185 14602 40243 14636
rect 40185 14568 40197 14602
rect 40231 14568 40243 14602
rect 40185 14534 40243 14568
rect 40185 14500 40197 14534
rect 40231 14500 40243 14534
rect 40185 14466 40243 14500
rect 40185 14432 40197 14466
rect 40231 14432 40243 14466
rect 40185 14398 40243 14432
rect 40185 14364 40197 14398
rect 40231 14364 40243 14398
rect 40185 14330 40243 14364
rect 40185 14296 40197 14330
rect 40231 14296 40243 14330
rect 40185 14262 40243 14296
rect 40185 14228 40197 14262
rect 40231 14228 40243 14262
rect 40185 14194 40243 14228
rect 40185 14160 40197 14194
rect 40231 14160 40243 14194
rect 40185 14126 40243 14160
rect 40185 14092 40197 14126
rect 40231 14092 40243 14126
rect 40185 14058 40243 14092
rect 40185 14024 40197 14058
rect 40231 14024 40243 14058
rect 40185 13990 40243 14024
rect 40185 13956 40197 13990
rect 40231 13956 40243 13990
rect 40185 13922 40243 13956
rect 40185 13888 40197 13922
rect 40231 13888 40243 13922
rect 40185 13854 40243 13888
rect 40185 13820 40197 13854
rect 40231 13820 40243 13854
rect 40185 13786 40243 13820
rect 40185 13752 40197 13786
rect 40231 13752 40243 13786
rect 40185 13718 40243 13752
rect 40185 13684 40197 13718
rect 40231 13684 40243 13718
rect 40185 13650 40243 13684
rect 40185 13616 40197 13650
rect 40231 13616 40243 13650
rect 40185 13585 40243 13616
rect 40443 15554 40501 15585
rect 40443 15520 40455 15554
rect 40489 15520 40501 15554
rect 40443 15486 40501 15520
rect 40443 15452 40455 15486
rect 40489 15452 40501 15486
rect 40443 15418 40501 15452
rect 40443 15384 40455 15418
rect 40489 15384 40501 15418
rect 40443 15350 40501 15384
rect 40443 15316 40455 15350
rect 40489 15316 40501 15350
rect 40443 15282 40501 15316
rect 40443 15248 40455 15282
rect 40489 15248 40501 15282
rect 40443 15214 40501 15248
rect 40443 15180 40455 15214
rect 40489 15180 40501 15214
rect 40443 15146 40501 15180
rect 40443 15112 40455 15146
rect 40489 15112 40501 15146
rect 40443 15078 40501 15112
rect 40443 15044 40455 15078
rect 40489 15044 40501 15078
rect 40443 15010 40501 15044
rect 40443 14976 40455 15010
rect 40489 14976 40501 15010
rect 40443 14942 40501 14976
rect 40443 14908 40455 14942
rect 40489 14908 40501 14942
rect 40443 14874 40501 14908
rect 40443 14840 40455 14874
rect 40489 14840 40501 14874
rect 40443 14806 40501 14840
rect 40443 14772 40455 14806
rect 40489 14772 40501 14806
rect 40443 14738 40501 14772
rect 40443 14704 40455 14738
rect 40489 14704 40501 14738
rect 40443 14670 40501 14704
rect 40443 14636 40455 14670
rect 40489 14636 40501 14670
rect 40443 14602 40501 14636
rect 40443 14568 40455 14602
rect 40489 14568 40501 14602
rect 40443 14534 40501 14568
rect 40443 14500 40455 14534
rect 40489 14500 40501 14534
rect 40443 14466 40501 14500
rect 40443 14432 40455 14466
rect 40489 14432 40501 14466
rect 40443 14398 40501 14432
rect 40443 14364 40455 14398
rect 40489 14364 40501 14398
rect 40443 14330 40501 14364
rect 40443 14296 40455 14330
rect 40489 14296 40501 14330
rect 40443 14262 40501 14296
rect 40443 14228 40455 14262
rect 40489 14228 40501 14262
rect 40443 14194 40501 14228
rect 40443 14160 40455 14194
rect 40489 14160 40501 14194
rect 40443 14126 40501 14160
rect 40443 14092 40455 14126
rect 40489 14092 40501 14126
rect 40443 14058 40501 14092
rect 40443 14024 40455 14058
rect 40489 14024 40501 14058
rect 40443 13990 40501 14024
rect 40443 13956 40455 13990
rect 40489 13956 40501 13990
rect 40443 13922 40501 13956
rect 40443 13888 40455 13922
rect 40489 13888 40501 13922
rect 40443 13854 40501 13888
rect 40443 13820 40455 13854
rect 40489 13820 40501 13854
rect 40443 13786 40501 13820
rect 40443 13752 40455 13786
rect 40489 13752 40501 13786
rect 40443 13718 40501 13752
rect 40443 13684 40455 13718
rect 40489 13684 40501 13718
rect 40443 13650 40501 13684
rect 40443 13616 40455 13650
rect 40489 13616 40501 13650
rect 40443 13585 40501 13616
rect 40701 15554 40759 15585
rect 40701 15520 40713 15554
rect 40747 15520 40759 15554
rect 40701 15486 40759 15520
rect 40701 15452 40713 15486
rect 40747 15452 40759 15486
rect 40701 15418 40759 15452
rect 40701 15384 40713 15418
rect 40747 15384 40759 15418
rect 40701 15350 40759 15384
rect 40701 15316 40713 15350
rect 40747 15316 40759 15350
rect 40701 15282 40759 15316
rect 40701 15248 40713 15282
rect 40747 15248 40759 15282
rect 40701 15214 40759 15248
rect 40701 15180 40713 15214
rect 40747 15180 40759 15214
rect 40701 15146 40759 15180
rect 40701 15112 40713 15146
rect 40747 15112 40759 15146
rect 40701 15078 40759 15112
rect 40701 15044 40713 15078
rect 40747 15044 40759 15078
rect 40701 15010 40759 15044
rect 40701 14976 40713 15010
rect 40747 14976 40759 15010
rect 40701 14942 40759 14976
rect 40701 14908 40713 14942
rect 40747 14908 40759 14942
rect 40701 14874 40759 14908
rect 40701 14840 40713 14874
rect 40747 14840 40759 14874
rect 40701 14806 40759 14840
rect 40701 14772 40713 14806
rect 40747 14772 40759 14806
rect 40701 14738 40759 14772
rect 40701 14704 40713 14738
rect 40747 14704 40759 14738
rect 40701 14670 40759 14704
rect 40701 14636 40713 14670
rect 40747 14636 40759 14670
rect 40701 14602 40759 14636
rect 40701 14568 40713 14602
rect 40747 14568 40759 14602
rect 40701 14534 40759 14568
rect 40701 14500 40713 14534
rect 40747 14500 40759 14534
rect 40701 14466 40759 14500
rect 40701 14432 40713 14466
rect 40747 14432 40759 14466
rect 40701 14398 40759 14432
rect 40701 14364 40713 14398
rect 40747 14364 40759 14398
rect 40701 14330 40759 14364
rect 40701 14296 40713 14330
rect 40747 14296 40759 14330
rect 40701 14262 40759 14296
rect 40701 14228 40713 14262
rect 40747 14228 40759 14262
rect 40701 14194 40759 14228
rect 40701 14160 40713 14194
rect 40747 14160 40759 14194
rect 40701 14126 40759 14160
rect 40701 14092 40713 14126
rect 40747 14092 40759 14126
rect 40701 14058 40759 14092
rect 40701 14024 40713 14058
rect 40747 14024 40759 14058
rect 40701 13990 40759 14024
rect 40701 13956 40713 13990
rect 40747 13956 40759 13990
rect 40701 13922 40759 13956
rect 40701 13888 40713 13922
rect 40747 13888 40759 13922
rect 40701 13854 40759 13888
rect 40701 13820 40713 13854
rect 40747 13820 40759 13854
rect 40701 13786 40759 13820
rect 40701 13752 40713 13786
rect 40747 13752 40759 13786
rect 40701 13718 40759 13752
rect 40701 13684 40713 13718
rect 40747 13684 40759 13718
rect 40701 13650 40759 13684
rect 40701 13616 40713 13650
rect 40747 13616 40759 13650
rect 40701 13585 40759 13616
rect 23130 11816 24130 11828
rect 23130 11782 23171 11816
rect 23205 11782 23239 11816
rect 23273 11782 23307 11816
rect 23341 11782 23375 11816
rect 23409 11782 23443 11816
rect 23477 11782 23511 11816
rect 23545 11782 23579 11816
rect 23613 11782 23647 11816
rect 23681 11782 23715 11816
rect 23749 11782 23783 11816
rect 23817 11782 23851 11816
rect 23885 11782 23919 11816
rect 23953 11782 23987 11816
rect 24021 11782 24055 11816
rect 24089 11782 24130 11816
rect 23130 11770 24130 11782
rect 23130 10758 24130 10770
rect 23130 10724 23171 10758
rect 23205 10724 23239 10758
rect 23273 10724 23307 10758
rect 23341 10724 23375 10758
rect 23409 10724 23443 10758
rect 23477 10724 23511 10758
rect 23545 10724 23579 10758
rect 23613 10724 23647 10758
rect 23681 10724 23715 10758
rect 23749 10724 23783 10758
rect 23817 10724 23851 10758
rect 23885 10724 23919 10758
rect 23953 10724 23987 10758
rect 24021 10724 24055 10758
rect 24089 10724 24130 10758
rect 23130 10712 24130 10724
rect 23610 7880 24610 7892
rect 23610 7846 23651 7880
rect 23685 7846 23719 7880
rect 23753 7846 23787 7880
rect 23821 7846 23855 7880
rect 23889 7846 23923 7880
rect 23957 7846 23991 7880
rect 24025 7846 24059 7880
rect 24093 7846 24127 7880
rect 24161 7846 24195 7880
rect 24229 7846 24263 7880
rect 24297 7846 24331 7880
rect 24365 7846 24399 7880
rect 24433 7846 24467 7880
rect 24501 7846 24535 7880
rect 24569 7846 24610 7880
rect 23610 7834 24610 7846
rect 23610 6822 24610 6834
rect 23610 6788 23651 6822
rect 23685 6788 23719 6822
rect 23753 6788 23787 6822
rect 23821 6788 23855 6822
rect 23889 6788 23923 6822
rect 23957 6788 23991 6822
rect 24025 6788 24059 6822
rect 24093 6788 24127 6822
rect 24161 6788 24195 6822
rect 24229 6788 24263 6822
rect 24297 6788 24331 6822
rect 24365 6788 24399 6822
rect 24433 6788 24467 6822
rect 24501 6788 24535 6822
rect 24569 6788 24610 6822
rect 23610 6776 24610 6788
rect 23610 5764 24610 5776
rect 23610 5730 23651 5764
rect 23685 5730 23719 5764
rect 23753 5730 23787 5764
rect 23821 5730 23855 5764
rect 23889 5730 23923 5764
rect 23957 5730 23991 5764
rect 24025 5730 24059 5764
rect 24093 5730 24127 5764
rect 24161 5730 24195 5764
rect 24229 5730 24263 5764
rect 24297 5730 24331 5764
rect 24365 5730 24399 5764
rect 24433 5730 24467 5764
rect 24501 5730 24535 5764
rect 24569 5730 24610 5764
rect 23610 5718 24610 5730
rect 23610 4706 24610 4718
rect 23610 4672 23651 4706
rect 23685 4672 23719 4706
rect 23753 4672 23787 4706
rect 23821 4672 23855 4706
rect 23889 4672 23923 4706
rect 23957 4672 23991 4706
rect 24025 4672 24059 4706
rect 24093 4672 24127 4706
rect 24161 4672 24195 4706
rect 24229 4672 24263 4706
rect 24297 4672 24331 4706
rect 24365 4672 24399 4706
rect 24433 4672 24467 4706
rect 24501 4672 24535 4706
rect 24569 4672 24610 4706
rect 23610 4660 24610 4672
rect 23610 3648 24610 3660
rect 23610 3614 23651 3648
rect 23685 3614 23719 3648
rect 23753 3614 23787 3648
rect 23821 3614 23855 3648
rect 23889 3614 23923 3648
rect 23957 3614 23991 3648
rect 24025 3614 24059 3648
rect 24093 3614 24127 3648
rect 24161 3614 24195 3648
rect 24229 3614 24263 3648
rect 24297 3614 24331 3648
rect 24365 3614 24399 3648
rect 24433 3614 24467 3648
rect 24501 3614 24535 3648
rect 24569 3614 24610 3648
rect 23610 3602 24610 3614
rect 25110 7880 26110 7892
rect 25110 7846 25151 7880
rect 25185 7846 25219 7880
rect 25253 7846 25287 7880
rect 25321 7846 25355 7880
rect 25389 7846 25423 7880
rect 25457 7846 25491 7880
rect 25525 7846 25559 7880
rect 25593 7846 25627 7880
rect 25661 7846 25695 7880
rect 25729 7846 25763 7880
rect 25797 7846 25831 7880
rect 25865 7846 25899 7880
rect 25933 7846 25967 7880
rect 26001 7846 26035 7880
rect 26069 7846 26110 7880
rect 25110 7834 26110 7846
rect 25110 6822 26110 6834
rect 25110 6788 25151 6822
rect 25185 6788 25219 6822
rect 25253 6788 25287 6822
rect 25321 6788 25355 6822
rect 25389 6788 25423 6822
rect 25457 6788 25491 6822
rect 25525 6788 25559 6822
rect 25593 6788 25627 6822
rect 25661 6788 25695 6822
rect 25729 6788 25763 6822
rect 25797 6788 25831 6822
rect 25865 6788 25899 6822
rect 25933 6788 25967 6822
rect 26001 6788 26035 6822
rect 26069 6788 26110 6822
rect 25110 6776 26110 6788
rect 25110 5764 26110 5776
rect 25110 5730 25151 5764
rect 25185 5730 25219 5764
rect 25253 5730 25287 5764
rect 25321 5730 25355 5764
rect 25389 5730 25423 5764
rect 25457 5730 25491 5764
rect 25525 5730 25559 5764
rect 25593 5730 25627 5764
rect 25661 5730 25695 5764
rect 25729 5730 25763 5764
rect 25797 5730 25831 5764
rect 25865 5730 25899 5764
rect 25933 5730 25967 5764
rect 26001 5730 26035 5764
rect 26069 5730 26110 5764
rect 25110 5718 26110 5730
rect 25110 4706 26110 4718
rect 25110 4672 25151 4706
rect 25185 4672 25219 4706
rect 25253 4672 25287 4706
rect 25321 4672 25355 4706
rect 25389 4672 25423 4706
rect 25457 4672 25491 4706
rect 25525 4672 25559 4706
rect 25593 4672 25627 4706
rect 25661 4672 25695 4706
rect 25729 4672 25763 4706
rect 25797 4672 25831 4706
rect 25865 4672 25899 4706
rect 25933 4672 25967 4706
rect 26001 4672 26035 4706
rect 26069 4672 26110 4706
rect 25110 4660 26110 4672
rect 25110 3648 26110 3660
rect 25110 3614 25151 3648
rect 25185 3614 25219 3648
rect 25253 3614 25287 3648
rect 25321 3614 25355 3648
rect 25389 3614 25423 3648
rect 25457 3614 25491 3648
rect 25525 3614 25559 3648
rect 25593 3614 25627 3648
rect 25661 3614 25695 3648
rect 25729 3614 25763 3648
rect 25797 3614 25831 3648
rect 25865 3614 25899 3648
rect 25933 3614 25967 3648
rect 26001 3614 26035 3648
rect 26069 3614 26110 3648
rect 25110 3602 26110 3614
rect 36765 11873 36823 11914
rect 36765 11839 36777 11873
rect 36811 11839 36823 11873
rect 36765 11805 36823 11839
rect 36765 11771 36777 11805
rect 36811 11771 36823 11805
rect 36765 11737 36823 11771
rect 36765 11703 36777 11737
rect 36811 11703 36823 11737
rect 36765 11669 36823 11703
rect 36765 11635 36777 11669
rect 36811 11635 36823 11669
rect 36765 11601 36823 11635
rect 36765 11567 36777 11601
rect 36811 11567 36823 11601
rect 36765 11533 36823 11567
rect 36765 11499 36777 11533
rect 36811 11499 36823 11533
rect 36765 11465 36823 11499
rect 36765 11431 36777 11465
rect 36811 11431 36823 11465
rect 36765 11397 36823 11431
rect 36765 11363 36777 11397
rect 36811 11363 36823 11397
rect 36765 11329 36823 11363
rect 36765 11295 36777 11329
rect 36811 11295 36823 11329
rect 36765 11261 36823 11295
rect 36765 11227 36777 11261
rect 36811 11227 36823 11261
rect 36765 11193 36823 11227
rect 36765 11159 36777 11193
rect 36811 11159 36823 11193
rect 36765 11125 36823 11159
rect 36765 11091 36777 11125
rect 36811 11091 36823 11125
rect 36765 11057 36823 11091
rect 36765 11023 36777 11057
rect 36811 11023 36823 11057
rect 36765 10989 36823 11023
rect 36765 10955 36777 10989
rect 36811 10955 36823 10989
rect 36765 10914 36823 10955
rect 37023 11873 37081 11914
rect 37023 11839 37035 11873
rect 37069 11839 37081 11873
rect 37023 11805 37081 11839
rect 37023 11771 37035 11805
rect 37069 11771 37081 11805
rect 37023 11737 37081 11771
rect 37023 11703 37035 11737
rect 37069 11703 37081 11737
rect 37023 11669 37081 11703
rect 37023 11635 37035 11669
rect 37069 11635 37081 11669
rect 37023 11601 37081 11635
rect 37023 11567 37035 11601
rect 37069 11567 37081 11601
rect 37023 11533 37081 11567
rect 37023 11499 37035 11533
rect 37069 11499 37081 11533
rect 37023 11465 37081 11499
rect 37023 11431 37035 11465
rect 37069 11431 37081 11465
rect 37023 11397 37081 11431
rect 37023 11363 37035 11397
rect 37069 11363 37081 11397
rect 37023 11329 37081 11363
rect 37023 11295 37035 11329
rect 37069 11295 37081 11329
rect 37023 11261 37081 11295
rect 37023 11227 37035 11261
rect 37069 11227 37081 11261
rect 37023 11193 37081 11227
rect 37023 11159 37035 11193
rect 37069 11159 37081 11193
rect 37023 11125 37081 11159
rect 37023 11091 37035 11125
rect 37069 11091 37081 11125
rect 37023 11057 37081 11091
rect 37023 11023 37035 11057
rect 37069 11023 37081 11057
rect 37023 10989 37081 11023
rect 37023 10955 37035 10989
rect 37069 10955 37081 10989
rect 37023 10914 37081 10955
rect 37281 11873 37339 11914
rect 37281 11839 37293 11873
rect 37327 11839 37339 11873
rect 37281 11805 37339 11839
rect 37281 11771 37293 11805
rect 37327 11771 37339 11805
rect 37281 11737 37339 11771
rect 37281 11703 37293 11737
rect 37327 11703 37339 11737
rect 37281 11669 37339 11703
rect 37281 11635 37293 11669
rect 37327 11635 37339 11669
rect 37281 11601 37339 11635
rect 37281 11567 37293 11601
rect 37327 11567 37339 11601
rect 37281 11533 37339 11567
rect 37281 11499 37293 11533
rect 37327 11499 37339 11533
rect 37281 11465 37339 11499
rect 37281 11431 37293 11465
rect 37327 11431 37339 11465
rect 37281 11397 37339 11431
rect 37281 11363 37293 11397
rect 37327 11363 37339 11397
rect 37281 11329 37339 11363
rect 37281 11295 37293 11329
rect 37327 11295 37339 11329
rect 37281 11261 37339 11295
rect 37281 11227 37293 11261
rect 37327 11227 37339 11261
rect 37281 11193 37339 11227
rect 37281 11159 37293 11193
rect 37327 11159 37339 11193
rect 37281 11125 37339 11159
rect 37281 11091 37293 11125
rect 37327 11091 37339 11125
rect 37281 11057 37339 11091
rect 37281 11023 37293 11057
rect 37327 11023 37339 11057
rect 37281 10989 37339 11023
rect 37281 10955 37293 10989
rect 37327 10955 37339 10989
rect 37281 10914 37339 10955
rect 37539 11873 37597 11914
rect 37539 11839 37551 11873
rect 37585 11839 37597 11873
rect 37539 11805 37597 11839
rect 37539 11771 37551 11805
rect 37585 11771 37597 11805
rect 37539 11737 37597 11771
rect 37539 11703 37551 11737
rect 37585 11703 37597 11737
rect 37539 11669 37597 11703
rect 37539 11635 37551 11669
rect 37585 11635 37597 11669
rect 37539 11601 37597 11635
rect 37539 11567 37551 11601
rect 37585 11567 37597 11601
rect 37539 11533 37597 11567
rect 37539 11499 37551 11533
rect 37585 11499 37597 11533
rect 37539 11465 37597 11499
rect 37539 11431 37551 11465
rect 37585 11431 37597 11465
rect 37539 11397 37597 11431
rect 37539 11363 37551 11397
rect 37585 11363 37597 11397
rect 37539 11329 37597 11363
rect 37539 11295 37551 11329
rect 37585 11295 37597 11329
rect 37539 11261 37597 11295
rect 37539 11227 37551 11261
rect 37585 11227 37597 11261
rect 37539 11193 37597 11227
rect 37539 11159 37551 11193
rect 37585 11159 37597 11193
rect 37539 11125 37597 11159
rect 37539 11091 37551 11125
rect 37585 11091 37597 11125
rect 37539 11057 37597 11091
rect 37539 11023 37551 11057
rect 37585 11023 37597 11057
rect 37539 10989 37597 11023
rect 37539 10955 37551 10989
rect 37585 10955 37597 10989
rect 37539 10914 37597 10955
rect 37797 11873 37855 11914
rect 37797 11839 37809 11873
rect 37843 11839 37855 11873
rect 37797 11805 37855 11839
rect 37797 11771 37809 11805
rect 37843 11771 37855 11805
rect 37797 11737 37855 11771
rect 37797 11703 37809 11737
rect 37843 11703 37855 11737
rect 37797 11669 37855 11703
rect 37797 11635 37809 11669
rect 37843 11635 37855 11669
rect 37797 11601 37855 11635
rect 37797 11567 37809 11601
rect 37843 11567 37855 11601
rect 37797 11533 37855 11567
rect 37797 11499 37809 11533
rect 37843 11499 37855 11533
rect 37797 11465 37855 11499
rect 37797 11431 37809 11465
rect 37843 11431 37855 11465
rect 37797 11397 37855 11431
rect 37797 11363 37809 11397
rect 37843 11363 37855 11397
rect 37797 11329 37855 11363
rect 37797 11295 37809 11329
rect 37843 11295 37855 11329
rect 37797 11261 37855 11295
rect 37797 11227 37809 11261
rect 37843 11227 37855 11261
rect 37797 11193 37855 11227
rect 37797 11159 37809 11193
rect 37843 11159 37855 11193
rect 37797 11125 37855 11159
rect 37797 11091 37809 11125
rect 37843 11091 37855 11125
rect 37797 11057 37855 11091
rect 37797 11023 37809 11057
rect 37843 11023 37855 11057
rect 37797 10989 37855 11023
rect 37797 10955 37809 10989
rect 37843 10955 37855 10989
rect 37797 10914 37855 10955
rect 38055 11873 38113 11914
rect 38055 11839 38067 11873
rect 38101 11839 38113 11873
rect 38055 11805 38113 11839
rect 38055 11771 38067 11805
rect 38101 11771 38113 11805
rect 38055 11737 38113 11771
rect 38055 11703 38067 11737
rect 38101 11703 38113 11737
rect 38055 11669 38113 11703
rect 38055 11635 38067 11669
rect 38101 11635 38113 11669
rect 38055 11601 38113 11635
rect 38055 11567 38067 11601
rect 38101 11567 38113 11601
rect 38055 11533 38113 11567
rect 38055 11499 38067 11533
rect 38101 11499 38113 11533
rect 38055 11465 38113 11499
rect 38055 11431 38067 11465
rect 38101 11431 38113 11465
rect 38055 11397 38113 11431
rect 38055 11363 38067 11397
rect 38101 11363 38113 11397
rect 38055 11329 38113 11363
rect 38055 11295 38067 11329
rect 38101 11295 38113 11329
rect 38055 11261 38113 11295
rect 38055 11227 38067 11261
rect 38101 11227 38113 11261
rect 38055 11193 38113 11227
rect 38055 11159 38067 11193
rect 38101 11159 38113 11193
rect 38055 11125 38113 11159
rect 38055 11091 38067 11125
rect 38101 11091 38113 11125
rect 38055 11057 38113 11091
rect 38055 11023 38067 11057
rect 38101 11023 38113 11057
rect 38055 10989 38113 11023
rect 38055 10955 38067 10989
rect 38101 10955 38113 10989
rect 38055 10914 38113 10955
rect 38313 11873 38371 11914
rect 38313 11839 38325 11873
rect 38359 11839 38371 11873
rect 38313 11805 38371 11839
rect 38313 11771 38325 11805
rect 38359 11771 38371 11805
rect 38313 11737 38371 11771
rect 38313 11703 38325 11737
rect 38359 11703 38371 11737
rect 38313 11669 38371 11703
rect 38313 11635 38325 11669
rect 38359 11635 38371 11669
rect 38313 11601 38371 11635
rect 38313 11567 38325 11601
rect 38359 11567 38371 11601
rect 38313 11533 38371 11567
rect 38313 11499 38325 11533
rect 38359 11499 38371 11533
rect 38313 11465 38371 11499
rect 38313 11431 38325 11465
rect 38359 11431 38371 11465
rect 38313 11397 38371 11431
rect 38313 11363 38325 11397
rect 38359 11363 38371 11397
rect 38313 11329 38371 11363
rect 38313 11295 38325 11329
rect 38359 11295 38371 11329
rect 38313 11261 38371 11295
rect 38313 11227 38325 11261
rect 38359 11227 38371 11261
rect 38313 11193 38371 11227
rect 38313 11159 38325 11193
rect 38359 11159 38371 11193
rect 38313 11125 38371 11159
rect 38313 11091 38325 11125
rect 38359 11091 38371 11125
rect 38313 11057 38371 11091
rect 38313 11023 38325 11057
rect 38359 11023 38371 11057
rect 38313 10989 38371 11023
rect 38313 10955 38325 10989
rect 38359 10955 38371 10989
rect 38313 10914 38371 10955
rect 38571 11873 38629 11914
rect 38571 11839 38583 11873
rect 38617 11839 38629 11873
rect 38571 11805 38629 11839
rect 38571 11771 38583 11805
rect 38617 11771 38629 11805
rect 38571 11737 38629 11771
rect 38571 11703 38583 11737
rect 38617 11703 38629 11737
rect 38571 11669 38629 11703
rect 38571 11635 38583 11669
rect 38617 11635 38629 11669
rect 38571 11601 38629 11635
rect 38571 11567 38583 11601
rect 38617 11567 38629 11601
rect 38571 11533 38629 11567
rect 38571 11499 38583 11533
rect 38617 11499 38629 11533
rect 38571 11465 38629 11499
rect 38571 11431 38583 11465
rect 38617 11431 38629 11465
rect 38571 11397 38629 11431
rect 38571 11363 38583 11397
rect 38617 11363 38629 11397
rect 38571 11329 38629 11363
rect 38571 11295 38583 11329
rect 38617 11295 38629 11329
rect 38571 11261 38629 11295
rect 38571 11227 38583 11261
rect 38617 11227 38629 11261
rect 38571 11193 38629 11227
rect 38571 11159 38583 11193
rect 38617 11159 38629 11193
rect 38571 11125 38629 11159
rect 38571 11091 38583 11125
rect 38617 11091 38629 11125
rect 38571 11057 38629 11091
rect 38571 11023 38583 11057
rect 38617 11023 38629 11057
rect 38571 10989 38629 11023
rect 38571 10955 38583 10989
rect 38617 10955 38629 10989
rect 38571 10914 38629 10955
rect 38829 11873 38887 11914
rect 38829 11839 38841 11873
rect 38875 11839 38887 11873
rect 38829 11805 38887 11839
rect 38829 11771 38841 11805
rect 38875 11771 38887 11805
rect 38829 11737 38887 11771
rect 38829 11703 38841 11737
rect 38875 11703 38887 11737
rect 38829 11669 38887 11703
rect 38829 11635 38841 11669
rect 38875 11635 38887 11669
rect 38829 11601 38887 11635
rect 38829 11567 38841 11601
rect 38875 11567 38887 11601
rect 38829 11533 38887 11567
rect 38829 11499 38841 11533
rect 38875 11499 38887 11533
rect 38829 11465 38887 11499
rect 38829 11431 38841 11465
rect 38875 11431 38887 11465
rect 38829 11397 38887 11431
rect 38829 11363 38841 11397
rect 38875 11363 38887 11397
rect 38829 11329 38887 11363
rect 38829 11295 38841 11329
rect 38875 11295 38887 11329
rect 38829 11261 38887 11295
rect 38829 11227 38841 11261
rect 38875 11227 38887 11261
rect 38829 11193 38887 11227
rect 38829 11159 38841 11193
rect 38875 11159 38887 11193
rect 38829 11125 38887 11159
rect 38829 11091 38841 11125
rect 38875 11091 38887 11125
rect 38829 11057 38887 11091
rect 38829 11023 38841 11057
rect 38875 11023 38887 11057
rect 38829 10989 38887 11023
rect 38829 10955 38841 10989
rect 38875 10955 38887 10989
rect 38829 10914 38887 10955
rect 39087 11873 39145 11914
rect 39087 11839 39099 11873
rect 39133 11839 39145 11873
rect 39087 11805 39145 11839
rect 39087 11771 39099 11805
rect 39133 11771 39145 11805
rect 39087 11737 39145 11771
rect 39087 11703 39099 11737
rect 39133 11703 39145 11737
rect 39087 11669 39145 11703
rect 39087 11635 39099 11669
rect 39133 11635 39145 11669
rect 39087 11601 39145 11635
rect 39087 11567 39099 11601
rect 39133 11567 39145 11601
rect 39087 11533 39145 11567
rect 39087 11499 39099 11533
rect 39133 11499 39145 11533
rect 39087 11465 39145 11499
rect 39087 11431 39099 11465
rect 39133 11431 39145 11465
rect 39087 11397 39145 11431
rect 39087 11363 39099 11397
rect 39133 11363 39145 11397
rect 39087 11329 39145 11363
rect 39087 11295 39099 11329
rect 39133 11295 39145 11329
rect 39087 11261 39145 11295
rect 39087 11227 39099 11261
rect 39133 11227 39145 11261
rect 39087 11193 39145 11227
rect 39087 11159 39099 11193
rect 39133 11159 39145 11193
rect 39087 11125 39145 11159
rect 39087 11091 39099 11125
rect 39133 11091 39145 11125
rect 39087 11057 39145 11091
rect 39087 11023 39099 11057
rect 39133 11023 39145 11057
rect 39087 10989 39145 11023
rect 39087 10955 39099 10989
rect 39133 10955 39145 10989
rect 39087 10914 39145 10955
rect 39345 11873 39403 11914
rect 39345 11839 39357 11873
rect 39391 11839 39403 11873
rect 39345 11805 39403 11839
rect 39345 11771 39357 11805
rect 39391 11771 39403 11805
rect 39345 11737 39403 11771
rect 39345 11703 39357 11737
rect 39391 11703 39403 11737
rect 39345 11669 39403 11703
rect 39345 11635 39357 11669
rect 39391 11635 39403 11669
rect 39345 11601 39403 11635
rect 39345 11567 39357 11601
rect 39391 11567 39403 11601
rect 39345 11533 39403 11567
rect 39345 11499 39357 11533
rect 39391 11499 39403 11533
rect 39345 11465 39403 11499
rect 39345 11431 39357 11465
rect 39391 11431 39403 11465
rect 39345 11397 39403 11431
rect 39345 11363 39357 11397
rect 39391 11363 39403 11397
rect 39345 11329 39403 11363
rect 39345 11295 39357 11329
rect 39391 11295 39403 11329
rect 39345 11261 39403 11295
rect 39345 11227 39357 11261
rect 39391 11227 39403 11261
rect 39345 11193 39403 11227
rect 39345 11159 39357 11193
rect 39391 11159 39403 11193
rect 39345 11125 39403 11159
rect 39345 11091 39357 11125
rect 39391 11091 39403 11125
rect 39345 11057 39403 11091
rect 39345 11023 39357 11057
rect 39391 11023 39403 11057
rect 39345 10989 39403 11023
rect 39345 10955 39357 10989
rect 39391 10955 39403 10989
rect 39345 10914 39403 10955
rect 39603 11873 39661 11914
rect 39603 11839 39615 11873
rect 39649 11839 39661 11873
rect 39603 11805 39661 11839
rect 39603 11771 39615 11805
rect 39649 11771 39661 11805
rect 39603 11737 39661 11771
rect 39603 11703 39615 11737
rect 39649 11703 39661 11737
rect 39603 11669 39661 11703
rect 39603 11635 39615 11669
rect 39649 11635 39661 11669
rect 39603 11601 39661 11635
rect 39603 11567 39615 11601
rect 39649 11567 39661 11601
rect 39603 11533 39661 11567
rect 39603 11499 39615 11533
rect 39649 11499 39661 11533
rect 39603 11465 39661 11499
rect 39603 11431 39615 11465
rect 39649 11431 39661 11465
rect 39603 11397 39661 11431
rect 39603 11363 39615 11397
rect 39649 11363 39661 11397
rect 39603 11329 39661 11363
rect 39603 11295 39615 11329
rect 39649 11295 39661 11329
rect 39603 11261 39661 11295
rect 39603 11227 39615 11261
rect 39649 11227 39661 11261
rect 39603 11193 39661 11227
rect 39603 11159 39615 11193
rect 39649 11159 39661 11193
rect 39603 11125 39661 11159
rect 39603 11091 39615 11125
rect 39649 11091 39661 11125
rect 39603 11057 39661 11091
rect 39603 11023 39615 11057
rect 39649 11023 39661 11057
rect 39603 10989 39661 11023
rect 39603 10955 39615 10989
rect 39649 10955 39661 10989
rect 39603 10914 39661 10955
rect 39861 11873 39919 11914
rect 39861 11839 39873 11873
rect 39907 11839 39919 11873
rect 39861 11805 39919 11839
rect 39861 11771 39873 11805
rect 39907 11771 39919 11805
rect 39861 11737 39919 11771
rect 39861 11703 39873 11737
rect 39907 11703 39919 11737
rect 39861 11669 39919 11703
rect 39861 11635 39873 11669
rect 39907 11635 39919 11669
rect 39861 11601 39919 11635
rect 39861 11567 39873 11601
rect 39907 11567 39919 11601
rect 39861 11533 39919 11567
rect 39861 11499 39873 11533
rect 39907 11499 39919 11533
rect 39861 11465 39919 11499
rect 39861 11431 39873 11465
rect 39907 11431 39919 11465
rect 39861 11397 39919 11431
rect 39861 11363 39873 11397
rect 39907 11363 39919 11397
rect 39861 11329 39919 11363
rect 39861 11295 39873 11329
rect 39907 11295 39919 11329
rect 39861 11261 39919 11295
rect 39861 11227 39873 11261
rect 39907 11227 39919 11261
rect 39861 11193 39919 11227
rect 39861 11159 39873 11193
rect 39907 11159 39919 11193
rect 39861 11125 39919 11159
rect 39861 11091 39873 11125
rect 39907 11091 39919 11125
rect 39861 11057 39919 11091
rect 39861 11023 39873 11057
rect 39907 11023 39919 11057
rect 39861 10989 39919 11023
rect 39861 10955 39873 10989
rect 39907 10955 39919 10989
rect 39861 10914 39919 10955
rect 40119 11873 40177 11914
rect 40119 11839 40131 11873
rect 40165 11839 40177 11873
rect 40119 11805 40177 11839
rect 40119 11771 40131 11805
rect 40165 11771 40177 11805
rect 40119 11737 40177 11771
rect 40119 11703 40131 11737
rect 40165 11703 40177 11737
rect 40119 11669 40177 11703
rect 40119 11635 40131 11669
rect 40165 11635 40177 11669
rect 40119 11601 40177 11635
rect 40119 11567 40131 11601
rect 40165 11567 40177 11601
rect 40119 11533 40177 11567
rect 40119 11499 40131 11533
rect 40165 11499 40177 11533
rect 40119 11465 40177 11499
rect 40119 11431 40131 11465
rect 40165 11431 40177 11465
rect 40119 11397 40177 11431
rect 40119 11363 40131 11397
rect 40165 11363 40177 11397
rect 40119 11329 40177 11363
rect 40119 11295 40131 11329
rect 40165 11295 40177 11329
rect 40119 11261 40177 11295
rect 40119 11227 40131 11261
rect 40165 11227 40177 11261
rect 40119 11193 40177 11227
rect 40119 11159 40131 11193
rect 40165 11159 40177 11193
rect 40119 11125 40177 11159
rect 40119 11091 40131 11125
rect 40165 11091 40177 11125
rect 40119 11057 40177 11091
rect 40119 11023 40131 11057
rect 40165 11023 40177 11057
rect 40119 10989 40177 11023
rect 40119 10955 40131 10989
rect 40165 10955 40177 10989
rect 40119 10914 40177 10955
rect 40377 11873 40435 11914
rect 40377 11839 40389 11873
rect 40423 11839 40435 11873
rect 40377 11805 40435 11839
rect 40377 11771 40389 11805
rect 40423 11771 40435 11805
rect 40377 11737 40435 11771
rect 40377 11703 40389 11737
rect 40423 11703 40435 11737
rect 40377 11669 40435 11703
rect 40377 11635 40389 11669
rect 40423 11635 40435 11669
rect 40377 11601 40435 11635
rect 40377 11567 40389 11601
rect 40423 11567 40435 11601
rect 40377 11533 40435 11567
rect 40377 11499 40389 11533
rect 40423 11499 40435 11533
rect 40377 11465 40435 11499
rect 40377 11431 40389 11465
rect 40423 11431 40435 11465
rect 40377 11397 40435 11431
rect 40377 11363 40389 11397
rect 40423 11363 40435 11397
rect 40377 11329 40435 11363
rect 40377 11295 40389 11329
rect 40423 11295 40435 11329
rect 40377 11261 40435 11295
rect 40377 11227 40389 11261
rect 40423 11227 40435 11261
rect 40377 11193 40435 11227
rect 40377 11159 40389 11193
rect 40423 11159 40435 11193
rect 40377 11125 40435 11159
rect 40377 11091 40389 11125
rect 40423 11091 40435 11125
rect 40377 11057 40435 11091
rect 40377 11023 40389 11057
rect 40423 11023 40435 11057
rect 40377 10989 40435 11023
rect 40377 10955 40389 10989
rect 40423 10955 40435 10989
rect 40377 10914 40435 10955
rect 40635 11873 40693 11914
rect 40635 11839 40647 11873
rect 40681 11839 40693 11873
rect 40635 11805 40693 11839
rect 40635 11771 40647 11805
rect 40681 11771 40693 11805
rect 40635 11737 40693 11771
rect 40635 11703 40647 11737
rect 40681 11703 40693 11737
rect 40635 11669 40693 11703
rect 40635 11635 40647 11669
rect 40681 11635 40693 11669
rect 40635 11601 40693 11635
rect 40635 11567 40647 11601
rect 40681 11567 40693 11601
rect 40635 11533 40693 11567
rect 40635 11499 40647 11533
rect 40681 11499 40693 11533
rect 40635 11465 40693 11499
rect 40635 11431 40647 11465
rect 40681 11431 40693 11465
rect 40635 11397 40693 11431
rect 40635 11363 40647 11397
rect 40681 11363 40693 11397
rect 40635 11329 40693 11363
rect 40635 11295 40647 11329
rect 40681 11295 40693 11329
rect 40635 11261 40693 11295
rect 40635 11227 40647 11261
rect 40681 11227 40693 11261
rect 40635 11193 40693 11227
rect 40635 11159 40647 11193
rect 40681 11159 40693 11193
rect 40635 11125 40693 11159
rect 40635 11091 40647 11125
rect 40681 11091 40693 11125
rect 40635 11057 40693 11091
rect 40635 11023 40647 11057
rect 40681 11023 40693 11057
rect 40635 10989 40693 11023
rect 40635 10955 40647 10989
rect 40681 10955 40693 10989
rect 40635 10914 40693 10955
rect 40893 11873 40951 11914
rect 40893 11839 40905 11873
rect 40939 11839 40951 11873
rect 40893 11805 40951 11839
rect 40893 11771 40905 11805
rect 40939 11771 40951 11805
rect 40893 11737 40951 11771
rect 40893 11703 40905 11737
rect 40939 11703 40951 11737
rect 40893 11669 40951 11703
rect 40893 11635 40905 11669
rect 40939 11635 40951 11669
rect 40893 11601 40951 11635
rect 40893 11567 40905 11601
rect 40939 11567 40951 11601
rect 40893 11533 40951 11567
rect 40893 11499 40905 11533
rect 40939 11499 40951 11533
rect 40893 11465 40951 11499
rect 40893 11431 40905 11465
rect 40939 11431 40951 11465
rect 40893 11397 40951 11431
rect 40893 11363 40905 11397
rect 40939 11363 40951 11397
rect 40893 11329 40951 11363
rect 40893 11295 40905 11329
rect 40939 11295 40951 11329
rect 40893 11261 40951 11295
rect 40893 11227 40905 11261
rect 40939 11227 40951 11261
rect 40893 11193 40951 11227
rect 40893 11159 40905 11193
rect 40939 11159 40951 11193
rect 40893 11125 40951 11159
rect 40893 11091 40905 11125
rect 40939 11091 40951 11125
rect 40893 11057 40951 11091
rect 40893 11023 40905 11057
rect 40939 11023 40951 11057
rect 40893 10989 40951 11023
rect 40893 10955 40905 10989
rect 40939 10955 40951 10989
rect 40893 10914 40951 10955
rect 41151 11873 41209 11914
rect 41151 11839 41163 11873
rect 41197 11839 41209 11873
rect 41151 11805 41209 11839
rect 41151 11771 41163 11805
rect 41197 11771 41209 11805
rect 41151 11737 41209 11771
rect 41151 11703 41163 11737
rect 41197 11703 41209 11737
rect 41151 11669 41209 11703
rect 41151 11635 41163 11669
rect 41197 11635 41209 11669
rect 41151 11601 41209 11635
rect 41151 11567 41163 11601
rect 41197 11567 41209 11601
rect 41151 11533 41209 11567
rect 41151 11499 41163 11533
rect 41197 11499 41209 11533
rect 41151 11465 41209 11499
rect 41151 11431 41163 11465
rect 41197 11431 41209 11465
rect 41151 11397 41209 11431
rect 41151 11363 41163 11397
rect 41197 11363 41209 11397
rect 41151 11329 41209 11363
rect 41151 11295 41163 11329
rect 41197 11295 41209 11329
rect 41151 11261 41209 11295
rect 41151 11227 41163 11261
rect 41197 11227 41209 11261
rect 41151 11193 41209 11227
rect 41151 11159 41163 11193
rect 41197 11159 41209 11193
rect 41151 11125 41209 11159
rect 41151 11091 41163 11125
rect 41197 11091 41209 11125
rect 41151 11057 41209 11091
rect 41151 11023 41163 11057
rect 41197 11023 41209 11057
rect 41151 10989 41209 11023
rect 41151 10955 41163 10989
rect 41197 10955 41209 10989
rect 41151 10914 41209 10955
rect 41409 11873 41467 11914
rect 41409 11839 41421 11873
rect 41455 11839 41467 11873
rect 41409 11805 41467 11839
rect 41409 11771 41421 11805
rect 41455 11771 41467 11805
rect 41409 11737 41467 11771
rect 41409 11703 41421 11737
rect 41455 11703 41467 11737
rect 41409 11669 41467 11703
rect 41409 11635 41421 11669
rect 41455 11635 41467 11669
rect 41409 11601 41467 11635
rect 41409 11567 41421 11601
rect 41455 11567 41467 11601
rect 41409 11533 41467 11567
rect 41409 11499 41421 11533
rect 41455 11499 41467 11533
rect 41409 11465 41467 11499
rect 41409 11431 41421 11465
rect 41455 11431 41467 11465
rect 41409 11397 41467 11431
rect 41409 11363 41421 11397
rect 41455 11363 41467 11397
rect 41409 11329 41467 11363
rect 41409 11295 41421 11329
rect 41455 11295 41467 11329
rect 41409 11261 41467 11295
rect 41409 11227 41421 11261
rect 41455 11227 41467 11261
rect 41409 11193 41467 11227
rect 41409 11159 41421 11193
rect 41455 11159 41467 11193
rect 41409 11125 41467 11159
rect 41409 11091 41421 11125
rect 41455 11091 41467 11125
rect 41409 11057 41467 11091
rect 41409 11023 41421 11057
rect 41455 11023 41467 11057
rect 41409 10989 41467 11023
rect 41409 10955 41421 10989
rect 41455 10955 41467 10989
rect 41409 10914 41467 10955
rect 41667 11873 41725 11914
rect 41667 11839 41679 11873
rect 41713 11839 41725 11873
rect 41667 11805 41725 11839
rect 41667 11771 41679 11805
rect 41713 11771 41725 11805
rect 41667 11737 41725 11771
rect 41667 11703 41679 11737
rect 41713 11703 41725 11737
rect 41667 11669 41725 11703
rect 41667 11635 41679 11669
rect 41713 11635 41725 11669
rect 41667 11601 41725 11635
rect 41667 11567 41679 11601
rect 41713 11567 41725 11601
rect 41667 11533 41725 11567
rect 41667 11499 41679 11533
rect 41713 11499 41725 11533
rect 41667 11465 41725 11499
rect 41667 11431 41679 11465
rect 41713 11431 41725 11465
rect 41667 11397 41725 11431
rect 41667 11363 41679 11397
rect 41713 11363 41725 11397
rect 41667 11329 41725 11363
rect 41667 11295 41679 11329
rect 41713 11295 41725 11329
rect 41667 11261 41725 11295
rect 41667 11227 41679 11261
rect 41713 11227 41725 11261
rect 41667 11193 41725 11227
rect 41667 11159 41679 11193
rect 41713 11159 41725 11193
rect 41667 11125 41725 11159
rect 41667 11091 41679 11125
rect 41713 11091 41725 11125
rect 41667 11057 41725 11091
rect 41667 11023 41679 11057
rect 41713 11023 41725 11057
rect 41667 10989 41725 11023
rect 41667 10955 41679 10989
rect 41713 10955 41725 10989
rect 41667 10914 41725 10955
rect 41925 11873 41983 11914
rect 41925 11839 41937 11873
rect 41971 11839 41983 11873
rect 41925 11805 41983 11839
rect 41925 11771 41937 11805
rect 41971 11771 41983 11805
rect 41925 11737 41983 11771
rect 41925 11703 41937 11737
rect 41971 11703 41983 11737
rect 41925 11669 41983 11703
rect 41925 11635 41937 11669
rect 41971 11635 41983 11669
rect 41925 11601 41983 11635
rect 41925 11567 41937 11601
rect 41971 11567 41983 11601
rect 41925 11533 41983 11567
rect 41925 11499 41937 11533
rect 41971 11499 41983 11533
rect 41925 11465 41983 11499
rect 41925 11431 41937 11465
rect 41971 11431 41983 11465
rect 41925 11397 41983 11431
rect 41925 11363 41937 11397
rect 41971 11363 41983 11397
rect 41925 11329 41983 11363
rect 41925 11295 41937 11329
rect 41971 11295 41983 11329
rect 41925 11261 41983 11295
rect 41925 11227 41937 11261
rect 41971 11227 41983 11261
rect 41925 11193 41983 11227
rect 41925 11159 41937 11193
rect 41971 11159 41983 11193
rect 41925 11125 41983 11159
rect 41925 11091 41937 11125
rect 41971 11091 41983 11125
rect 41925 11057 41983 11091
rect 41925 11023 41937 11057
rect 41971 11023 41983 11057
rect 41925 10989 41983 11023
rect 41925 10955 41937 10989
rect 41971 10955 41983 10989
rect 41925 10914 41983 10955
rect 37800 10508 37858 10549
rect 37800 10474 37812 10508
rect 37846 10474 37858 10508
rect 37800 10440 37858 10474
rect 37800 10406 37812 10440
rect 37846 10406 37858 10440
rect 37800 10372 37858 10406
rect 37800 10338 37812 10372
rect 37846 10338 37858 10372
rect 37800 10304 37858 10338
rect 37800 10270 37812 10304
rect 37846 10270 37858 10304
rect 37800 10236 37858 10270
rect 37800 10202 37812 10236
rect 37846 10202 37858 10236
rect 37800 10168 37858 10202
rect 37800 10134 37812 10168
rect 37846 10134 37858 10168
rect 37800 10100 37858 10134
rect 37800 10066 37812 10100
rect 37846 10066 37858 10100
rect 37800 10032 37858 10066
rect 37800 9998 37812 10032
rect 37846 9998 37858 10032
rect 37800 9964 37858 9998
rect 37800 9930 37812 9964
rect 37846 9930 37858 9964
rect 37800 9896 37858 9930
rect 37800 9862 37812 9896
rect 37846 9862 37858 9896
rect 37800 9828 37858 9862
rect 37800 9794 37812 9828
rect 37846 9794 37858 9828
rect 37800 9760 37858 9794
rect 37800 9726 37812 9760
rect 37846 9726 37858 9760
rect 37800 9692 37858 9726
rect 37800 9658 37812 9692
rect 37846 9658 37858 9692
rect 37800 9624 37858 9658
rect 37800 9590 37812 9624
rect 37846 9590 37858 9624
rect 37800 9549 37858 9590
rect 38058 10508 38116 10549
rect 38058 10474 38070 10508
rect 38104 10474 38116 10508
rect 38058 10440 38116 10474
rect 38058 10406 38070 10440
rect 38104 10406 38116 10440
rect 38058 10372 38116 10406
rect 38058 10338 38070 10372
rect 38104 10338 38116 10372
rect 38058 10304 38116 10338
rect 38058 10270 38070 10304
rect 38104 10270 38116 10304
rect 38058 10236 38116 10270
rect 38058 10202 38070 10236
rect 38104 10202 38116 10236
rect 38058 10168 38116 10202
rect 38058 10134 38070 10168
rect 38104 10134 38116 10168
rect 38058 10100 38116 10134
rect 38058 10066 38070 10100
rect 38104 10066 38116 10100
rect 38058 10032 38116 10066
rect 38058 9998 38070 10032
rect 38104 9998 38116 10032
rect 38058 9964 38116 9998
rect 38058 9930 38070 9964
rect 38104 9930 38116 9964
rect 38058 9896 38116 9930
rect 38058 9862 38070 9896
rect 38104 9862 38116 9896
rect 38058 9828 38116 9862
rect 38058 9794 38070 9828
rect 38104 9794 38116 9828
rect 38058 9760 38116 9794
rect 38058 9726 38070 9760
rect 38104 9726 38116 9760
rect 38058 9692 38116 9726
rect 38058 9658 38070 9692
rect 38104 9658 38116 9692
rect 38058 9624 38116 9658
rect 38058 9590 38070 9624
rect 38104 9590 38116 9624
rect 38058 9549 38116 9590
rect 38266 10508 38324 10549
rect 38266 10474 38278 10508
rect 38312 10474 38324 10508
rect 38266 10440 38324 10474
rect 38266 10406 38278 10440
rect 38312 10406 38324 10440
rect 38266 10372 38324 10406
rect 38266 10338 38278 10372
rect 38312 10338 38324 10372
rect 38266 10304 38324 10338
rect 38266 10270 38278 10304
rect 38312 10270 38324 10304
rect 38266 10236 38324 10270
rect 38266 10202 38278 10236
rect 38312 10202 38324 10236
rect 38266 10168 38324 10202
rect 38266 10134 38278 10168
rect 38312 10134 38324 10168
rect 38266 10100 38324 10134
rect 38266 10066 38278 10100
rect 38312 10066 38324 10100
rect 38266 10032 38324 10066
rect 38266 9998 38278 10032
rect 38312 9998 38324 10032
rect 38266 9964 38324 9998
rect 38266 9930 38278 9964
rect 38312 9930 38324 9964
rect 38266 9896 38324 9930
rect 38266 9862 38278 9896
rect 38312 9862 38324 9896
rect 38266 9828 38324 9862
rect 38266 9794 38278 9828
rect 38312 9794 38324 9828
rect 38266 9760 38324 9794
rect 38266 9726 38278 9760
rect 38312 9726 38324 9760
rect 38266 9692 38324 9726
rect 38266 9658 38278 9692
rect 38312 9658 38324 9692
rect 38266 9624 38324 9658
rect 38266 9590 38278 9624
rect 38312 9590 38324 9624
rect 38266 9549 38324 9590
rect 38524 10508 38582 10549
rect 38524 10474 38536 10508
rect 38570 10474 38582 10508
rect 38524 10440 38582 10474
rect 38524 10406 38536 10440
rect 38570 10406 38582 10440
rect 38524 10372 38582 10406
rect 38524 10338 38536 10372
rect 38570 10338 38582 10372
rect 38524 10304 38582 10338
rect 38524 10270 38536 10304
rect 38570 10270 38582 10304
rect 38524 10236 38582 10270
rect 38524 10202 38536 10236
rect 38570 10202 38582 10236
rect 38524 10168 38582 10202
rect 38524 10134 38536 10168
rect 38570 10134 38582 10168
rect 38524 10100 38582 10134
rect 38524 10066 38536 10100
rect 38570 10066 38582 10100
rect 38524 10032 38582 10066
rect 38524 9998 38536 10032
rect 38570 9998 38582 10032
rect 38524 9964 38582 9998
rect 38524 9930 38536 9964
rect 38570 9930 38582 9964
rect 38524 9896 38582 9930
rect 38524 9862 38536 9896
rect 38570 9862 38582 9896
rect 38524 9828 38582 9862
rect 38524 9794 38536 9828
rect 38570 9794 38582 9828
rect 38524 9760 38582 9794
rect 38524 9726 38536 9760
rect 38570 9726 38582 9760
rect 38524 9692 38582 9726
rect 38524 9658 38536 9692
rect 38570 9658 38582 9692
rect 38524 9624 38582 9658
rect 38524 9590 38536 9624
rect 38570 9590 38582 9624
rect 38524 9549 38582 9590
rect 38782 10508 38840 10549
rect 38782 10474 38794 10508
rect 38828 10474 38840 10508
rect 38782 10440 38840 10474
rect 38782 10406 38794 10440
rect 38828 10406 38840 10440
rect 38782 10372 38840 10406
rect 38782 10338 38794 10372
rect 38828 10338 38840 10372
rect 38782 10304 38840 10338
rect 38782 10270 38794 10304
rect 38828 10270 38840 10304
rect 38782 10236 38840 10270
rect 38782 10202 38794 10236
rect 38828 10202 38840 10236
rect 38782 10168 38840 10202
rect 38782 10134 38794 10168
rect 38828 10134 38840 10168
rect 38782 10100 38840 10134
rect 38782 10066 38794 10100
rect 38828 10066 38840 10100
rect 38782 10032 38840 10066
rect 38782 9998 38794 10032
rect 38828 9998 38840 10032
rect 38782 9964 38840 9998
rect 38782 9930 38794 9964
rect 38828 9930 38840 9964
rect 38782 9896 38840 9930
rect 38782 9862 38794 9896
rect 38828 9862 38840 9896
rect 38782 9828 38840 9862
rect 38782 9794 38794 9828
rect 38828 9794 38840 9828
rect 38782 9760 38840 9794
rect 38782 9726 38794 9760
rect 38828 9726 38840 9760
rect 38782 9692 38840 9726
rect 38782 9658 38794 9692
rect 38828 9658 38840 9692
rect 38782 9624 38840 9658
rect 38782 9590 38794 9624
rect 38828 9590 38840 9624
rect 38782 9549 38840 9590
rect 39040 10508 39098 10549
rect 39040 10474 39052 10508
rect 39086 10474 39098 10508
rect 39040 10440 39098 10474
rect 39040 10406 39052 10440
rect 39086 10406 39098 10440
rect 39040 10372 39098 10406
rect 39040 10338 39052 10372
rect 39086 10338 39098 10372
rect 39040 10304 39098 10338
rect 39040 10270 39052 10304
rect 39086 10270 39098 10304
rect 39040 10236 39098 10270
rect 39040 10202 39052 10236
rect 39086 10202 39098 10236
rect 39040 10168 39098 10202
rect 39040 10134 39052 10168
rect 39086 10134 39098 10168
rect 39040 10100 39098 10134
rect 39040 10066 39052 10100
rect 39086 10066 39098 10100
rect 39040 10032 39098 10066
rect 39040 9998 39052 10032
rect 39086 9998 39098 10032
rect 39040 9964 39098 9998
rect 39040 9930 39052 9964
rect 39086 9930 39098 9964
rect 39040 9896 39098 9930
rect 39040 9862 39052 9896
rect 39086 9862 39098 9896
rect 39040 9828 39098 9862
rect 39040 9794 39052 9828
rect 39086 9794 39098 9828
rect 39040 9760 39098 9794
rect 39040 9726 39052 9760
rect 39086 9726 39098 9760
rect 39040 9692 39098 9726
rect 39040 9658 39052 9692
rect 39086 9658 39098 9692
rect 39040 9624 39098 9658
rect 39040 9590 39052 9624
rect 39086 9590 39098 9624
rect 39040 9549 39098 9590
rect 39298 10508 39356 10549
rect 39298 10474 39310 10508
rect 39344 10474 39356 10508
rect 39298 10440 39356 10474
rect 39298 10406 39310 10440
rect 39344 10406 39356 10440
rect 39298 10372 39356 10406
rect 39298 10338 39310 10372
rect 39344 10338 39356 10372
rect 39298 10304 39356 10338
rect 39298 10270 39310 10304
rect 39344 10270 39356 10304
rect 39298 10236 39356 10270
rect 39298 10202 39310 10236
rect 39344 10202 39356 10236
rect 39298 10168 39356 10202
rect 39298 10134 39310 10168
rect 39344 10134 39356 10168
rect 39298 10100 39356 10134
rect 39298 10066 39310 10100
rect 39344 10066 39356 10100
rect 39298 10032 39356 10066
rect 39298 9998 39310 10032
rect 39344 9998 39356 10032
rect 39298 9964 39356 9998
rect 39298 9930 39310 9964
rect 39344 9930 39356 9964
rect 39298 9896 39356 9930
rect 39298 9862 39310 9896
rect 39344 9862 39356 9896
rect 39298 9828 39356 9862
rect 39298 9794 39310 9828
rect 39344 9794 39356 9828
rect 39298 9760 39356 9794
rect 39298 9726 39310 9760
rect 39344 9726 39356 9760
rect 39298 9692 39356 9726
rect 39298 9658 39310 9692
rect 39344 9658 39356 9692
rect 39298 9624 39356 9658
rect 39298 9590 39310 9624
rect 39344 9590 39356 9624
rect 39298 9549 39356 9590
rect 39556 10508 39614 10549
rect 39556 10474 39568 10508
rect 39602 10474 39614 10508
rect 39556 10440 39614 10474
rect 39556 10406 39568 10440
rect 39602 10406 39614 10440
rect 39556 10372 39614 10406
rect 39556 10338 39568 10372
rect 39602 10338 39614 10372
rect 39556 10304 39614 10338
rect 39556 10270 39568 10304
rect 39602 10270 39614 10304
rect 39556 10236 39614 10270
rect 39556 10202 39568 10236
rect 39602 10202 39614 10236
rect 39556 10168 39614 10202
rect 39556 10134 39568 10168
rect 39602 10134 39614 10168
rect 39556 10100 39614 10134
rect 39556 10066 39568 10100
rect 39602 10066 39614 10100
rect 39556 10032 39614 10066
rect 39556 9998 39568 10032
rect 39602 9998 39614 10032
rect 39556 9964 39614 9998
rect 39556 9930 39568 9964
rect 39602 9930 39614 9964
rect 39556 9896 39614 9930
rect 39556 9862 39568 9896
rect 39602 9862 39614 9896
rect 39556 9828 39614 9862
rect 39556 9794 39568 9828
rect 39602 9794 39614 9828
rect 39556 9760 39614 9794
rect 39556 9726 39568 9760
rect 39602 9726 39614 9760
rect 39556 9692 39614 9726
rect 39556 9658 39568 9692
rect 39602 9658 39614 9692
rect 39556 9624 39614 9658
rect 39556 9590 39568 9624
rect 39602 9590 39614 9624
rect 39556 9549 39614 9590
rect 39814 10508 39872 10549
rect 39814 10474 39826 10508
rect 39860 10474 39872 10508
rect 39814 10440 39872 10474
rect 39814 10406 39826 10440
rect 39860 10406 39872 10440
rect 39814 10372 39872 10406
rect 39814 10338 39826 10372
rect 39860 10338 39872 10372
rect 39814 10304 39872 10338
rect 39814 10270 39826 10304
rect 39860 10270 39872 10304
rect 39814 10236 39872 10270
rect 39814 10202 39826 10236
rect 39860 10202 39872 10236
rect 39814 10168 39872 10202
rect 39814 10134 39826 10168
rect 39860 10134 39872 10168
rect 39814 10100 39872 10134
rect 39814 10066 39826 10100
rect 39860 10066 39872 10100
rect 39814 10032 39872 10066
rect 39814 9998 39826 10032
rect 39860 9998 39872 10032
rect 39814 9964 39872 9998
rect 39814 9930 39826 9964
rect 39860 9930 39872 9964
rect 39814 9896 39872 9930
rect 39814 9862 39826 9896
rect 39860 9862 39872 9896
rect 39814 9828 39872 9862
rect 39814 9794 39826 9828
rect 39860 9794 39872 9828
rect 39814 9760 39872 9794
rect 39814 9726 39826 9760
rect 39860 9726 39872 9760
rect 39814 9692 39872 9726
rect 39814 9658 39826 9692
rect 39860 9658 39872 9692
rect 39814 9624 39872 9658
rect 39814 9590 39826 9624
rect 39860 9590 39872 9624
rect 39814 9549 39872 9590
rect 40072 10508 40130 10549
rect 40072 10474 40084 10508
rect 40118 10474 40130 10508
rect 40072 10440 40130 10474
rect 40072 10406 40084 10440
rect 40118 10406 40130 10440
rect 40072 10372 40130 10406
rect 40072 10338 40084 10372
rect 40118 10338 40130 10372
rect 40072 10304 40130 10338
rect 40072 10270 40084 10304
rect 40118 10270 40130 10304
rect 40072 10236 40130 10270
rect 40072 10202 40084 10236
rect 40118 10202 40130 10236
rect 40072 10168 40130 10202
rect 40072 10134 40084 10168
rect 40118 10134 40130 10168
rect 40072 10100 40130 10134
rect 40072 10066 40084 10100
rect 40118 10066 40130 10100
rect 40072 10032 40130 10066
rect 40072 9998 40084 10032
rect 40118 9998 40130 10032
rect 40072 9964 40130 9998
rect 40072 9930 40084 9964
rect 40118 9930 40130 9964
rect 40072 9896 40130 9930
rect 40072 9862 40084 9896
rect 40118 9862 40130 9896
rect 40072 9828 40130 9862
rect 40072 9794 40084 9828
rect 40118 9794 40130 9828
rect 40072 9760 40130 9794
rect 40072 9726 40084 9760
rect 40118 9726 40130 9760
rect 40072 9692 40130 9726
rect 40072 9658 40084 9692
rect 40118 9658 40130 9692
rect 40072 9624 40130 9658
rect 40072 9590 40084 9624
rect 40118 9590 40130 9624
rect 40072 9549 40130 9590
rect 40330 10508 40388 10549
rect 40330 10474 40342 10508
rect 40376 10474 40388 10508
rect 40330 10440 40388 10474
rect 40330 10406 40342 10440
rect 40376 10406 40388 10440
rect 40330 10372 40388 10406
rect 40330 10338 40342 10372
rect 40376 10338 40388 10372
rect 40330 10304 40388 10338
rect 40330 10270 40342 10304
rect 40376 10270 40388 10304
rect 40330 10236 40388 10270
rect 40330 10202 40342 10236
rect 40376 10202 40388 10236
rect 40330 10168 40388 10202
rect 40330 10134 40342 10168
rect 40376 10134 40388 10168
rect 40330 10100 40388 10134
rect 40330 10066 40342 10100
rect 40376 10066 40388 10100
rect 40330 10032 40388 10066
rect 40330 9998 40342 10032
rect 40376 9998 40388 10032
rect 40330 9964 40388 9998
rect 40330 9930 40342 9964
rect 40376 9930 40388 9964
rect 40330 9896 40388 9930
rect 40330 9862 40342 9896
rect 40376 9862 40388 9896
rect 40330 9828 40388 9862
rect 40330 9794 40342 9828
rect 40376 9794 40388 9828
rect 40330 9760 40388 9794
rect 40330 9726 40342 9760
rect 40376 9726 40388 9760
rect 40330 9692 40388 9726
rect 40330 9658 40342 9692
rect 40376 9658 40388 9692
rect 40330 9624 40388 9658
rect 40330 9590 40342 9624
rect 40376 9590 40388 9624
rect 40330 9549 40388 9590
rect 40588 10508 40646 10549
rect 40588 10474 40600 10508
rect 40634 10474 40646 10508
rect 40588 10440 40646 10474
rect 40588 10406 40600 10440
rect 40634 10406 40646 10440
rect 40588 10372 40646 10406
rect 40588 10338 40600 10372
rect 40634 10338 40646 10372
rect 40588 10304 40646 10338
rect 40588 10270 40600 10304
rect 40634 10270 40646 10304
rect 40588 10236 40646 10270
rect 40588 10202 40600 10236
rect 40634 10202 40646 10236
rect 40588 10168 40646 10202
rect 40588 10134 40600 10168
rect 40634 10134 40646 10168
rect 40588 10100 40646 10134
rect 40588 10066 40600 10100
rect 40634 10066 40646 10100
rect 40588 10032 40646 10066
rect 40588 9998 40600 10032
rect 40634 9998 40646 10032
rect 40588 9964 40646 9998
rect 40588 9930 40600 9964
rect 40634 9930 40646 9964
rect 40588 9896 40646 9930
rect 40588 9862 40600 9896
rect 40634 9862 40646 9896
rect 40588 9828 40646 9862
rect 40588 9794 40600 9828
rect 40634 9794 40646 9828
rect 40588 9760 40646 9794
rect 40588 9726 40600 9760
rect 40634 9726 40646 9760
rect 40588 9692 40646 9726
rect 40588 9658 40600 9692
rect 40634 9658 40646 9692
rect 40588 9624 40646 9658
rect 40588 9590 40600 9624
rect 40634 9590 40646 9624
rect 40588 9549 40646 9590
rect 40846 10508 40904 10549
rect 40846 10474 40858 10508
rect 40892 10474 40904 10508
rect 40846 10440 40904 10474
rect 40846 10406 40858 10440
rect 40892 10406 40904 10440
rect 40846 10372 40904 10406
rect 40846 10338 40858 10372
rect 40892 10338 40904 10372
rect 40846 10304 40904 10338
rect 40846 10270 40858 10304
rect 40892 10270 40904 10304
rect 40846 10236 40904 10270
rect 40846 10202 40858 10236
rect 40892 10202 40904 10236
rect 40846 10168 40904 10202
rect 40846 10134 40858 10168
rect 40892 10134 40904 10168
rect 40846 10100 40904 10134
rect 40846 10066 40858 10100
rect 40892 10066 40904 10100
rect 40846 10032 40904 10066
rect 40846 9998 40858 10032
rect 40892 9998 40904 10032
rect 40846 9964 40904 9998
rect 40846 9930 40858 9964
rect 40892 9930 40904 9964
rect 40846 9896 40904 9930
rect 40846 9862 40858 9896
rect 40892 9862 40904 9896
rect 40846 9828 40904 9862
rect 40846 9794 40858 9828
rect 40892 9794 40904 9828
rect 40846 9760 40904 9794
rect 40846 9726 40858 9760
rect 40892 9726 40904 9760
rect 40846 9692 40904 9726
rect 40846 9658 40858 9692
rect 40892 9658 40904 9692
rect 40846 9624 40904 9658
rect 40846 9590 40858 9624
rect 40892 9590 40904 9624
rect 40846 9549 40904 9590
rect 37800 8257 37858 8288
rect 37800 8223 37812 8257
rect 37846 8223 37858 8257
rect 37800 8189 37858 8223
rect 37800 8155 37812 8189
rect 37846 8155 37858 8189
rect 37800 8121 37858 8155
rect 37800 8087 37812 8121
rect 37846 8087 37858 8121
rect 37800 8053 37858 8087
rect 37800 8019 37812 8053
rect 37846 8019 37858 8053
rect 37800 7985 37858 8019
rect 37800 7951 37812 7985
rect 37846 7951 37858 7985
rect 37800 7917 37858 7951
rect 37800 7883 37812 7917
rect 37846 7883 37858 7917
rect 37800 7849 37858 7883
rect 37800 7815 37812 7849
rect 37846 7815 37858 7849
rect 37800 7781 37858 7815
rect 37800 7747 37812 7781
rect 37846 7747 37858 7781
rect 37800 7713 37858 7747
rect 37800 7679 37812 7713
rect 37846 7679 37858 7713
rect 37800 7645 37858 7679
rect 37800 7611 37812 7645
rect 37846 7611 37858 7645
rect 37800 7577 37858 7611
rect 37800 7543 37812 7577
rect 37846 7543 37858 7577
rect 37800 7509 37858 7543
rect 37800 7475 37812 7509
rect 37846 7475 37858 7509
rect 37800 7441 37858 7475
rect 37800 7407 37812 7441
rect 37846 7407 37858 7441
rect 37800 7373 37858 7407
rect 37800 7339 37812 7373
rect 37846 7339 37858 7373
rect 37800 7305 37858 7339
rect 37800 7271 37812 7305
rect 37846 7271 37858 7305
rect 37800 7237 37858 7271
rect 37800 7203 37812 7237
rect 37846 7203 37858 7237
rect 37800 7169 37858 7203
rect 37800 7135 37812 7169
rect 37846 7135 37858 7169
rect 37800 7101 37858 7135
rect 37800 7067 37812 7101
rect 37846 7067 37858 7101
rect 37800 7033 37858 7067
rect 37800 6999 37812 7033
rect 37846 6999 37858 7033
rect 37800 6965 37858 6999
rect 37800 6931 37812 6965
rect 37846 6931 37858 6965
rect 37800 6897 37858 6931
rect 37800 6863 37812 6897
rect 37846 6863 37858 6897
rect 37800 6829 37858 6863
rect 37800 6795 37812 6829
rect 37846 6795 37858 6829
rect 37800 6761 37858 6795
rect 37800 6727 37812 6761
rect 37846 6727 37858 6761
rect 37800 6693 37858 6727
rect 37800 6659 37812 6693
rect 37846 6659 37858 6693
rect 37800 6625 37858 6659
rect 37800 6591 37812 6625
rect 37846 6591 37858 6625
rect 37800 6557 37858 6591
rect 37800 6523 37812 6557
rect 37846 6523 37858 6557
rect 37800 6489 37858 6523
rect 37800 6455 37812 6489
rect 37846 6455 37858 6489
rect 37800 6421 37858 6455
rect 37800 6387 37812 6421
rect 37846 6387 37858 6421
rect 37800 6353 37858 6387
rect 37800 6319 37812 6353
rect 37846 6319 37858 6353
rect 37800 6288 37858 6319
rect 38058 8257 38116 8288
rect 38058 8223 38070 8257
rect 38104 8223 38116 8257
rect 38058 8189 38116 8223
rect 38058 8155 38070 8189
rect 38104 8155 38116 8189
rect 38058 8121 38116 8155
rect 38058 8087 38070 8121
rect 38104 8087 38116 8121
rect 38058 8053 38116 8087
rect 38058 8019 38070 8053
rect 38104 8019 38116 8053
rect 38058 7985 38116 8019
rect 38058 7951 38070 7985
rect 38104 7951 38116 7985
rect 38058 7917 38116 7951
rect 38058 7883 38070 7917
rect 38104 7883 38116 7917
rect 38058 7849 38116 7883
rect 38058 7815 38070 7849
rect 38104 7815 38116 7849
rect 38058 7781 38116 7815
rect 38058 7747 38070 7781
rect 38104 7747 38116 7781
rect 38058 7713 38116 7747
rect 38058 7679 38070 7713
rect 38104 7679 38116 7713
rect 38058 7645 38116 7679
rect 38058 7611 38070 7645
rect 38104 7611 38116 7645
rect 38058 7577 38116 7611
rect 38058 7543 38070 7577
rect 38104 7543 38116 7577
rect 38058 7509 38116 7543
rect 38058 7475 38070 7509
rect 38104 7475 38116 7509
rect 38058 7441 38116 7475
rect 38058 7407 38070 7441
rect 38104 7407 38116 7441
rect 38058 7373 38116 7407
rect 38058 7339 38070 7373
rect 38104 7339 38116 7373
rect 38058 7305 38116 7339
rect 38058 7271 38070 7305
rect 38104 7271 38116 7305
rect 38058 7237 38116 7271
rect 38058 7203 38070 7237
rect 38104 7203 38116 7237
rect 38058 7169 38116 7203
rect 38058 7135 38070 7169
rect 38104 7135 38116 7169
rect 38058 7101 38116 7135
rect 38058 7067 38070 7101
rect 38104 7067 38116 7101
rect 38058 7033 38116 7067
rect 38058 6999 38070 7033
rect 38104 6999 38116 7033
rect 38058 6965 38116 6999
rect 38058 6931 38070 6965
rect 38104 6931 38116 6965
rect 38058 6897 38116 6931
rect 38058 6863 38070 6897
rect 38104 6863 38116 6897
rect 38058 6829 38116 6863
rect 38058 6795 38070 6829
rect 38104 6795 38116 6829
rect 38058 6761 38116 6795
rect 38058 6727 38070 6761
rect 38104 6727 38116 6761
rect 38058 6693 38116 6727
rect 38058 6659 38070 6693
rect 38104 6659 38116 6693
rect 38058 6625 38116 6659
rect 38058 6591 38070 6625
rect 38104 6591 38116 6625
rect 38058 6557 38116 6591
rect 38058 6523 38070 6557
rect 38104 6523 38116 6557
rect 38058 6489 38116 6523
rect 38058 6455 38070 6489
rect 38104 6455 38116 6489
rect 38058 6421 38116 6455
rect 38058 6387 38070 6421
rect 38104 6387 38116 6421
rect 38058 6353 38116 6387
rect 38058 6319 38070 6353
rect 38104 6319 38116 6353
rect 38058 6288 38116 6319
rect 38316 8257 38374 8288
rect 38316 8223 38328 8257
rect 38362 8223 38374 8257
rect 38316 8189 38374 8223
rect 38316 8155 38328 8189
rect 38362 8155 38374 8189
rect 38316 8121 38374 8155
rect 38316 8087 38328 8121
rect 38362 8087 38374 8121
rect 38316 8053 38374 8087
rect 38316 8019 38328 8053
rect 38362 8019 38374 8053
rect 38316 7985 38374 8019
rect 38316 7951 38328 7985
rect 38362 7951 38374 7985
rect 38316 7917 38374 7951
rect 38316 7883 38328 7917
rect 38362 7883 38374 7917
rect 38316 7849 38374 7883
rect 38316 7815 38328 7849
rect 38362 7815 38374 7849
rect 38316 7781 38374 7815
rect 38316 7747 38328 7781
rect 38362 7747 38374 7781
rect 38316 7713 38374 7747
rect 38316 7679 38328 7713
rect 38362 7679 38374 7713
rect 38316 7645 38374 7679
rect 38316 7611 38328 7645
rect 38362 7611 38374 7645
rect 38316 7577 38374 7611
rect 38316 7543 38328 7577
rect 38362 7543 38374 7577
rect 38316 7509 38374 7543
rect 38316 7475 38328 7509
rect 38362 7475 38374 7509
rect 38316 7441 38374 7475
rect 38316 7407 38328 7441
rect 38362 7407 38374 7441
rect 38316 7373 38374 7407
rect 38316 7339 38328 7373
rect 38362 7339 38374 7373
rect 38316 7305 38374 7339
rect 38316 7271 38328 7305
rect 38362 7271 38374 7305
rect 38316 7237 38374 7271
rect 38316 7203 38328 7237
rect 38362 7203 38374 7237
rect 38316 7169 38374 7203
rect 38316 7135 38328 7169
rect 38362 7135 38374 7169
rect 38316 7101 38374 7135
rect 38316 7067 38328 7101
rect 38362 7067 38374 7101
rect 38316 7033 38374 7067
rect 38316 6999 38328 7033
rect 38362 6999 38374 7033
rect 38316 6965 38374 6999
rect 38316 6931 38328 6965
rect 38362 6931 38374 6965
rect 38316 6897 38374 6931
rect 38316 6863 38328 6897
rect 38362 6863 38374 6897
rect 38316 6829 38374 6863
rect 38316 6795 38328 6829
rect 38362 6795 38374 6829
rect 38316 6761 38374 6795
rect 38316 6727 38328 6761
rect 38362 6727 38374 6761
rect 38316 6693 38374 6727
rect 38316 6659 38328 6693
rect 38362 6659 38374 6693
rect 38316 6625 38374 6659
rect 38316 6591 38328 6625
rect 38362 6591 38374 6625
rect 38316 6557 38374 6591
rect 38316 6523 38328 6557
rect 38362 6523 38374 6557
rect 38316 6489 38374 6523
rect 38316 6455 38328 6489
rect 38362 6455 38374 6489
rect 38316 6421 38374 6455
rect 38316 6387 38328 6421
rect 38362 6387 38374 6421
rect 38316 6353 38374 6387
rect 38316 6319 38328 6353
rect 38362 6319 38374 6353
rect 38316 6288 38374 6319
rect 38574 8257 38632 8288
rect 38574 8223 38586 8257
rect 38620 8223 38632 8257
rect 38574 8189 38632 8223
rect 38574 8155 38586 8189
rect 38620 8155 38632 8189
rect 38574 8121 38632 8155
rect 38574 8087 38586 8121
rect 38620 8087 38632 8121
rect 38574 8053 38632 8087
rect 38574 8019 38586 8053
rect 38620 8019 38632 8053
rect 38574 7985 38632 8019
rect 38574 7951 38586 7985
rect 38620 7951 38632 7985
rect 38574 7917 38632 7951
rect 38574 7883 38586 7917
rect 38620 7883 38632 7917
rect 38574 7849 38632 7883
rect 38574 7815 38586 7849
rect 38620 7815 38632 7849
rect 38574 7781 38632 7815
rect 38574 7747 38586 7781
rect 38620 7747 38632 7781
rect 38574 7713 38632 7747
rect 38574 7679 38586 7713
rect 38620 7679 38632 7713
rect 38574 7645 38632 7679
rect 38574 7611 38586 7645
rect 38620 7611 38632 7645
rect 38574 7577 38632 7611
rect 38574 7543 38586 7577
rect 38620 7543 38632 7577
rect 38574 7509 38632 7543
rect 38574 7475 38586 7509
rect 38620 7475 38632 7509
rect 38574 7441 38632 7475
rect 38574 7407 38586 7441
rect 38620 7407 38632 7441
rect 38574 7373 38632 7407
rect 38574 7339 38586 7373
rect 38620 7339 38632 7373
rect 38574 7305 38632 7339
rect 38574 7271 38586 7305
rect 38620 7271 38632 7305
rect 38574 7237 38632 7271
rect 38574 7203 38586 7237
rect 38620 7203 38632 7237
rect 38574 7169 38632 7203
rect 38574 7135 38586 7169
rect 38620 7135 38632 7169
rect 38574 7101 38632 7135
rect 38574 7067 38586 7101
rect 38620 7067 38632 7101
rect 38574 7033 38632 7067
rect 38574 6999 38586 7033
rect 38620 6999 38632 7033
rect 38574 6965 38632 6999
rect 38574 6931 38586 6965
rect 38620 6931 38632 6965
rect 38574 6897 38632 6931
rect 38574 6863 38586 6897
rect 38620 6863 38632 6897
rect 38574 6829 38632 6863
rect 38574 6795 38586 6829
rect 38620 6795 38632 6829
rect 38574 6761 38632 6795
rect 38574 6727 38586 6761
rect 38620 6727 38632 6761
rect 38574 6693 38632 6727
rect 38574 6659 38586 6693
rect 38620 6659 38632 6693
rect 38574 6625 38632 6659
rect 38574 6591 38586 6625
rect 38620 6591 38632 6625
rect 38574 6557 38632 6591
rect 38574 6523 38586 6557
rect 38620 6523 38632 6557
rect 38574 6489 38632 6523
rect 38574 6455 38586 6489
rect 38620 6455 38632 6489
rect 38574 6421 38632 6455
rect 38574 6387 38586 6421
rect 38620 6387 38632 6421
rect 38574 6353 38632 6387
rect 38574 6319 38586 6353
rect 38620 6319 38632 6353
rect 38574 6288 38632 6319
rect 38832 8257 38890 8288
rect 38832 8223 38844 8257
rect 38878 8223 38890 8257
rect 38832 8189 38890 8223
rect 38832 8155 38844 8189
rect 38878 8155 38890 8189
rect 38832 8121 38890 8155
rect 38832 8087 38844 8121
rect 38878 8087 38890 8121
rect 38832 8053 38890 8087
rect 38832 8019 38844 8053
rect 38878 8019 38890 8053
rect 38832 7985 38890 8019
rect 38832 7951 38844 7985
rect 38878 7951 38890 7985
rect 38832 7917 38890 7951
rect 38832 7883 38844 7917
rect 38878 7883 38890 7917
rect 38832 7849 38890 7883
rect 38832 7815 38844 7849
rect 38878 7815 38890 7849
rect 38832 7781 38890 7815
rect 38832 7747 38844 7781
rect 38878 7747 38890 7781
rect 38832 7713 38890 7747
rect 38832 7679 38844 7713
rect 38878 7679 38890 7713
rect 38832 7645 38890 7679
rect 38832 7611 38844 7645
rect 38878 7611 38890 7645
rect 38832 7577 38890 7611
rect 38832 7543 38844 7577
rect 38878 7543 38890 7577
rect 38832 7509 38890 7543
rect 38832 7475 38844 7509
rect 38878 7475 38890 7509
rect 38832 7441 38890 7475
rect 38832 7407 38844 7441
rect 38878 7407 38890 7441
rect 38832 7373 38890 7407
rect 38832 7339 38844 7373
rect 38878 7339 38890 7373
rect 38832 7305 38890 7339
rect 38832 7271 38844 7305
rect 38878 7271 38890 7305
rect 38832 7237 38890 7271
rect 38832 7203 38844 7237
rect 38878 7203 38890 7237
rect 38832 7169 38890 7203
rect 38832 7135 38844 7169
rect 38878 7135 38890 7169
rect 38832 7101 38890 7135
rect 38832 7067 38844 7101
rect 38878 7067 38890 7101
rect 38832 7033 38890 7067
rect 38832 6999 38844 7033
rect 38878 6999 38890 7033
rect 38832 6965 38890 6999
rect 38832 6931 38844 6965
rect 38878 6931 38890 6965
rect 38832 6897 38890 6931
rect 38832 6863 38844 6897
rect 38878 6863 38890 6897
rect 38832 6829 38890 6863
rect 38832 6795 38844 6829
rect 38878 6795 38890 6829
rect 38832 6761 38890 6795
rect 38832 6727 38844 6761
rect 38878 6727 38890 6761
rect 38832 6693 38890 6727
rect 38832 6659 38844 6693
rect 38878 6659 38890 6693
rect 38832 6625 38890 6659
rect 38832 6591 38844 6625
rect 38878 6591 38890 6625
rect 38832 6557 38890 6591
rect 38832 6523 38844 6557
rect 38878 6523 38890 6557
rect 38832 6489 38890 6523
rect 38832 6455 38844 6489
rect 38878 6455 38890 6489
rect 38832 6421 38890 6455
rect 38832 6387 38844 6421
rect 38878 6387 38890 6421
rect 38832 6353 38890 6387
rect 38832 6319 38844 6353
rect 38878 6319 38890 6353
rect 38832 6288 38890 6319
rect 39090 8257 39148 8288
rect 39090 8223 39102 8257
rect 39136 8223 39148 8257
rect 39090 8189 39148 8223
rect 39090 8155 39102 8189
rect 39136 8155 39148 8189
rect 39090 8121 39148 8155
rect 39090 8087 39102 8121
rect 39136 8087 39148 8121
rect 39090 8053 39148 8087
rect 39090 8019 39102 8053
rect 39136 8019 39148 8053
rect 39090 7985 39148 8019
rect 39090 7951 39102 7985
rect 39136 7951 39148 7985
rect 39090 7917 39148 7951
rect 39090 7883 39102 7917
rect 39136 7883 39148 7917
rect 39090 7849 39148 7883
rect 39090 7815 39102 7849
rect 39136 7815 39148 7849
rect 39090 7781 39148 7815
rect 39090 7747 39102 7781
rect 39136 7747 39148 7781
rect 39090 7713 39148 7747
rect 39090 7679 39102 7713
rect 39136 7679 39148 7713
rect 39090 7645 39148 7679
rect 39090 7611 39102 7645
rect 39136 7611 39148 7645
rect 39090 7577 39148 7611
rect 39090 7543 39102 7577
rect 39136 7543 39148 7577
rect 39090 7509 39148 7543
rect 39090 7475 39102 7509
rect 39136 7475 39148 7509
rect 39090 7441 39148 7475
rect 39090 7407 39102 7441
rect 39136 7407 39148 7441
rect 39090 7373 39148 7407
rect 39090 7339 39102 7373
rect 39136 7339 39148 7373
rect 39090 7305 39148 7339
rect 39090 7271 39102 7305
rect 39136 7271 39148 7305
rect 39090 7237 39148 7271
rect 39090 7203 39102 7237
rect 39136 7203 39148 7237
rect 39090 7169 39148 7203
rect 39090 7135 39102 7169
rect 39136 7135 39148 7169
rect 39090 7101 39148 7135
rect 39090 7067 39102 7101
rect 39136 7067 39148 7101
rect 39090 7033 39148 7067
rect 39090 6999 39102 7033
rect 39136 6999 39148 7033
rect 39090 6965 39148 6999
rect 39090 6931 39102 6965
rect 39136 6931 39148 6965
rect 39090 6897 39148 6931
rect 39090 6863 39102 6897
rect 39136 6863 39148 6897
rect 39090 6829 39148 6863
rect 39090 6795 39102 6829
rect 39136 6795 39148 6829
rect 39090 6761 39148 6795
rect 39090 6727 39102 6761
rect 39136 6727 39148 6761
rect 39090 6693 39148 6727
rect 39090 6659 39102 6693
rect 39136 6659 39148 6693
rect 39090 6625 39148 6659
rect 39090 6591 39102 6625
rect 39136 6591 39148 6625
rect 39090 6557 39148 6591
rect 39090 6523 39102 6557
rect 39136 6523 39148 6557
rect 39090 6489 39148 6523
rect 39090 6455 39102 6489
rect 39136 6455 39148 6489
rect 39090 6421 39148 6455
rect 39090 6387 39102 6421
rect 39136 6387 39148 6421
rect 39090 6353 39148 6387
rect 39090 6319 39102 6353
rect 39136 6319 39148 6353
rect 39090 6288 39148 6319
rect 39348 8257 39406 8288
rect 39348 8223 39360 8257
rect 39394 8223 39406 8257
rect 39348 8189 39406 8223
rect 39348 8155 39360 8189
rect 39394 8155 39406 8189
rect 39348 8121 39406 8155
rect 39348 8087 39360 8121
rect 39394 8087 39406 8121
rect 39348 8053 39406 8087
rect 39348 8019 39360 8053
rect 39394 8019 39406 8053
rect 39348 7985 39406 8019
rect 39348 7951 39360 7985
rect 39394 7951 39406 7985
rect 39348 7917 39406 7951
rect 39348 7883 39360 7917
rect 39394 7883 39406 7917
rect 39348 7849 39406 7883
rect 39348 7815 39360 7849
rect 39394 7815 39406 7849
rect 39348 7781 39406 7815
rect 39348 7747 39360 7781
rect 39394 7747 39406 7781
rect 39348 7713 39406 7747
rect 39348 7679 39360 7713
rect 39394 7679 39406 7713
rect 39348 7645 39406 7679
rect 39348 7611 39360 7645
rect 39394 7611 39406 7645
rect 39348 7577 39406 7611
rect 39348 7543 39360 7577
rect 39394 7543 39406 7577
rect 39348 7509 39406 7543
rect 39348 7475 39360 7509
rect 39394 7475 39406 7509
rect 39348 7441 39406 7475
rect 39348 7407 39360 7441
rect 39394 7407 39406 7441
rect 39348 7373 39406 7407
rect 39348 7339 39360 7373
rect 39394 7339 39406 7373
rect 39348 7305 39406 7339
rect 39348 7271 39360 7305
rect 39394 7271 39406 7305
rect 39348 7237 39406 7271
rect 39348 7203 39360 7237
rect 39394 7203 39406 7237
rect 39348 7169 39406 7203
rect 39348 7135 39360 7169
rect 39394 7135 39406 7169
rect 39348 7101 39406 7135
rect 39348 7067 39360 7101
rect 39394 7067 39406 7101
rect 39348 7033 39406 7067
rect 39348 6999 39360 7033
rect 39394 6999 39406 7033
rect 39348 6965 39406 6999
rect 39348 6931 39360 6965
rect 39394 6931 39406 6965
rect 39348 6897 39406 6931
rect 39348 6863 39360 6897
rect 39394 6863 39406 6897
rect 39348 6829 39406 6863
rect 39348 6795 39360 6829
rect 39394 6795 39406 6829
rect 39348 6761 39406 6795
rect 39348 6727 39360 6761
rect 39394 6727 39406 6761
rect 39348 6693 39406 6727
rect 39348 6659 39360 6693
rect 39394 6659 39406 6693
rect 39348 6625 39406 6659
rect 39348 6591 39360 6625
rect 39394 6591 39406 6625
rect 39348 6557 39406 6591
rect 39348 6523 39360 6557
rect 39394 6523 39406 6557
rect 39348 6489 39406 6523
rect 39348 6455 39360 6489
rect 39394 6455 39406 6489
rect 39348 6421 39406 6455
rect 39348 6387 39360 6421
rect 39394 6387 39406 6421
rect 39348 6353 39406 6387
rect 39348 6319 39360 6353
rect 39394 6319 39406 6353
rect 39348 6288 39406 6319
rect 39606 8257 39664 8288
rect 39606 8223 39618 8257
rect 39652 8223 39664 8257
rect 39606 8189 39664 8223
rect 39606 8155 39618 8189
rect 39652 8155 39664 8189
rect 39606 8121 39664 8155
rect 39606 8087 39618 8121
rect 39652 8087 39664 8121
rect 39606 8053 39664 8087
rect 39606 8019 39618 8053
rect 39652 8019 39664 8053
rect 39606 7985 39664 8019
rect 39606 7951 39618 7985
rect 39652 7951 39664 7985
rect 39606 7917 39664 7951
rect 39606 7883 39618 7917
rect 39652 7883 39664 7917
rect 39606 7849 39664 7883
rect 39606 7815 39618 7849
rect 39652 7815 39664 7849
rect 39606 7781 39664 7815
rect 39606 7747 39618 7781
rect 39652 7747 39664 7781
rect 39606 7713 39664 7747
rect 39606 7679 39618 7713
rect 39652 7679 39664 7713
rect 39606 7645 39664 7679
rect 39606 7611 39618 7645
rect 39652 7611 39664 7645
rect 39606 7577 39664 7611
rect 39606 7543 39618 7577
rect 39652 7543 39664 7577
rect 39606 7509 39664 7543
rect 39606 7475 39618 7509
rect 39652 7475 39664 7509
rect 39606 7441 39664 7475
rect 39606 7407 39618 7441
rect 39652 7407 39664 7441
rect 39606 7373 39664 7407
rect 39606 7339 39618 7373
rect 39652 7339 39664 7373
rect 39606 7305 39664 7339
rect 39606 7271 39618 7305
rect 39652 7271 39664 7305
rect 39606 7237 39664 7271
rect 39606 7203 39618 7237
rect 39652 7203 39664 7237
rect 39606 7169 39664 7203
rect 39606 7135 39618 7169
rect 39652 7135 39664 7169
rect 39606 7101 39664 7135
rect 39606 7067 39618 7101
rect 39652 7067 39664 7101
rect 39606 7033 39664 7067
rect 39606 6999 39618 7033
rect 39652 6999 39664 7033
rect 39606 6965 39664 6999
rect 39606 6931 39618 6965
rect 39652 6931 39664 6965
rect 39606 6897 39664 6931
rect 39606 6863 39618 6897
rect 39652 6863 39664 6897
rect 39606 6829 39664 6863
rect 39606 6795 39618 6829
rect 39652 6795 39664 6829
rect 39606 6761 39664 6795
rect 39606 6727 39618 6761
rect 39652 6727 39664 6761
rect 39606 6693 39664 6727
rect 39606 6659 39618 6693
rect 39652 6659 39664 6693
rect 39606 6625 39664 6659
rect 39606 6591 39618 6625
rect 39652 6591 39664 6625
rect 39606 6557 39664 6591
rect 39606 6523 39618 6557
rect 39652 6523 39664 6557
rect 39606 6489 39664 6523
rect 39606 6455 39618 6489
rect 39652 6455 39664 6489
rect 39606 6421 39664 6455
rect 39606 6387 39618 6421
rect 39652 6387 39664 6421
rect 39606 6353 39664 6387
rect 39606 6319 39618 6353
rect 39652 6319 39664 6353
rect 39606 6288 39664 6319
rect 39864 8257 39922 8288
rect 39864 8223 39876 8257
rect 39910 8223 39922 8257
rect 39864 8189 39922 8223
rect 39864 8155 39876 8189
rect 39910 8155 39922 8189
rect 39864 8121 39922 8155
rect 39864 8087 39876 8121
rect 39910 8087 39922 8121
rect 39864 8053 39922 8087
rect 39864 8019 39876 8053
rect 39910 8019 39922 8053
rect 39864 7985 39922 8019
rect 39864 7951 39876 7985
rect 39910 7951 39922 7985
rect 39864 7917 39922 7951
rect 39864 7883 39876 7917
rect 39910 7883 39922 7917
rect 39864 7849 39922 7883
rect 39864 7815 39876 7849
rect 39910 7815 39922 7849
rect 39864 7781 39922 7815
rect 39864 7747 39876 7781
rect 39910 7747 39922 7781
rect 39864 7713 39922 7747
rect 39864 7679 39876 7713
rect 39910 7679 39922 7713
rect 39864 7645 39922 7679
rect 39864 7611 39876 7645
rect 39910 7611 39922 7645
rect 39864 7577 39922 7611
rect 39864 7543 39876 7577
rect 39910 7543 39922 7577
rect 39864 7509 39922 7543
rect 39864 7475 39876 7509
rect 39910 7475 39922 7509
rect 39864 7441 39922 7475
rect 39864 7407 39876 7441
rect 39910 7407 39922 7441
rect 39864 7373 39922 7407
rect 39864 7339 39876 7373
rect 39910 7339 39922 7373
rect 39864 7305 39922 7339
rect 39864 7271 39876 7305
rect 39910 7271 39922 7305
rect 39864 7237 39922 7271
rect 39864 7203 39876 7237
rect 39910 7203 39922 7237
rect 39864 7169 39922 7203
rect 39864 7135 39876 7169
rect 39910 7135 39922 7169
rect 39864 7101 39922 7135
rect 39864 7067 39876 7101
rect 39910 7067 39922 7101
rect 39864 7033 39922 7067
rect 39864 6999 39876 7033
rect 39910 6999 39922 7033
rect 39864 6965 39922 6999
rect 39864 6931 39876 6965
rect 39910 6931 39922 6965
rect 39864 6897 39922 6931
rect 39864 6863 39876 6897
rect 39910 6863 39922 6897
rect 39864 6829 39922 6863
rect 39864 6795 39876 6829
rect 39910 6795 39922 6829
rect 39864 6761 39922 6795
rect 39864 6727 39876 6761
rect 39910 6727 39922 6761
rect 39864 6693 39922 6727
rect 39864 6659 39876 6693
rect 39910 6659 39922 6693
rect 39864 6625 39922 6659
rect 39864 6591 39876 6625
rect 39910 6591 39922 6625
rect 39864 6557 39922 6591
rect 39864 6523 39876 6557
rect 39910 6523 39922 6557
rect 39864 6489 39922 6523
rect 39864 6455 39876 6489
rect 39910 6455 39922 6489
rect 39864 6421 39922 6455
rect 39864 6387 39876 6421
rect 39910 6387 39922 6421
rect 39864 6353 39922 6387
rect 39864 6319 39876 6353
rect 39910 6319 39922 6353
rect 39864 6288 39922 6319
rect 40122 8257 40180 8288
rect 40122 8223 40134 8257
rect 40168 8223 40180 8257
rect 40122 8189 40180 8223
rect 40122 8155 40134 8189
rect 40168 8155 40180 8189
rect 40122 8121 40180 8155
rect 40122 8087 40134 8121
rect 40168 8087 40180 8121
rect 40122 8053 40180 8087
rect 40122 8019 40134 8053
rect 40168 8019 40180 8053
rect 40122 7985 40180 8019
rect 40122 7951 40134 7985
rect 40168 7951 40180 7985
rect 40122 7917 40180 7951
rect 40122 7883 40134 7917
rect 40168 7883 40180 7917
rect 40122 7849 40180 7883
rect 40122 7815 40134 7849
rect 40168 7815 40180 7849
rect 40122 7781 40180 7815
rect 40122 7747 40134 7781
rect 40168 7747 40180 7781
rect 40122 7713 40180 7747
rect 40122 7679 40134 7713
rect 40168 7679 40180 7713
rect 40122 7645 40180 7679
rect 40122 7611 40134 7645
rect 40168 7611 40180 7645
rect 40122 7577 40180 7611
rect 40122 7543 40134 7577
rect 40168 7543 40180 7577
rect 40122 7509 40180 7543
rect 40122 7475 40134 7509
rect 40168 7475 40180 7509
rect 40122 7441 40180 7475
rect 40122 7407 40134 7441
rect 40168 7407 40180 7441
rect 40122 7373 40180 7407
rect 40122 7339 40134 7373
rect 40168 7339 40180 7373
rect 40122 7305 40180 7339
rect 40122 7271 40134 7305
rect 40168 7271 40180 7305
rect 40122 7237 40180 7271
rect 40122 7203 40134 7237
rect 40168 7203 40180 7237
rect 40122 7169 40180 7203
rect 40122 7135 40134 7169
rect 40168 7135 40180 7169
rect 40122 7101 40180 7135
rect 40122 7067 40134 7101
rect 40168 7067 40180 7101
rect 40122 7033 40180 7067
rect 40122 6999 40134 7033
rect 40168 6999 40180 7033
rect 40122 6965 40180 6999
rect 40122 6931 40134 6965
rect 40168 6931 40180 6965
rect 40122 6897 40180 6931
rect 40122 6863 40134 6897
rect 40168 6863 40180 6897
rect 40122 6829 40180 6863
rect 40122 6795 40134 6829
rect 40168 6795 40180 6829
rect 40122 6761 40180 6795
rect 40122 6727 40134 6761
rect 40168 6727 40180 6761
rect 40122 6693 40180 6727
rect 40122 6659 40134 6693
rect 40168 6659 40180 6693
rect 40122 6625 40180 6659
rect 40122 6591 40134 6625
rect 40168 6591 40180 6625
rect 40122 6557 40180 6591
rect 40122 6523 40134 6557
rect 40168 6523 40180 6557
rect 40122 6489 40180 6523
rect 40122 6455 40134 6489
rect 40168 6455 40180 6489
rect 40122 6421 40180 6455
rect 40122 6387 40134 6421
rect 40168 6387 40180 6421
rect 40122 6353 40180 6387
rect 40122 6319 40134 6353
rect 40168 6319 40180 6353
rect 40122 6288 40180 6319
rect 40380 8257 40438 8288
rect 40380 8223 40392 8257
rect 40426 8223 40438 8257
rect 40380 8189 40438 8223
rect 40380 8155 40392 8189
rect 40426 8155 40438 8189
rect 40380 8121 40438 8155
rect 40380 8087 40392 8121
rect 40426 8087 40438 8121
rect 40380 8053 40438 8087
rect 40380 8019 40392 8053
rect 40426 8019 40438 8053
rect 40380 7985 40438 8019
rect 40380 7951 40392 7985
rect 40426 7951 40438 7985
rect 40380 7917 40438 7951
rect 40380 7883 40392 7917
rect 40426 7883 40438 7917
rect 40380 7849 40438 7883
rect 40380 7815 40392 7849
rect 40426 7815 40438 7849
rect 40380 7781 40438 7815
rect 40380 7747 40392 7781
rect 40426 7747 40438 7781
rect 40380 7713 40438 7747
rect 40380 7679 40392 7713
rect 40426 7679 40438 7713
rect 40380 7645 40438 7679
rect 40380 7611 40392 7645
rect 40426 7611 40438 7645
rect 40380 7577 40438 7611
rect 40380 7543 40392 7577
rect 40426 7543 40438 7577
rect 40380 7509 40438 7543
rect 40380 7475 40392 7509
rect 40426 7475 40438 7509
rect 40380 7441 40438 7475
rect 40380 7407 40392 7441
rect 40426 7407 40438 7441
rect 40380 7373 40438 7407
rect 40380 7339 40392 7373
rect 40426 7339 40438 7373
rect 40380 7305 40438 7339
rect 40380 7271 40392 7305
rect 40426 7271 40438 7305
rect 40380 7237 40438 7271
rect 40380 7203 40392 7237
rect 40426 7203 40438 7237
rect 40380 7169 40438 7203
rect 40380 7135 40392 7169
rect 40426 7135 40438 7169
rect 40380 7101 40438 7135
rect 40380 7067 40392 7101
rect 40426 7067 40438 7101
rect 40380 7033 40438 7067
rect 40380 6999 40392 7033
rect 40426 6999 40438 7033
rect 40380 6965 40438 6999
rect 40380 6931 40392 6965
rect 40426 6931 40438 6965
rect 40380 6897 40438 6931
rect 40380 6863 40392 6897
rect 40426 6863 40438 6897
rect 40380 6829 40438 6863
rect 40380 6795 40392 6829
rect 40426 6795 40438 6829
rect 40380 6761 40438 6795
rect 40380 6727 40392 6761
rect 40426 6727 40438 6761
rect 40380 6693 40438 6727
rect 40380 6659 40392 6693
rect 40426 6659 40438 6693
rect 40380 6625 40438 6659
rect 40380 6591 40392 6625
rect 40426 6591 40438 6625
rect 40380 6557 40438 6591
rect 40380 6523 40392 6557
rect 40426 6523 40438 6557
rect 40380 6489 40438 6523
rect 40380 6455 40392 6489
rect 40426 6455 40438 6489
rect 40380 6421 40438 6455
rect 40380 6387 40392 6421
rect 40426 6387 40438 6421
rect 40380 6353 40438 6387
rect 40380 6319 40392 6353
rect 40426 6319 40438 6353
rect 40380 6288 40438 6319
rect 40638 8257 40696 8288
rect 40638 8223 40650 8257
rect 40684 8223 40696 8257
rect 40638 8189 40696 8223
rect 40638 8155 40650 8189
rect 40684 8155 40696 8189
rect 40638 8121 40696 8155
rect 40638 8087 40650 8121
rect 40684 8087 40696 8121
rect 40638 8053 40696 8087
rect 40638 8019 40650 8053
rect 40684 8019 40696 8053
rect 40638 7985 40696 8019
rect 40638 7951 40650 7985
rect 40684 7951 40696 7985
rect 40638 7917 40696 7951
rect 40638 7883 40650 7917
rect 40684 7883 40696 7917
rect 40638 7849 40696 7883
rect 40638 7815 40650 7849
rect 40684 7815 40696 7849
rect 40638 7781 40696 7815
rect 40638 7747 40650 7781
rect 40684 7747 40696 7781
rect 40638 7713 40696 7747
rect 40638 7679 40650 7713
rect 40684 7679 40696 7713
rect 40638 7645 40696 7679
rect 40638 7611 40650 7645
rect 40684 7611 40696 7645
rect 40638 7577 40696 7611
rect 40638 7543 40650 7577
rect 40684 7543 40696 7577
rect 40638 7509 40696 7543
rect 40638 7475 40650 7509
rect 40684 7475 40696 7509
rect 40638 7441 40696 7475
rect 40638 7407 40650 7441
rect 40684 7407 40696 7441
rect 40638 7373 40696 7407
rect 40638 7339 40650 7373
rect 40684 7339 40696 7373
rect 40638 7305 40696 7339
rect 40638 7271 40650 7305
rect 40684 7271 40696 7305
rect 40638 7237 40696 7271
rect 40638 7203 40650 7237
rect 40684 7203 40696 7237
rect 40638 7169 40696 7203
rect 40638 7135 40650 7169
rect 40684 7135 40696 7169
rect 40638 7101 40696 7135
rect 40638 7067 40650 7101
rect 40684 7067 40696 7101
rect 40638 7033 40696 7067
rect 40638 6999 40650 7033
rect 40684 6999 40696 7033
rect 40638 6965 40696 6999
rect 40638 6931 40650 6965
rect 40684 6931 40696 6965
rect 40638 6897 40696 6931
rect 40638 6863 40650 6897
rect 40684 6863 40696 6897
rect 40638 6829 40696 6863
rect 40638 6795 40650 6829
rect 40684 6795 40696 6829
rect 40638 6761 40696 6795
rect 40638 6727 40650 6761
rect 40684 6727 40696 6761
rect 40638 6693 40696 6727
rect 40638 6659 40650 6693
rect 40684 6659 40696 6693
rect 40638 6625 40696 6659
rect 40638 6591 40650 6625
rect 40684 6591 40696 6625
rect 40638 6557 40696 6591
rect 40638 6523 40650 6557
rect 40684 6523 40696 6557
rect 40638 6489 40696 6523
rect 40638 6455 40650 6489
rect 40684 6455 40696 6489
rect 40638 6421 40696 6455
rect 40638 6387 40650 6421
rect 40684 6387 40696 6421
rect 40638 6353 40696 6387
rect 40638 6319 40650 6353
rect 40684 6319 40696 6353
rect 40638 6288 40696 6319
rect 40896 8257 40954 8288
rect 40896 8223 40908 8257
rect 40942 8223 40954 8257
rect 40896 8189 40954 8223
rect 40896 8155 40908 8189
rect 40942 8155 40954 8189
rect 40896 8121 40954 8155
rect 40896 8087 40908 8121
rect 40942 8087 40954 8121
rect 40896 8053 40954 8087
rect 40896 8019 40908 8053
rect 40942 8019 40954 8053
rect 40896 7985 40954 8019
rect 40896 7951 40908 7985
rect 40942 7951 40954 7985
rect 40896 7917 40954 7951
rect 40896 7883 40908 7917
rect 40942 7883 40954 7917
rect 40896 7849 40954 7883
rect 40896 7815 40908 7849
rect 40942 7815 40954 7849
rect 40896 7781 40954 7815
rect 40896 7747 40908 7781
rect 40942 7747 40954 7781
rect 40896 7713 40954 7747
rect 40896 7679 40908 7713
rect 40942 7679 40954 7713
rect 40896 7645 40954 7679
rect 40896 7611 40908 7645
rect 40942 7611 40954 7645
rect 40896 7577 40954 7611
rect 40896 7543 40908 7577
rect 40942 7543 40954 7577
rect 40896 7509 40954 7543
rect 40896 7475 40908 7509
rect 40942 7475 40954 7509
rect 40896 7441 40954 7475
rect 40896 7407 40908 7441
rect 40942 7407 40954 7441
rect 40896 7373 40954 7407
rect 40896 7339 40908 7373
rect 40942 7339 40954 7373
rect 40896 7305 40954 7339
rect 40896 7271 40908 7305
rect 40942 7271 40954 7305
rect 40896 7237 40954 7271
rect 40896 7203 40908 7237
rect 40942 7203 40954 7237
rect 40896 7169 40954 7203
rect 40896 7135 40908 7169
rect 40942 7135 40954 7169
rect 40896 7101 40954 7135
rect 40896 7067 40908 7101
rect 40942 7067 40954 7101
rect 40896 7033 40954 7067
rect 40896 6999 40908 7033
rect 40942 6999 40954 7033
rect 40896 6965 40954 6999
rect 40896 6931 40908 6965
rect 40942 6931 40954 6965
rect 40896 6897 40954 6931
rect 40896 6863 40908 6897
rect 40942 6863 40954 6897
rect 40896 6829 40954 6863
rect 40896 6795 40908 6829
rect 40942 6795 40954 6829
rect 40896 6761 40954 6795
rect 40896 6727 40908 6761
rect 40942 6727 40954 6761
rect 40896 6693 40954 6727
rect 40896 6659 40908 6693
rect 40942 6659 40954 6693
rect 40896 6625 40954 6659
rect 40896 6591 40908 6625
rect 40942 6591 40954 6625
rect 40896 6557 40954 6591
rect 40896 6523 40908 6557
rect 40942 6523 40954 6557
rect 40896 6489 40954 6523
rect 40896 6455 40908 6489
rect 40942 6455 40954 6489
rect 40896 6421 40954 6455
rect 40896 6387 40908 6421
rect 40942 6387 40954 6421
rect 40896 6353 40954 6387
rect 40896 6319 40908 6353
rect 40942 6319 40954 6353
rect 40896 6288 40954 6319
rect 41154 8257 41212 8288
rect 41154 8223 41166 8257
rect 41200 8223 41212 8257
rect 41154 8189 41212 8223
rect 41154 8155 41166 8189
rect 41200 8155 41212 8189
rect 41154 8121 41212 8155
rect 41154 8087 41166 8121
rect 41200 8087 41212 8121
rect 41154 8053 41212 8087
rect 41154 8019 41166 8053
rect 41200 8019 41212 8053
rect 41154 7985 41212 8019
rect 41154 7951 41166 7985
rect 41200 7951 41212 7985
rect 41154 7917 41212 7951
rect 41154 7883 41166 7917
rect 41200 7883 41212 7917
rect 41154 7849 41212 7883
rect 41154 7815 41166 7849
rect 41200 7815 41212 7849
rect 41154 7781 41212 7815
rect 41154 7747 41166 7781
rect 41200 7747 41212 7781
rect 41154 7713 41212 7747
rect 41154 7679 41166 7713
rect 41200 7679 41212 7713
rect 41154 7645 41212 7679
rect 41154 7611 41166 7645
rect 41200 7611 41212 7645
rect 41154 7577 41212 7611
rect 41154 7543 41166 7577
rect 41200 7543 41212 7577
rect 41154 7509 41212 7543
rect 41154 7475 41166 7509
rect 41200 7475 41212 7509
rect 41154 7441 41212 7475
rect 41154 7407 41166 7441
rect 41200 7407 41212 7441
rect 41154 7373 41212 7407
rect 41154 7339 41166 7373
rect 41200 7339 41212 7373
rect 41154 7305 41212 7339
rect 41154 7271 41166 7305
rect 41200 7271 41212 7305
rect 41154 7237 41212 7271
rect 41154 7203 41166 7237
rect 41200 7203 41212 7237
rect 41154 7169 41212 7203
rect 41154 7135 41166 7169
rect 41200 7135 41212 7169
rect 41154 7101 41212 7135
rect 41154 7067 41166 7101
rect 41200 7067 41212 7101
rect 41154 7033 41212 7067
rect 41154 6999 41166 7033
rect 41200 6999 41212 7033
rect 41154 6965 41212 6999
rect 41154 6931 41166 6965
rect 41200 6931 41212 6965
rect 41154 6897 41212 6931
rect 41154 6863 41166 6897
rect 41200 6863 41212 6897
rect 41154 6829 41212 6863
rect 41154 6795 41166 6829
rect 41200 6795 41212 6829
rect 41154 6761 41212 6795
rect 41154 6727 41166 6761
rect 41200 6727 41212 6761
rect 41154 6693 41212 6727
rect 41154 6659 41166 6693
rect 41200 6659 41212 6693
rect 41154 6625 41212 6659
rect 41154 6591 41166 6625
rect 41200 6591 41212 6625
rect 41154 6557 41212 6591
rect 41154 6523 41166 6557
rect 41200 6523 41212 6557
rect 41154 6489 41212 6523
rect 41154 6455 41166 6489
rect 41200 6455 41212 6489
rect 41154 6421 41212 6455
rect 41154 6387 41166 6421
rect 41200 6387 41212 6421
rect 41154 6353 41212 6387
rect 41154 6319 41166 6353
rect 41200 6319 41212 6353
rect 41154 6288 41212 6319
rect 41412 8257 41470 8288
rect 41412 8223 41424 8257
rect 41458 8223 41470 8257
rect 41412 8189 41470 8223
rect 41412 8155 41424 8189
rect 41458 8155 41470 8189
rect 41412 8121 41470 8155
rect 41412 8087 41424 8121
rect 41458 8087 41470 8121
rect 41412 8053 41470 8087
rect 41412 8019 41424 8053
rect 41458 8019 41470 8053
rect 41412 7985 41470 8019
rect 41412 7951 41424 7985
rect 41458 7951 41470 7985
rect 41412 7917 41470 7951
rect 41412 7883 41424 7917
rect 41458 7883 41470 7917
rect 41412 7849 41470 7883
rect 41412 7815 41424 7849
rect 41458 7815 41470 7849
rect 41412 7781 41470 7815
rect 41412 7747 41424 7781
rect 41458 7747 41470 7781
rect 41412 7713 41470 7747
rect 41412 7679 41424 7713
rect 41458 7679 41470 7713
rect 41412 7645 41470 7679
rect 41412 7611 41424 7645
rect 41458 7611 41470 7645
rect 41412 7577 41470 7611
rect 41412 7543 41424 7577
rect 41458 7543 41470 7577
rect 41412 7509 41470 7543
rect 41412 7475 41424 7509
rect 41458 7475 41470 7509
rect 41412 7441 41470 7475
rect 41412 7407 41424 7441
rect 41458 7407 41470 7441
rect 41412 7373 41470 7407
rect 41412 7339 41424 7373
rect 41458 7339 41470 7373
rect 41412 7305 41470 7339
rect 41412 7271 41424 7305
rect 41458 7271 41470 7305
rect 41412 7237 41470 7271
rect 41412 7203 41424 7237
rect 41458 7203 41470 7237
rect 41412 7169 41470 7203
rect 41412 7135 41424 7169
rect 41458 7135 41470 7169
rect 41412 7101 41470 7135
rect 41412 7067 41424 7101
rect 41458 7067 41470 7101
rect 41412 7033 41470 7067
rect 41412 6999 41424 7033
rect 41458 6999 41470 7033
rect 41412 6965 41470 6999
rect 41412 6931 41424 6965
rect 41458 6931 41470 6965
rect 41412 6897 41470 6931
rect 41412 6863 41424 6897
rect 41458 6863 41470 6897
rect 41412 6829 41470 6863
rect 41412 6795 41424 6829
rect 41458 6795 41470 6829
rect 41412 6761 41470 6795
rect 41412 6727 41424 6761
rect 41458 6727 41470 6761
rect 41412 6693 41470 6727
rect 41412 6659 41424 6693
rect 41458 6659 41470 6693
rect 41412 6625 41470 6659
rect 41412 6591 41424 6625
rect 41458 6591 41470 6625
rect 41412 6557 41470 6591
rect 41412 6523 41424 6557
rect 41458 6523 41470 6557
rect 41412 6489 41470 6523
rect 41412 6455 41424 6489
rect 41458 6455 41470 6489
rect 41412 6421 41470 6455
rect 41412 6387 41424 6421
rect 41458 6387 41470 6421
rect 41412 6353 41470 6387
rect 41412 6319 41424 6353
rect 41458 6319 41470 6353
rect 41412 6288 41470 6319
rect 41670 8257 41728 8288
rect 41670 8223 41682 8257
rect 41716 8223 41728 8257
rect 41670 8189 41728 8223
rect 41670 8155 41682 8189
rect 41716 8155 41728 8189
rect 41670 8121 41728 8155
rect 41670 8087 41682 8121
rect 41716 8087 41728 8121
rect 41670 8053 41728 8087
rect 41670 8019 41682 8053
rect 41716 8019 41728 8053
rect 41670 7985 41728 8019
rect 41670 7951 41682 7985
rect 41716 7951 41728 7985
rect 41670 7917 41728 7951
rect 41670 7883 41682 7917
rect 41716 7883 41728 7917
rect 41670 7849 41728 7883
rect 41670 7815 41682 7849
rect 41716 7815 41728 7849
rect 41670 7781 41728 7815
rect 41670 7747 41682 7781
rect 41716 7747 41728 7781
rect 41670 7713 41728 7747
rect 41670 7679 41682 7713
rect 41716 7679 41728 7713
rect 41670 7645 41728 7679
rect 41670 7611 41682 7645
rect 41716 7611 41728 7645
rect 41670 7577 41728 7611
rect 41670 7543 41682 7577
rect 41716 7543 41728 7577
rect 41670 7509 41728 7543
rect 41670 7475 41682 7509
rect 41716 7475 41728 7509
rect 41670 7441 41728 7475
rect 41670 7407 41682 7441
rect 41716 7407 41728 7441
rect 41670 7373 41728 7407
rect 41670 7339 41682 7373
rect 41716 7339 41728 7373
rect 41670 7305 41728 7339
rect 41670 7271 41682 7305
rect 41716 7271 41728 7305
rect 41670 7237 41728 7271
rect 41670 7203 41682 7237
rect 41716 7203 41728 7237
rect 41670 7169 41728 7203
rect 41670 7135 41682 7169
rect 41716 7135 41728 7169
rect 41670 7101 41728 7135
rect 41670 7067 41682 7101
rect 41716 7067 41728 7101
rect 41670 7033 41728 7067
rect 41670 6999 41682 7033
rect 41716 6999 41728 7033
rect 41670 6965 41728 6999
rect 41670 6931 41682 6965
rect 41716 6931 41728 6965
rect 41670 6897 41728 6931
rect 41670 6863 41682 6897
rect 41716 6863 41728 6897
rect 41670 6829 41728 6863
rect 41670 6795 41682 6829
rect 41716 6795 41728 6829
rect 41670 6761 41728 6795
rect 41670 6727 41682 6761
rect 41716 6727 41728 6761
rect 41670 6693 41728 6727
rect 41670 6659 41682 6693
rect 41716 6659 41728 6693
rect 41670 6625 41728 6659
rect 41670 6591 41682 6625
rect 41716 6591 41728 6625
rect 41670 6557 41728 6591
rect 41670 6523 41682 6557
rect 41716 6523 41728 6557
rect 41670 6489 41728 6523
rect 41670 6455 41682 6489
rect 41716 6455 41728 6489
rect 41670 6421 41728 6455
rect 41670 6387 41682 6421
rect 41716 6387 41728 6421
rect 41670 6353 41728 6387
rect 41670 6319 41682 6353
rect 41716 6319 41728 6353
rect 41670 6288 41728 6319
rect 41928 8257 41986 8288
rect 41928 8223 41940 8257
rect 41974 8223 41986 8257
rect 41928 8189 41986 8223
rect 41928 8155 41940 8189
rect 41974 8155 41986 8189
rect 41928 8121 41986 8155
rect 41928 8087 41940 8121
rect 41974 8087 41986 8121
rect 41928 8053 41986 8087
rect 41928 8019 41940 8053
rect 41974 8019 41986 8053
rect 41928 7985 41986 8019
rect 41928 7951 41940 7985
rect 41974 7951 41986 7985
rect 41928 7917 41986 7951
rect 41928 7883 41940 7917
rect 41974 7883 41986 7917
rect 41928 7849 41986 7883
rect 41928 7815 41940 7849
rect 41974 7815 41986 7849
rect 41928 7781 41986 7815
rect 41928 7747 41940 7781
rect 41974 7747 41986 7781
rect 41928 7713 41986 7747
rect 41928 7679 41940 7713
rect 41974 7679 41986 7713
rect 41928 7645 41986 7679
rect 41928 7611 41940 7645
rect 41974 7611 41986 7645
rect 41928 7577 41986 7611
rect 41928 7543 41940 7577
rect 41974 7543 41986 7577
rect 41928 7509 41986 7543
rect 41928 7475 41940 7509
rect 41974 7475 41986 7509
rect 41928 7441 41986 7475
rect 41928 7407 41940 7441
rect 41974 7407 41986 7441
rect 41928 7373 41986 7407
rect 41928 7339 41940 7373
rect 41974 7339 41986 7373
rect 41928 7305 41986 7339
rect 41928 7271 41940 7305
rect 41974 7271 41986 7305
rect 41928 7237 41986 7271
rect 41928 7203 41940 7237
rect 41974 7203 41986 7237
rect 41928 7169 41986 7203
rect 41928 7135 41940 7169
rect 41974 7135 41986 7169
rect 41928 7101 41986 7135
rect 41928 7067 41940 7101
rect 41974 7067 41986 7101
rect 41928 7033 41986 7067
rect 41928 6999 41940 7033
rect 41974 6999 41986 7033
rect 41928 6965 41986 6999
rect 41928 6931 41940 6965
rect 41974 6931 41986 6965
rect 41928 6897 41986 6931
rect 41928 6863 41940 6897
rect 41974 6863 41986 6897
rect 41928 6829 41986 6863
rect 41928 6795 41940 6829
rect 41974 6795 41986 6829
rect 41928 6761 41986 6795
rect 41928 6727 41940 6761
rect 41974 6727 41986 6761
rect 41928 6693 41986 6727
rect 41928 6659 41940 6693
rect 41974 6659 41986 6693
rect 41928 6625 41986 6659
rect 41928 6591 41940 6625
rect 41974 6591 41986 6625
rect 41928 6557 41986 6591
rect 41928 6523 41940 6557
rect 41974 6523 41986 6557
rect 41928 6489 41986 6523
rect 41928 6455 41940 6489
rect 41974 6455 41986 6489
rect 41928 6421 41986 6455
rect 41928 6387 41940 6421
rect 41974 6387 41986 6421
rect 41928 6353 41986 6387
rect 41928 6319 41940 6353
rect 41974 6319 41986 6353
rect 41928 6288 41986 6319
<< mvpdiff >>
rect -6460 17183 -6402 17224
rect -6460 17149 -6448 17183
rect -6414 17149 -6402 17183
rect -6460 17115 -6402 17149
rect -6460 17081 -6448 17115
rect -6414 17081 -6402 17115
rect -6460 17047 -6402 17081
rect -6460 17013 -6448 17047
rect -6414 17013 -6402 17047
rect -6460 16979 -6402 17013
rect -6460 16945 -6448 16979
rect -6414 16945 -6402 16979
rect -6460 16911 -6402 16945
rect -6460 16877 -6448 16911
rect -6414 16877 -6402 16911
rect -6460 16843 -6402 16877
rect -6460 16809 -6448 16843
rect -6414 16809 -6402 16843
rect -6460 16775 -6402 16809
rect -6460 16741 -6448 16775
rect -6414 16741 -6402 16775
rect -6460 16707 -6402 16741
rect -6460 16673 -6448 16707
rect -6414 16673 -6402 16707
rect -6460 16639 -6402 16673
rect -6460 16605 -6448 16639
rect -6414 16605 -6402 16639
rect -6460 16571 -6402 16605
rect -6460 16537 -6448 16571
rect -6414 16537 -6402 16571
rect -6460 16503 -6402 16537
rect -6460 16469 -6448 16503
rect -6414 16469 -6402 16503
rect -6460 16435 -6402 16469
rect -6460 16401 -6448 16435
rect -6414 16401 -6402 16435
rect -6460 16367 -6402 16401
rect -6460 16333 -6448 16367
rect -6414 16333 -6402 16367
rect -6460 16299 -6402 16333
rect -6460 16265 -6448 16299
rect -6414 16265 -6402 16299
rect -6460 16224 -6402 16265
rect -6202 17183 -6144 17224
rect -6202 17149 -6190 17183
rect -6156 17149 -6144 17183
rect -6202 17115 -6144 17149
rect -6202 17081 -6190 17115
rect -6156 17081 -6144 17115
rect -6202 17047 -6144 17081
rect -6202 17013 -6190 17047
rect -6156 17013 -6144 17047
rect -6202 16979 -6144 17013
rect -6202 16945 -6190 16979
rect -6156 16945 -6144 16979
rect -6202 16911 -6144 16945
rect -6202 16877 -6190 16911
rect -6156 16877 -6144 16911
rect -6202 16843 -6144 16877
rect -6202 16809 -6190 16843
rect -6156 16809 -6144 16843
rect -6202 16775 -6144 16809
rect -6202 16741 -6190 16775
rect -6156 16741 -6144 16775
rect -6202 16707 -6144 16741
rect -6202 16673 -6190 16707
rect -6156 16673 -6144 16707
rect -6202 16639 -6144 16673
rect -6202 16605 -6190 16639
rect -6156 16605 -6144 16639
rect -6202 16571 -6144 16605
rect -6202 16537 -6190 16571
rect -6156 16537 -6144 16571
rect -6202 16503 -6144 16537
rect -6202 16469 -6190 16503
rect -6156 16469 -6144 16503
rect -6202 16435 -6144 16469
rect -6202 16401 -6190 16435
rect -6156 16401 -6144 16435
rect -6202 16367 -6144 16401
rect -6202 16333 -6190 16367
rect -6156 16333 -6144 16367
rect -6202 16299 -6144 16333
rect -6202 16265 -6190 16299
rect -6156 16265 -6144 16299
rect -6202 16224 -6144 16265
rect -5944 17183 -5886 17224
rect -5944 17149 -5932 17183
rect -5898 17149 -5886 17183
rect -5944 17115 -5886 17149
rect -5944 17081 -5932 17115
rect -5898 17081 -5886 17115
rect -5944 17047 -5886 17081
rect -5944 17013 -5932 17047
rect -5898 17013 -5886 17047
rect -5944 16979 -5886 17013
rect -5944 16945 -5932 16979
rect -5898 16945 -5886 16979
rect -5944 16911 -5886 16945
rect -5944 16877 -5932 16911
rect -5898 16877 -5886 16911
rect -5944 16843 -5886 16877
rect -5944 16809 -5932 16843
rect -5898 16809 -5886 16843
rect -5944 16775 -5886 16809
rect -5944 16741 -5932 16775
rect -5898 16741 -5886 16775
rect -5944 16707 -5886 16741
rect -5944 16673 -5932 16707
rect -5898 16673 -5886 16707
rect -5944 16639 -5886 16673
rect -5944 16605 -5932 16639
rect -5898 16605 -5886 16639
rect -5944 16571 -5886 16605
rect -5944 16537 -5932 16571
rect -5898 16537 -5886 16571
rect -5944 16503 -5886 16537
rect -5944 16469 -5932 16503
rect -5898 16469 -5886 16503
rect -5944 16435 -5886 16469
rect -5944 16401 -5932 16435
rect -5898 16401 -5886 16435
rect -5944 16367 -5886 16401
rect -5944 16333 -5932 16367
rect -5898 16333 -5886 16367
rect -5944 16299 -5886 16333
rect -5944 16265 -5932 16299
rect -5898 16265 -5886 16299
rect -5944 16224 -5886 16265
rect -2992 18062 -2934 18093
rect -2992 18028 -2980 18062
rect -2946 18028 -2934 18062
rect -2992 17994 -2934 18028
rect -2992 17960 -2980 17994
rect -2946 17960 -2934 17994
rect -2992 17926 -2934 17960
rect -2992 17892 -2980 17926
rect -2946 17892 -2934 17926
rect -2992 17858 -2934 17892
rect -2992 17824 -2980 17858
rect -2946 17824 -2934 17858
rect -2992 17790 -2934 17824
rect -2992 17756 -2980 17790
rect -2946 17756 -2934 17790
rect -2992 17722 -2934 17756
rect -2992 17688 -2980 17722
rect -2946 17688 -2934 17722
rect -2992 17654 -2934 17688
rect -2992 17620 -2980 17654
rect -2946 17620 -2934 17654
rect -2992 17586 -2934 17620
rect -2992 17552 -2980 17586
rect -2946 17552 -2934 17586
rect -2992 17518 -2934 17552
rect -2992 17484 -2980 17518
rect -2946 17484 -2934 17518
rect -2992 17450 -2934 17484
rect -2992 17416 -2980 17450
rect -2946 17416 -2934 17450
rect -2992 17382 -2934 17416
rect -2992 17348 -2980 17382
rect -2946 17348 -2934 17382
rect -2992 17314 -2934 17348
rect -2992 17280 -2980 17314
rect -2946 17280 -2934 17314
rect -2992 17246 -2934 17280
rect -2992 17212 -2980 17246
rect -2946 17212 -2934 17246
rect -2992 17178 -2934 17212
rect -2992 17144 -2980 17178
rect -2946 17144 -2934 17178
rect -2992 17110 -2934 17144
rect -2992 17076 -2980 17110
rect -2946 17076 -2934 17110
rect -2992 17042 -2934 17076
rect -2992 17008 -2980 17042
rect -2946 17008 -2934 17042
rect -2992 16974 -2934 17008
rect -2992 16940 -2980 16974
rect -2946 16940 -2934 16974
rect -2992 16906 -2934 16940
rect -2992 16872 -2980 16906
rect -2946 16872 -2934 16906
rect -2992 16838 -2934 16872
rect -2992 16804 -2980 16838
rect -2946 16804 -2934 16838
rect -2992 16770 -2934 16804
rect -2992 16736 -2980 16770
rect -2946 16736 -2934 16770
rect -2992 16702 -2934 16736
rect -2992 16668 -2980 16702
rect -2946 16668 -2934 16702
rect -2992 16634 -2934 16668
rect -2992 16600 -2980 16634
rect -2946 16600 -2934 16634
rect -2992 16566 -2934 16600
rect -2992 16532 -2980 16566
rect -2946 16532 -2934 16566
rect -2992 16498 -2934 16532
rect -2992 16464 -2980 16498
rect -2946 16464 -2934 16498
rect -2992 16430 -2934 16464
rect -2992 16396 -2980 16430
rect -2946 16396 -2934 16430
rect -2992 16362 -2934 16396
rect -2992 16328 -2980 16362
rect -2946 16328 -2934 16362
rect -2992 16294 -2934 16328
rect -2992 16260 -2980 16294
rect -2946 16260 -2934 16294
rect -2992 16226 -2934 16260
rect -2992 16192 -2980 16226
rect -2946 16192 -2934 16226
rect -2992 16158 -2934 16192
rect -2992 16124 -2980 16158
rect -2946 16124 -2934 16158
rect -2992 16093 -2934 16124
rect -2734 18062 -2676 18093
rect -2734 18028 -2722 18062
rect -2688 18028 -2676 18062
rect -2734 17994 -2676 18028
rect -2734 17960 -2722 17994
rect -2688 17960 -2676 17994
rect -2734 17926 -2676 17960
rect -2734 17892 -2722 17926
rect -2688 17892 -2676 17926
rect -2734 17858 -2676 17892
rect -2734 17824 -2722 17858
rect -2688 17824 -2676 17858
rect -2734 17790 -2676 17824
rect -2734 17756 -2722 17790
rect -2688 17756 -2676 17790
rect -2734 17722 -2676 17756
rect -2734 17688 -2722 17722
rect -2688 17688 -2676 17722
rect -2734 17654 -2676 17688
rect -2734 17620 -2722 17654
rect -2688 17620 -2676 17654
rect -2734 17586 -2676 17620
rect -2734 17552 -2722 17586
rect -2688 17552 -2676 17586
rect -2734 17518 -2676 17552
rect -2734 17484 -2722 17518
rect -2688 17484 -2676 17518
rect -2734 17450 -2676 17484
rect -2734 17416 -2722 17450
rect -2688 17416 -2676 17450
rect -2734 17382 -2676 17416
rect -2734 17348 -2722 17382
rect -2688 17348 -2676 17382
rect -2734 17314 -2676 17348
rect -2734 17280 -2722 17314
rect -2688 17280 -2676 17314
rect -2734 17246 -2676 17280
rect -2734 17212 -2722 17246
rect -2688 17212 -2676 17246
rect -2734 17178 -2676 17212
rect -2734 17144 -2722 17178
rect -2688 17144 -2676 17178
rect -2734 17110 -2676 17144
rect -2734 17076 -2722 17110
rect -2688 17076 -2676 17110
rect -2734 17042 -2676 17076
rect -2734 17008 -2722 17042
rect -2688 17008 -2676 17042
rect -2734 16974 -2676 17008
rect -2734 16940 -2722 16974
rect -2688 16940 -2676 16974
rect -2734 16906 -2676 16940
rect -2734 16872 -2722 16906
rect -2688 16872 -2676 16906
rect -2734 16838 -2676 16872
rect -2734 16804 -2722 16838
rect -2688 16804 -2676 16838
rect -2734 16770 -2676 16804
rect -2734 16736 -2722 16770
rect -2688 16736 -2676 16770
rect -2734 16702 -2676 16736
rect -2734 16668 -2722 16702
rect -2688 16668 -2676 16702
rect -2734 16634 -2676 16668
rect -2734 16600 -2722 16634
rect -2688 16600 -2676 16634
rect -2734 16566 -2676 16600
rect -2734 16532 -2722 16566
rect -2688 16532 -2676 16566
rect -2734 16498 -2676 16532
rect -2734 16464 -2722 16498
rect -2688 16464 -2676 16498
rect -2734 16430 -2676 16464
rect -2734 16396 -2722 16430
rect -2688 16396 -2676 16430
rect -2734 16362 -2676 16396
rect -2734 16328 -2722 16362
rect -2688 16328 -2676 16362
rect -2734 16294 -2676 16328
rect -2734 16260 -2722 16294
rect -2688 16260 -2676 16294
rect -2734 16226 -2676 16260
rect -2734 16192 -2722 16226
rect -2688 16192 -2676 16226
rect -2734 16158 -2676 16192
rect -2734 16124 -2722 16158
rect -2688 16124 -2676 16158
rect -2734 16093 -2676 16124
rect -2476 18062 -2418 18093
rect -2476 18028 -2464 18062
rect -2430 18028 -2418 18062
rect -2476 17994 -2418 18028
rect -2476 17960 -2464 17994
rect -2430 17960 -2418 17994
rect -2476 17926 -2418 17960
rect -2476 17892 -2464 17926
rect -2430 17892 -2418 17926
rect -2476 17858 -2418 17892
rect -2476 17824 -2464 17858
rect -2430 17824 -2418 17858
rect -2476 17790 -2418 17824
rect -2476 17756 -2464 17790
rect -2430 17756 -2418 17790
rect -2476 17722 -2418 17756
rect -2476 17688 -2464 17722
rect -2430 17688 -2418 17722
rect -2476 17654 -2418 17688
rect -2476 17620 -2464 17654
rect -2430 17620 -2418 17654
rect -2476 17586 -2418 17620
rect -2476 17552 -2464 17586
rect -2430 17552 -2418 17586
rect -2476 17518 -2418 17552
rect -2476 17484 -2464 17518
rect -2430 17484 -2418 17518
rect -2476 17450 -2418 17484
rect -2476 17416 -2464 17450
rect -2430 17416 -2418 17450
rect -2476 17382 -2418 17416
rect -2476 17348 -2464 17382
rect -2430 17348 -2418 17382
rect -2476 17314 -2418 17348
rect -2476 17280 -2464 17314
rect -2430 17280 -2418 17314
rect -2476 17246 -2418 17280
rect -2476 17212 -2464 17246
rect -2430 17212 -2418 17246
rect -2476 17178 -2418 17212
rect -2476 17144 -2464 17178
rect -2430 17144 -2418 17178
rect -2476 17110 -2418 17144
rect -2476 17076 -2464 17110
rect -2430 17076 -2418 17110
rect -2476 17042 -2418 17076
rect -2476 17008 -2464 17042
rect -2430 17008 -2418 17042
rect -2476 16974 -2418 17008
rect -2476 16940 -2464 16974
rect -2430 16940 -2418 16974
rect -2476 16906 -2418 16940
rect -2476 16872 -2464 16906
rect -2430 16872 -2418 16906
rect -2476 16838 -2418 16872
rect -2476 16804 -2464 16838
rect -2430 16804 -2418 16838
rect -2476 16770 -2418 16804
rect -2476 16736 -2464 16770
rect -2430 16736 -2418 16770
rect -2476 16702 -2418 16736
rect -2476 16668 -2464 16702
rect -2430 16668 -2418 16702
rect -2476 16634 -2418 16668
rect -2476 16600 -2464 16634
rect -2430 16600 -2418 16634
rect -2476 16566 -2418 16600
rect -2476 16532 -2464 16566
rect -2430 16532 -2418 16566
rect -2476 16498 -2418 16532
rect -2476 16464 -2464 16498
rect -2430 16464 -2418 16498
rect -2476 16430 -2418 16464
rect -2476 16396 -2464 16430
rect -2430 16396 -2418 16430
rect -2476 16362 -2418 16396
rect -2476 16328 -2464 16362
rect -2430 16328 -2418 16362
rect -2476 16294 -2418 16328
rect -2476 16260 -2464 16294
rect -2430 16260 -2418 16294
rect -2476 16226 -2418 16260
rect -2476 16192 -2464 16226
rect -2430 16192 -2418 16226
rect -2476 16158 -2418 16192
rect -2476 16124 -2464 16158
rect -2430 16124 -2418 16158
rect -2476 16093 -2418 16124
rect -2218 18062 -2160 18093
rect -2218 18028 -2206 18062
rect -2172 18028 -2160 18062
rect -2218 17994 -2160 18028
rect -2218 17960 -2206 17994
rect -2172 17960 -2160 17994
rect -2218 17926 -2160 17960
rect -2218 17892 -2206 17926
rect -2172 17892 -2160 17926
rect -2218 17858 -2160 17892
rect -2218 17824 -2206 17858
rect -2172 17824 -2160 17858
rect -2218 17790 -2160 17824
rect -2218 17756 -2206 17790
rect -2172 17756 -2160 17790
rect -2218 17722 -2160 17756
rect -2218 17688 -2206 17722
rect -2172 17688 -2160 17722
rect -2218 17654 -2160 17688
rect -2218 17620 -2206 17654
rect -2172 17620 -2160 17654
rect -2218 17586 -2160 17620
rect -2218 17552 -2206 17586
rect -2172 17552 -2160 17586
rect -2218 17518 -2160 17552
rect -2218 17484 -2206 17518
rect -2172 17484 -2160 17518
rect -2218 17450 -2160 17484
rect -2218 17416 -2206 17450
rect -2172 17416 -2160 17450
rect -2218 17382 -2160 17416
rect -2218 17348 -2206 17382
rect -2172 17348 -2160 17382
rect -2218 17314 -2160 17348
rect -2218 17280 -2206 17314
rect -2172 17280 -2160 17314
rect -2218 17246 -2160 17280
rect -2218 17212 -2206 17246
rect -2172 17212 -2160 17246
rect -2218 17178 -2160 17212
rect -2218 17144 -2206 17178
rect -2172 17144 -2160 17178
rect -2218 17110 -2160 17144
rect -2218 17076 -2206 17110
rect -2172 17076 -2160 17110
rect -2218 17042 -2160 17076
rect -2218 17008 -2206 17042
rect -2172 17008 -2160 17042
rect -2218 16974 -2160 17008
rect -2218 16940 -2206 16974
rect -2172 16940 -2160 16974
rect -2218 16906 -2160 16940
rect -2218 16872 -2206 16906
rect -2172 16872 -2160 16906
rect -2218 16838 -2160 16872
rect -2218 16804 -2206 16838
rect -2172 16804 -2160 16838
rect -2218 16770 -2160 16804
rect -2218 16736 -2206 16770
rect -2172 16736 -2160 16770
rect -2218 16702 -2160 16736
rect -2218 16668 -2206 16702
rect -2172 16668 -2160 16702
rect -2218 16634 -2160 16668
rect -2218 16600 -2206 16634
rect -2172 16600 -2160 16634
rect -2218 16566 -2160 16600
rect -2218 16532 -2206 16566
rect -2172 16532 -2160 16566
rect -2218 16498 -2160 16532
rect -2218 16464 -2206 16498
rect -2172 16464 -2160 16498
rect -2218 16430 -2160 16464
rect -2218 16396 -2206 16430
rect -2172 16396 -2160 16430
rect -2218 16362 -2160 16396
rect -2218 16328 -2206 16362
rect -2172 16328 -2160 16362
rect -2218 16294 -2160 16328
rect -2218 16260 -2206 16294
rect -2172 16260 -2160 16294
rect -2218 16226 -2160 16260
rect -2218 16192 -2206 16226
rect -2172 16192 -2160 16226
rect -2218 16158 -2160 16192
rect -2218 16124 -2206 16158
rect -2172 16124 -2160 16158
rect -2218 16093 -2160 16124
rect -1960 18062 -1902 18093
rect -1960 18028 -1948 18062
rect -1914 18028 -1902 18062
rect -1960 17994 -1902 18028
rect -1960 17960 -1948 17994
rect -1914 17960 -1902 17994
rect -1960 17926 -1902 17960
rect -1960 17892 -1948 17926
rect -1914 17892 -1902 17926
rect -1960 17858 -1902 17892
rect -1960 17824 -1948 17858
rect -1914 17824 -1902 17858
rect -1960 17790 -1902 17824
rect -1960 17756 -1948 17790
rect -1914 17756 -1902 17790
rect -1960 17722 -1902 17756
rect -1960 17688 -1948 17722
rect -1914 17688 -1902 17722
rect -1960 17654 -1902 17688
rect -1960 17620 -1948 17654
rect -1914 17620 -1902 17654
rect -1960 17586 -1902 17620
rect -1960 17552 -1948 17586
rect -1914 17552 -1902 17586
rect -1960 17518 -1902 17552
rect -1960 17484 -1948 17518
rect -1914 17484 -1902 17518
rect -1960 17450 -1902 17484
rect -1960 17416 -1948 17450
rect -1914 17416 -1902 17450
rect -1960 17382 -1902 17416
rect -1960 17348 -1948 17382
rect -1914 17348 -1902 17382
rect -1960 17314 -1902 17348
rect -1960 17280 -1948 17314
rect -1914 17280 -1902 17314
rect -1960 17246 -1902 17280
rect -1960 17212 -1948 17246
rect -1914 17212 -1902 17246
rect -1960 17178 -1902 17212
rect -1960 17144 -1948 17178
rect -1914 17144 -1902 17178
rect -1960 17110 -1902 17144
rect -1960 17076 -1948 17110
rect -1914 17076 -1902 17110
rect -1960 17042 -1902 17076
rect -1960 17008 -1948 17042
rect -1914 17008 -1902 17042
rect -1960 16974 -1902 17008
rect -1960 16940 -1948 16974
rect -1914 16940 -1902 16974
rect -1960 16906 -1902 16940
rect -1960 16872 -1948 16906
rect -1914 16872 -1902 16906
rect -1960 16838 -1902 16872
rect -1960 16804 -1948 16838
rect -1914 16804 -1902 16838
rect -1960 16770 -1902 16804
rect -1960 16736 -1948 16770
rect -1914 16736 -1902 16770
rect -1960 16702 -1902 16736
rect -1960 16668 -1948 16702
rect -1914 16668 -1902 16702
rect -1960 16634 -1902 16668
rect -1960 16600 -1948 16634
rect -1914 16600 -1902 16634
rect -1960 16566 -1902 16600
rect -1960 16532 -1948 16566
rect -1914 16532 -1902 16566
rect -1960 16498 -1902 16532
rect -1960 16464 -1948 16498
rect -1914 16464 -1902 16498
rect -1960 16430 -1902 16464
rect -1960 16396 -1948 16430
rect -1914 16396 -1902 16430
rect -1960 16362 -1902 16396
rect -1960 16328 -1948 16362
rect -1914 16328 -1902 16362
rect -1960 16294 -1902 16328
rect -1960 16260 -1948 16294
rect -1914 16260 -1902 16294
rect -1960 16226 -1902 16260
rect -1960 16192 -1948 16226
rect -1914 16192 -1902 16226
rect -1960 16158 -1902 16192
rect -1960 16124 -1948 16158
rect -1914 16124 -1902 16158
rect -1960 16093 -1902 16124
rect -1702 18062 -1644 18093
rect -1702 18028 -1690 18062
rect -1656 18028 -1644 18062
rect -1702 17994 -1644 18028
rect -1702 17960 -1690 17994
rect -1656 17960 -1644 17994
rect -1702 17926 -1644 17960
rect -1702 17892 -1690 17926
rect -1656 17892 -1644 17926
rect -1702 17858 -1644 17892
rect -1702 17824 -1690 17858
rect -1656 17824 -1644 17858
rect -1702 17790 -1644 17824
rect -1702 17756 -1690 17790
rect -1656 17756 -1644 17790
rect -1702 17722 -1644 17756
rect -1702 17688 -1690 17722
rect -1656 17688 -1644 17722
rect -1702 17654 -1644 17688
rect -1702 17620 -1690 17654
rect -1656 17620 -1644 17654
rect -1702 17586 -1644 17620
rect -1702 17552 -1690 17586
rect -1656 17552 -1644 17586
rect -1702 17518 -1644 17552
rect -1702 17484 -1690 17518
rect -1656 17484 -1644 17518
rect -1702 17450 -1644 17484
rect -1702 17416 -1690 17450
rect -1656 17416 -1644 17450
rect -1702 17382 -1644 17416
rect -1702 17348 -1690 17382
rect -1656 17348 -1644 17382
rect -1702 17314 -1644 17348
rect -1702 17280 -1690 17314
rect -1656 17280 -1644 17314
rect -1702 17246 -1644 17280
rect -1702 17212 -1690 17246
rect -1656 17212 -1644 17246
rect -1702 17178 -1644 17212
rect -1702 17144 -1690 17178
rect -1656 17144 -1644 17178
rect -1702 17110 -1644 17144
rect -1702 17076 -1690 17110
rect -1656 17076 -1644 17110
rect -1702 17042 -1644 17076
rect -1702 17008 -1690 17042
rect -1656 17008 -1644 17042
rect -1702 16974 -1644 17008
rect -1702 16940 -1690 16974
rect -1656 16940 -1644 16974
rect -1702 16906 -1644 16940
rect -1702 16872 -1690 16906
rect -1656 16872 -1644 16906
rect -1702 16838 -1644 16872
rect -1702 16804 -1690 16838
rect -1656 16804 -1644 16838
rect -1702 16770 -1644 16804
rect -1702 16736 -1690 16770
rect -1656 16736 -1644 16770
rect -1702 16702 -1644 16736
rect -1702 16668 -1690 16702
rect -1656 16668 -1644 16702
rect -1702 16634 -1644 16668
rect -1702 16600 -1690 16634
rect -1656 16600 -1644 16634
rect -1702 16566 -1644 16600
rect -1702 16532 -1690 16566
rect -1656 16532 -1644 16566
rect -1702 16498 -1644 16532
rect -1702 16464 -1690 16498
rect -1656 16464 -1644 16498
rect -1702 16430 -1644 16464
rect -1702 16396 -1690 16430
rect -1656 16396 -1644 16430
rect -1702 16362 -1644 16396
rect -1702 16328 -1690 16362
rect -1656 16328 -1644 16362
rect -1702 16294 -1644 16328
rect -1702 16260 -1690 16294
rect -1656 16260 -1644 16294
rect -1702 16226 -1644 16260
rect -1702 16192 -1690 16226
rect -1656 16192 -1644 16226
rect -1702 16158 -1644 16192
rect -1702 16124 -1690 16158
rect -1656 16124 -1644 16158
rect -1702 16093 -1644 16124
rect -1444 18062 -1386 18093
rect -1444 18028 -1432 18062
rect -1398 18028 -1386 18062
rect -1444 17994 -1386 18028
rect -1444 17960 -1432 17994
rect -1398 17960 -1386 17994
rect -1444 17926 -1386 17960
rect -1444 17892 -1432 17926
rect -1398 17892 -1386 17926
rect -1444 17858 -1386 17892
rect -1444 17824 -1432 17858
rect -1398 17824 -1386 17858
rect -1444 17790 -1386 17824
rect -1444 17756 -1432 17790
rect -1398 17756 -1386 17790
rect -1444 17722 -1386 17756
rect -1444 17688 -1432 17722
rect -1398 17688 -1386 17722
rect -1444 17654 -1386 17688
rect -1444 17620 -1432 17654
rect -1398 17620 -1386 17654
rect -1444 17586 -1386 17620
rect -1444 17552 -1432 17586
rect -1398 17552 -1386 17586
rect -1444 17518 -1386 17552
rect -1444 17484 -1432 17518
rect -1398 17484 -1386 17518
rect -1444 17450 -1386 17484
rect -1444 17416 -1432 17450
rect -1398 17416 -1386 17450
rect -1444 17382 -1386 17416
rect -1444 17348 -1432 17382
rect -1398 17348 -1386 17382
rect -1444 17314 -1386 17348
rect -1444 17280 -1432 17314
rect -1398 17280 -1386 17314
rect -1444 17246 -1386 17280
rect -1444 17212 -1432 17246
rect -1398 17212 -1386 17246
rect -1444 17178 -1386 17212
rect -1444 17144 -1432 17178
rect -1398 17144 -1386 17178
rect -1444 17110 -1386 17144
rect -1444 17076 -1432 17110
rect -1398 17076 -1386 17110
rect -1444 17042 -1386 17076
rect -1444 17008 -1432 17042
rect -1398 17008 -1386 17042
rect -1444 16974 -1386 17008
rect -1444 16940 -1432 16974
rect -1398 16940 -1386 16974
rect -1444 16906 -1386 16940
rect -1444 16872 -1432 16906
rect -1398 16872 -1386 16906
rect -1444 16838 -1386 16872
rect -1444 16804 -1432 16838
rect -1398 16804 -1386 16838
rect -1444 16770 -1386 16804
rect -1444 16736 -1432 16770
rect -1398 16736 -1386 16770
rect -1444 16702 -1386 16736
rect -1444 16668 -1432 16702
rect -1398 16668 -1386 16702
rect -1444 16634 -1386 16668
rect -1444 16600 -1432 16634
rect -1398 16600 -1386 16634
rect -1444 16566 -1386 16600
rect -1444 16532 -1432 16566
rect -1398 16532 -1386 16566
rect -1444 16498 -1386 16532
rect -1444 16464 -1432 16498
rect -1398 16464 -1386 16498
rect -1444 16430 -1386 16464
rect -1444 16396 -1432 16430
rect -1398 16396 -1386 16430
rect -1444 16362 -1386 16396
rect -1444 16328 -1432 16362
rect -1398 16328 -1386 16362
rect -1444 16294 -1386 16328
rect -1444 16260 -1432 16294
rect -1398 16260 -1386 16294
rect -1444 16226 -1386 16260
rect -1444 16192 -1432 16226
rect -1398 16192 -1386 16226
rect -1444 16158 -1386 16192
rect -1444 16124 -1432 16158
rect -1398 16124 -1386 16158
rect -1444 16093 -1386 16124
rect -1186 18062 -1128 18093
rect -1186 18028 -1174 18062
rect -1140 18028 -1128 18062
rect -1186 17994 -1128 18028
rect -1186 17960 -1174 17994
rect -1140 17960 -1128 17994
rect -1186 17926 -1128 17960
rect -1186 17892 -1174 17926
rect -1140 17892 -1128 17926
rect -1186 17858 -1128 17892
rect -1186 17824 -1174 17858
rect -1140 17824 -1128 17858
rect -1186 17790 -1128 17824
rect -1186 17756 -1174 17790
rect -1140 17756 -1128 17790
rect -1186 17722 -1128 17756
rect -1186 17688 -1174 17722
rect -1140 17688 -1128 17722
rect -1186 17654 -1128 17688
rect -1186 17620 -1174 17654
rect -1140 17620 -1128 17654
rect -1186 17586 -1128 17620
rect -1186 17552 -1174 17586
rect -1140 17552 -1128 17586
rect -1186 17518 -1128 17552
rect -1186 17484 -1174 17518
rect -1140 17484 -1128 17518
rect -1186 17450 -1128 17484
rect -1186 17416 -1174 17450
rect -1140 17416 -1128 17450
rect -1186 17382 -1128 17416
rect -1186 17348 -1174 17382
rect -1140 17348 -1128 17382
rect -1186 17314 -1128 17348
rect -1186 17280 -1174 17314
rect -1140 17280 -1128 17314
rect -1186 17246 -1128 17280
rect -1186 17212 -1174 17246
rect -1140 17212 -1128 17246
rect -1186 17178 -1128 17212
rect -1186 17144 -1174 17178
rect -1140 17144 -1128 17178
rect -1186 17110 -1128 17144
rect -1186 17076 -1174 17110
rect -1140 17076 -1128 17110
rect -1186 17042 -1128 17076
rect -1186 17008 -1174 17042
rect -1140 17008 -1128 17042
rect -1186 16974 -1128 17008
rect -1186 16940 -1174 16974
rect -1140 16940 -1128 16974
rect -1186 16906 -1128 16940
rect -1186 16872 -1174 16906
rect -1140 16872 -1128 16906
rect -1186 16838 -1128 16872
rect -1186 16804 -1174 16838
rect -1140 16804 -1128 16838
rect -1186 16770 -1128 16804
rect -1186 16736 -1174 16770
rect -1140 16736 -1128 16770
rect -1186 16702 -1128 16736
rect -1186 16668 -1174 16702
rect -1140 16668 -1128 16702
rect -1186 16634 -1128 16668
rect -1186 16600 -1174 16634
rect -1140 16600 -1128 16634
rect -1186 16566 -1128 16600
rect -1186 16532 -1174 16566
rect -1140 16532 -1128 16566
rect -1186 16498 -1128 16532
rect -1186 16464 -1174 16498
rect -1140 16464 -1128 16498
rect -1186 16430 -1128 16464
rect -1186 16396 -1174 16430
rect -1140 16396 -1128 16430
rect -1186 16362 -1128 16396
rect -1186 16328 -1174 16362
rect -1140 16328 -1128 16362
rect -1186 16294 -1128 16328
rect -1186 16260 -1174 16294
rect -1140 16260 -1128 16294
rect -1186 16226 -1128 16260
rect -1186 16192 -1174 16226
rect -1140 16192 -1128 16226
rect -1186 16158 -1128 16192
rect -1186 16124 -1174 16158
rect -1140 16124 -1128 16158
rect -1186 16093 -1128 16124
rect -928 18062 -870 18093
rect -928 18028 -916 18062
rect -882 18028 -870 18062
rect -928 17994 -870 18028
rect -928 17960 -916 17994
rect -882 17960 -870 17994
rect -928 17926 -870 17960
rect -928 17892 -916 17926
rect -882 17892 -870 17926
rect -928 17858 -870 17892
rect -928 17824 -916 17858
rect -882 17824 -870 17858
rect -928 17790 -870 17824
rect -928 17756 -916 17790
rect -882 17756 -870 17790
rect -928 17722 -870 17756
rect -928 17688 -916 17722
rect -882 17688 -870 17722
rect -928 17654 -870 17688
rect -928 17620 -916 17654
rect -882 17620 -870 17654
rect -928 17586 -870 17620
rect -928 17552 -916 17586
rect -882 17552 -870 17586
rect -928 17518 -870 17552
rect -928 17484 -916 17518
rect -882 17484 -870 17518
rect -928 17450 -870 17484
rect -928 17416 -916 17450
rect -882 17416 -870 17450
rect -928 17382 -870 17416
rect -928 17348 -916 17382
rect -882 17348 -870 17382
rect -928 17314 -870 17348
rect -928 17280 -916 17314
rect -882 17280 -870 17314
rect -928 17246 -870 17280
rect -928 17212 -916 17246
rect -882 17212 -870 17246
rect -928 17178 -870 17212
rect -928 17144 -916 17178
rect -882 17144 -870 17178
rect -928 17110 -870 17144
rect -928 17076 -916 17110
rect -882 17076 -870 17110
rect -928 17042 -870 17076
rect -928 17008 -916 17042
rect -882 17008 -870 17042
rect -928 16974 -870 17008
rect -928 16940 -916 16974
rect -882 16940 -870 16974
rect -928 16906 -870 16940
rect -928 16872 -916 16906
rect -882 16872 -870 16906
rect -928 16838 -870 16872
rect -928 16804 -916 16838
rect -882 16804 -870 16838
rect -928 16770 -870 16804
rect -928 16736 -916 16770
rect -882 16736 -870 16770
rect -928 16702 -870 16736
rect -928 16668 -916 16702
rect -882 16668 -870 16702
rect -928 16634 -870 16668
rect -928 16600 -916 16634
rect -882 16600 -870 16634
rect -928 16566 -870 16600
rect -928 16532 -916 16566
rect -882 16532 -870 16566
rect -928 16498 -870 16532
rect -928 16464 -916 16498
rect -882 16464 -870 16498
rect -928 16430 -870 16464
rect -928 16396 -916 16430
rect -882 16396 -870 16430
rect -928 16362 -870 16396
rect -928 16328 -916 16362
rect -882 16328 -870 16362
rect -928 16294 -870 16328
rect -928 16260 -916 16294
rect -882 16260 -870 16294
rect -928 16226 -870 16260
rect -928 16192 -916 16226
rect -882 16192 -870 16226
rect -928 16158 -870 16192
rect -928 16124 -916 16158
rect -882 16124 -870 16158
rect -928 16093 -870 16124
rect -670 18062 -612 18093
rect -670 18028 -658 18062
rect -624 18028 -612 18062
rect -670 17994 -612 18028
rect -670 17960 -658 17994
rect -624 17960 -612 17994
rect -670 17926 -612 17960
rect -670 17892 -658 17926
rect -624 17892 -612 17926
rect -670 17858 -612 17892
rect -670 17824 -658 17858
rect -624 17824 -612 17858
rect -670 17790 -612 17824
rect -670 17756 -658 17790
rect -624 17756 -612 17790
rect -670 17722 -612 17756
rect -670 17688 -658 17722
rect -624 17688 -612 17722
rect -670 17654 -612 17688
rect -670 17620 -658 17654
rect -624 17620 -612 17654
rect -670 17586 -612 17620
rect -670 17552 -658 17586
rect -624 17552 -612 17586
rect -670 17518 -612 17552
rect -670 17484 -658 17518
rect -624 17484 -612 17518
rect -670 17450 -612 17484
rect -670 17416 -658 17450
rect -624 17416 -612 17450
rect -670 17382 -612 17416
rect -670 17348 -658 17382
rect -624 17348 -612 17382
rect -670 17314 -612 17348
rect -670 17280 -658 17314
rect -624 17280 -612 17314
rect -670 17246 -612 17280
rect -670 17212 -658 17246
rect -624 17212 -612 17246
rect -670 17178 -612 17212
rect -670 17144 -658 17178
rect -624 17144 -612 17178
rect -670 17110 -612 17144
rect -670 17076 -658 17110
rect -624 17076 -612 17110
rect -670 17042 -612 17076
rect -670 17008 -658 17042
rect -624 17008 -612 17042
rect -670 16974 -612 17008
rect -670 16940 -658 16974
rect -624 16940 -612 16974
rect -670 16906 -612 16940
rect -670 16872 -658 16906
rect -624 16872 -612 16906
rect -670 16838 -612 16872
rect -670 16804 -658 16838
rect -624 16804 -612 16838
rect -670 16770 -612 16804
rect -670 16736 -658 16770
rect -624 16736 -612 16770
rect -670 16702 -612 16736
rect -670 16668 -658 16702
rect -624 16668 -612 16702
rect -670 16634 -612 16668
rect -670 16600 -658 16634
rect -624 16600 -612 16634
rect -670 16566 -612 16600
rect -670 16532 -658 16566
rect -624 16532 -612 16566
rect -670 16498 -612 16532
rect -670 16464 -658 16498
rect -624 16464 -612 16498
rect -670 16430 -612 16464
rect -670 16396 -658 16430
rect -624 16396 -612 16430
rect -670 16362 -612 16396
rect -670 16328 -658 16362
rect -624 16328 -612 16362
rect -670 16294 -612 16328
rect -670 16260 -658 16294
rect -624 16260 -612 16294
rect -670 16226 -612 16260
rect -670 16192 -658 16226
rect -624 16192 -612 16226
rect -670 16158 -612 16192
rect -670 16124 -658 16158
rect -624 16124 -612 16158
rect -670 16093 -612 16124
rect -412 18062 -354 18093
rect -412 18028 -400 18062
rect -366 18028 -354 18062
rect -412 17994 -354 18028
rect -412 17960 -400 17994
rect -366 17960 -354 17994
rect -412 17926 -354 17960
rect -412 17892 -400 17926
rect -366 17892 -354 17926
rect -412 17858 -354 17892
rect -412 17824 -400 17858
rect -366 17824 -354 17858
rect -412 17790 -354 17824
rect -412 17756 -400 17790
rect -366 17756 -354 17790
rect -412 17722 -354 17756
rect -412 17688 -400 17722
rect -366 17688 -354 17722
rect -412 17654 -354 17688
rect -412 17620 -400 17654
rect -366 17620 -354 17654
rect -412 17586 -354 17620
rect -412 17552 -400 17586
rect -366 17552 -354 17586
rect -412 17518 -354 17552
rect -412 17484 -400 17518
rect -366 17484 -354 17518
rect -412 17450 -354 17484
rect -412 17416 -400 17450
rect -366 17416 -354 17450
rect -412 17382 -354 17416
rect -412 17348 -400 17382
rect -366 17348 -354 17382
rect -412 17314 -354 17348
rect -412 17280 -400 17314
rect -366 17280 -354 17314
rect -412 17246 -354 17280
rect -412 17212 -400 17246
rect -366 17212 -354 17246
rect -412 17178 -354 17212
rect -412 17144 -400 17178
rect -366 17144 -354 17178
rect -412 17110 -354 17144
rect -412 17076 -400 17110
rect -366 17076 -354 17110
rect -412 17042 -354 17076
rect -412 17008 -400 17042
rect -366 17008 -354 17042
rect -412 16974 -354 17008
rect -412 16940 -400 16974
rect -366 16940 -354 16974
rect -412 16906 -354 16940
rect -412 16872 -400 16906
rect -366 16872 -354 16906
rect -412 16838 -354 16872
rect -412 16804 -400 16838
rect -366 16804 -354 16838
rect -412 16770 -354 16804
rect -412 16736 -400 16770
rect -366 16736 -354 16770
rect -412 16702 -354 16736
rect -412 16668 -400 16702
rect -366 16668 -354 16702
rect -412 16634 -354 16668
rect -412 16600 -400 16634
rect -366 16600 -354 16634
rect -412 16566 -354 16600
rect -412 16532 -400 16566
rect -366 16532 -354 16566
rect -412 16498 -354 16532
rect -412 16464 -400 16498
rect -366 16464 -354 16498
rect -412 16430 -354 16464
rect -412 16396 -400 16430
rect -366 16396 -354 16430
rect -412 16362 -354 16396
rect -412 16328 -400 16362
rect -366 16328 -354 16362
rect -412 16294 -354 16328
rect -412 16260 -400 16294
rect -366 16260 -354 16294
rect -412 16226 -354 16260
rect -412 16192 -400 16226
rect -366 16192 -354 16226
rect -412 16158 -354 16192
rect -412 16124 -400 16158
rect -366 16124 -354 16158
rect -412 16093 -354 16124
rect 23164 18706 23222 18747
rect 23164 18672 23176 18706
rect 23210 18672 23222 18706
rect 23164 18638 23222 18672
rect 23164 18604 23176 18638
rect 23210 18604 23222 18638
rect 23164 18570 23222 18604
rect 23164 18536 23176 18570
rect 23210 18536 23222 18570
rect 23164 18502 23222 18536
rect 23164 18468 23176 18502
rect 23210 18468 23222 18502
rect 23164 18434 23222 18468
rect 23164 18400 23176 18434
rect 23210 18400 23222 18434
rect 23164 18366 23222 18400
rect 23164 18332 23176 18366
rect 23210 18332 23222 18366
rect 23164 18298 23222 18332
rect 23164 18264 23176 18298
rect 23210 18264 23222 18298
rect 23164 18230 23222 18264
rect 23164 18196 23176 18230
rect 23210 18196 23222 18230
rect 23164 18162 23222 18196
rect 23164 18128 23176 18162
rect 23210 18128 23222 18162
rect 23164 18094 23222 18128
rect 23164 18060 23176 18094
rect 23210 18060 23222 18094
rect 23164 18026 23222 18060
rect 23164 17992 23176 18026
rect 23210 17992 23222 18026
rect 23164 17958 23222 17992
rect 23164 17924 23176 17958
rect 23210 17924 23222 17958
rect 23164 17890 23222 17924
rect 23164 17856 23176 17890
rect 23210 17856 23222 17890
rect 23164 17822 23222 17856
rect 23164 17788 23176 17822
rect 23210 17788 23222 17822
rect 23164 17747 23222 17788
rect 24222 18706 24280 18747
rect 24222 18672 24234 18706
rect 24268 18672 24280 18706
rect 24222 18638 24280 18672
rect 24222 18604 24234 18638
rect 24268 18604 24280 18638
rect 24222 18570 24280 18604
rect 24222 18536 24234 18570
rect 24268 18536 24280 18570
rect 24222 18502 24280 18536
rect 24222 18468 24234 18502
rect 24268 18468 24280 18502
rect 24222 18434 24280 18468
rect 24222 18400 24234 18434
rect 24268 18400 24280 18434
rect 24222 18366 24280 18400
rect 24222 18332 24234 18366
rect 24268 18332 24280 18366
rect 24222 18298 24280 18332
rect 24222 18264 24234 18298
rect 24268 18264 24280 18298
rect 24222 18230 24280 18264
rect 24222 18196 24234 18230
rect 24268 18196 24280 18230
rect 24222 18162 24280 18196
rect 24222 18128 24234 18162
rect 24268 18128 24280 18162
rect 24222 18094 24280 18128
rect 24222 18060 24234 18094
rect 24268 18060 24280 18094
rect 24222 18026 24280 18060
rect 24222 17992 24234 18026
rect 24268 17992 24280 18026
rect 24222 17958 24280 17992
rect 24222 17924 24234 17958
rect 24268 17924 24280 17958
rect 24222 17890 24280 17924
rect 24222 17856 24234 17890
rect 24268 17856 24280 17890
rect 24222 17822 24280 17856
rect 24222 17788 24234 17822
rect 24268 17788 24280 17822
rect 24222 17747 24280 17788
rect 24680 18712 24738 18747
rect 24680 18678 24692 18712
rect 24726 18678 24738 18712
rect 24680 18644 24738 18678
rect 24680 18610 24692 18644
rect 24726 18610 24738 18644
rect 24680 18576 24738 18610
rect 24680 18542 24692 18576
rect 24726 18542 24738 18576
rect 24680 18508 24738 18542
rect 24680 18474 24692 18508
rect 24726 18474 24738 18508
rect 24680 18440 24738 18474
rect 24680 18406 24692 18440
rect 24726 18406 24738 18440
rect 24680 18372 24738 18406
rect 24680 18338 24692 18372
rect 24726 18338 24738 18372
rect 24680 18304 24738 18338
rect 24680 18270 24692 18304
rect 24726 18270 24738 18304
rect 24680 18236 24738 18270
rect 24680 18202 24692 18236
rect 24726 18202 24738 18236
rect 24680 18168 24738 18202
rect 24680 18134 24692 18168
rect 24726 18134 24738 18168
rect 24680 18100 24738 18134
rect 24680 18066 24692 18100
rect 24726 18066 24738 18100
rect 24680 18032 24738 18066
rect 24680 17998 24692 18032
rect 24726 17998 24738 18032
rect 24680 17964 24738 17998
rect 24680 17930 24692 17964
rect 24726 17930 24738 17964
rect 24680 17896 24738 17930
rect 24680 17862 24692 17896
rect 24726 17862 24738 17896
rect 24680 17828 24738 17862
rect 24680 17794 24692 17828
rect 24726 17794 24738 17828
rect 24680 17760 24738 17794
rect 24680 17726 24692 17760
rect 24726 17726 24738 17760
rect 24680 17692 24738 17726
rect 24680 17658 24692 17692
rect 24726 17658 24738 17692
rect 24680 17624 24738 17658
rect 24680 17590 24692 17624
rect 24726 17590 24738 17624
rect 24680 17556 24738 17590
rect 24680 17522 24692 17556
rect 24726 17522 24738 17556
rect 24680 17488 24738 17522
rect 24680 17454 24692 17488
rect 24726 17454 24738 17488
rect 24680 17420 24738 17454
rect 24680 17386 24692 17420
rect 24726 17386 24738 17420
rect 24680 17352 24738 17386
rect 24680 17318 24692 17352
rect 24726 17318 24738 17352
rect 24680 17284 24738 17318
rect 24680 17250 24692 17284
rect 24726 17250 24738 17284
rect 24680 17216 24738 17250
rect 24680 17182 24692 17216
rect 24726 17182 24738 17216
rect 24680 17147 24738 17182
rect 25738 18712 25796 18747
rect 25738 18678 25750 18712
rect 25784 18678 25796 18712
rect 25738 18644 25796 18678
rect 25738 18610 25750 18644
rect 25784 18610 25796 18644
rect 25738 18576 25796 18610
rect 25738 18542 25750 18576
rect 25784 18542 25796 18576
rect 25738 18508 25796 18542
rect 25738 18474 25750 18508
rect 25784 18474 25796 18508
rect 25738 18440 25796 18474
rect 25738 18406 25750 18440
rect 25784 18406 25796 18440
rect 25738 18372 25796 18406
rect 25738 18338 25750 18372
rect 25784 18338 25796 18372
rect 25738 18304 25796 18338
rect 25738 18270 25750 18304
rect 25784 18270 25796 18304
rect 25738 18236 25796 18270
rect 25738 18202 25750 18236
rect 25784 18202 25796 18236
rect 25738 18168 25796 18202
rect 25738 18134 25750 18168
rect 25784 18134 25796 18168
rect 25738 18100 25796 18134
rect 25738 18066 25750 18100
rect 25784 18066 25796 18100
rect 25738 18032 25796 18066
rect 25738 17998 25750 18032
rect 25784 17998 25796 18032
rect 25738 17964 25796 17998
rect 25738 17930 25750 17964
rect 25784 17930 25796 17964
rect 25738 17896 25796 17930
rect 25738 17862 25750 17896
rect 25784 17862 25796 17896
rect 25738 17828 25796 17862
rect 25738 17794 25750 17828
rect 25784 17794 25796 17828
rect 25738 17760 25796 17794
rect 25738 17726 25750 17760
rect 25784 17726 25796 17760
rect 25738 17692 25796 17726
rect 25738 17658 25750 17692
rect 25784 17658 25796 17692
rect 25738 17624 25796 17658
rect 25738 17590 25750 17624
rect 25784 17590 25796 17624
rect 25738 17556 25796 17590
rect 25738 17522 25750 17556
rect 25784 17522 25796 17556
rect 25738 17488 25796 17522
rect 25738 17454 25750 17488
rect 25784 17454 25796 17488
rect 25738 17420 25796 17454
rect 25738 17386 25750 17420
rect 25784 17386 25796 17420
rect 25738 17352 25796 17386
rect 25738 17318 25750 17352
rect 25784 17318 25796 17352
rect 25738 17284 25796 17318
rect 25738 17250 25750 17284
rect 25784 17250 25796 17284
rect 25738 17216 25796 17250
rect 25738 17182 25750 17216
rect 25784 17182 25796 17216
rect 25738 17147 25796 17182
rect 26796 18712 26854 18747
rect 26796 18678 26808 18712
rect 26842 18678 26854 18712
rect 26796 18644 26854 18678
rect 26796 18610 26808 18644
rect 26842 18610 26854 18644
rect 26796 18576 26854 18610
rect 26796 18542 26808 18576
rect 26842 18542 26854 18576
rect 26796 18508 26854 18542
rect 26796 18474 26808 18508
rect 26842 18474 26854 18508
rect 26796 18440 26854 18474
rect 26796 18406 26808 18440
rect 26842 18406 26854 18440
rect 26796 18372 26854 18406
rect 26796 18338 26808 18372
rect 26842 18338 26854 18372
rect 26796 18304 26854 18338
rect 26796 18270 26808 18304
rect 26842 18270 26854 18304
rect 26796 18236 26854 18270
rect 26796 18202 26808 18236
rect 26842 18202 26854 18236
rect 26796 18168 26854 18202
rect 26796 18134 26808 18168
rect 26842 18134 26854 18168
rect 26796 18100 26854 18134
rect 26796 18066 26808 18100
rect 26842 18066 26854 18100
rect 26796 18032 26854 18066
rect 26796 17998 26808 18032
rect 26842 17998 26854 18032
rect 26796 17964 26854 17998
rect 26796 17930 26808 17964
rect 26842 17930 26854 17964
rect 26796 17896 26854 17930
rect 26796 17862 26808 17896
rect 26842 17862 26854 17896
rect 26796 17828 26854 17862
rect 26796 17794 26808 17828
rect 26842 17794 26854 17828
rect 26796 17760 26854 17794
rect 26796 17726 26808 17760
rect 26842 17726 26854 17760
rect 26796 17692 26854 17726
rect 26796 17658 26808 17692
rect 26842 17658 26854 17692
rect 26796 17624 26854 17658
rect 26796 17590 26808 17624
rect 26842 17590 26854 17624
rect 26796 17556 26854 17590
rect 26796 17522 26808 17556
rect 26842 17522 26854 17556
rect 26796 17488 26854 17522
rect 26796 17454 26808 17488
rect 26842 17454 26854 17488
rect 26796 17420 26854 17454
rect 26796 17386 26808 17420
rect 26842 17386 26854 17420
rect 26796 17352 26854 17386
rect 26796 17318 26808 17352
rect 26842 17318 26854 17352
rect 26796 17284 26854 17318
rect 26796 17250 26808 17284
rect 26842 17250 26854 17284
rect 26796 17216 26854 17250
rect 26796 17182 26808 17216
rect 26842 17182 26854 17216
rect 26796 17147 26854 17182
rect 27854 18712 27912 18747
rect 27854 18678 27866 18712
rect 27900 18678 27912 18712
rect 27854 18644 27912 18678
rect 27854 18610 27866 18644
rect 27900 18610 27912 18644
rect 27854 18576 27912 18610
rect 27854 18542 27866 18576
rect 27900 18542 27912 18576
rect 27854 18508 27912 18542
rect 27854 18474 27866 18508
rect 27900 18474 27912 18508
rect 27854 18440 27912 18474
rect 27854 18406 27866 18440
rect 27900 18406 27912 18440
rect 27854 18372 27912 18406
rect 27854 18338 27866 18372
rect 27900 18338 27912 18372
rect 27854 18304 27912 18338
rect 27854 18270 27866 18304
rect 27900 18270 27912 18304
rect 27854 18236 27912 18270
rect 27854 18202 27866 18236
rect 27900 18202 27912 18236
rect 27854 18168 27912 18202
rect 27854 18134 27866 18168
rect 27900 18134 27912 18168
rect 27854 18100 27912 18134
rect 27854 18066 27866 18100
rect 27900 18066 27912 18100
rect 27854 18032 27912 18066
rect 27854 17998 27866 18032
rect 27900 17998 27912 18032
rect 27854 17964 27912 17998
rect 27854 17930 27866 17964
rect 27900 17930 27912 17964
rect 27854 17896 27912 17930
rect 27854 17862 27866 17896
rect 27900 17862 27912 17896
rect 27854 17828 27912 17862
rect 27854 17794 27866 17828
rect 27900 17794 27912 17828
rect 27854 17760 27912 17794
rect 27854 17726 27866 17760
rect 27900 17726 27912 17760
rect 27854 17692 27912 17726
rect 27854 17658 27866 17692
rect 27900 17658 27912 17692
rect 27854 17624 27912 17658
rect 27854 17590 27866 17624
rect 27900 17590 27912 17624
rect 27854 17556 27912 17590
rect 27854 17522 27866 17556
rect 27900 17522 27912 17556
rect 27854 17488 27912 17522
rect 27854 17454 27866 17488
rect 27900 17454 27912 17488
rect 27854 17420 27912 17454
rect 27854 17386 27866 17420
rect 27900 17386 27912 17420
rect 27854 17352 27912 17386
rect 27854 17318 27866 17352
rect 27900 17318 27912 17352
rect 27854 17284 27912 17318
rect 27854 17250 27866 17284
rect 27900 17250 27912 17284
rect 27854 17216 27912 17250
rect 27854 17182 27866 17216
rect 27900 17182 27912 17216
rect 27854 17147 27912 17182
rect 39132 17933 39190 17974
rect 39132 17899 39144 17933
rect 39178 17899 39190 17933
rect 39132 17865 39190 17899
rect 39132 17831 39144 17865
rect 39178 17831 39190 17865
rect 39132 17797 39190 17831
rect 39132 17763 39144 17797
rect 39178 17763 39190 17797
rect 39132 17729 39190 17763
rect 39132 17695 39144 17729
rect 39178 17695 39190 17729
rect 39132 17661 39190 17695
rect 39132 17627 39144 17661
rect 39178 17627 39190 17661
rect 39132 17593 39190 17627
rect 39132 17559 39144 17593
rect 39178 17559 39190 17593
rect 39132 17525 39190 17559
rect 39132 17491 39144 17525
rect 39178 17491 39190 17525
rect 39132 17457 39190 17491
rect 39132 17423 39144 17457
rect 39178 17423 39190 17457
rect 39132 17389 39190 17423
rect 39132 17355 39144 17389
rect 39178 17355 39190 17389
rect 39132 17321 39190 17355
rect 39132 17287 39144 17321
rect 39178 17287 39190 17321
rect 39132 17253 39190 17287
rect 39132 17219 39144 17253
rect 39178 17219 39190 17253
rect 39132 17185 39190 17219
rect 39132 17151 39144 17185
rect 39178 17151 39190 17185
rect 39132 17117 39190 17151
rect 39132 17083 39144 17117
rect 39178 17083 39190 17117
rect 39132 17049 39190 17083
rect 39132 17015 39144 17049
rect 39178 17015 39190 17049
rect 39132 16974 39190 17015
rect 39390 17933 39448 17974
rect 39390 17899 39402 17933
rect 39436 17899 39448 17933
rect 39390 17865 39448 17899
rect 39390 17831 39402 17865
rect 39436 17831 39448 17865
rect 39390 17797 39448 17831
rect 39390 17763 39402 17797
rect 39436 17763 39448 17797
rect 39390 17729 39448 17763
rect 39390 17695 39402 17729
rect 39436 17695 39448 17729
rect 39390 17661 39448 17695
rect 39390 17627 39402 17661
rect 39436 17627 39448 17661
rect 39390 17593 39448 17627
rect 39390 17559 39402 17593
rect 39436 17559 39448 17593
rect 39390 17525 39448 17559
rect 39390 17491 39402 17525
rect 39436 17491 39448 17525
rect 39390 17457 39448 17491
rect 39390 17423 39402 17457
rect 39436 17423 39448 17457
rect 39390 17389 39448 17423
rect 39390 17355 39402 17389
rect 39436 17355 39448 17389
rect 39390 17321 39448 17355
rect 39390 17287 39402 17321
rect 39436 17287 39448 17321
rect 39390 17253 39448 17287
rect 39390 17219 39402 17253
rect 39436 17219 39448 17253
rect 39390 17185 39448 17219
rect 39390 17151 39402 17185
rect 39436 17151 39448 17185
rect 39390 17117 39448 17151
rect 39390 17083 39402 17117
rect 39436 17083 39448 17117
rect 39390 17049 39448 17083
rect 39390 17015 39402 17049
rect 39436 17015 39448 17049
rect 39390 16974 39448 17015
rect 39648 17933 39706 17974
rect 39648 17899 39660 17933
rect 39694 17899 39706 17933
rect 39648 17865 39706 17899
rect 39648 17831 39660 17865
rect 39694 17831 39706 17865
rect 39648 17797 39706 17831
rect 39648 17763 39660 17797
rect 39694 17763 39706 17797
rect 39648 17729 39706 17763
rect 39648 17695 39660 17729
rect 39694 17695 39706 17729
rect 39648 17661 39706 17695
rect 39648 17627 39660 17661
rect 39694 17627 39706 17661
rect 39648 17593 39706 17627
rect 39648 17559 39660 17593
rect 39694 17559 39706 17593
rect 39648 17525 39706 17559
rect 39648 17491 39660 17525
rect 39694 17491 39706 17525
rect 39648 17457 39706 17491
rect 39648 17423 39660 17457
rect 39694 17423 39706 17457
rect 39648 17389 39706 17423
rect 39648 17355 39660 17389
rect 39694 17355 39706 17389
rect 39648 17321 39706 17355
rect 39648 17287 39660 17321
rect 39694 17287 39706 17321
rect 39648 17253 39706 17287
rect 39648 17219 39660 17253
rect 39694 17219 39706 17253
rect 39648 17185 39706 17219
rect 39648 17151 39660 17185
rect 39694 17151 39706 17185
rect 39648 17117 39706 17151
rect 39648 17083 39660 17117
rect 39694 17083 39706 17117
rect 39648 17049 39706 17083
rect 39648 17015 39660 17049
rect 39694 17015 39706 17049
rect 39648 16974 39706 17015
rect 42600 18812 42658 18843
rect 42600 18778 42612 18812
rect 42646 18778 42658 18812
rect 42600 18744 42658 18778
rect 42600 18710 42612 18744
rect 42646 18710 42658 18744
rect 42600 18676 42658 18710
rect 42600 18642 42612 18676
rect 42646 18642 42658 18676
rect 42600 18608 42658 18642
rect 42600 18574 42612 18608
rect 42646 18574 42658 18608
rect 42600 18540 42658 18574
rect 42600 18506 42612 18540
rect 42646 18506 42658 18540
rect 42600 18472 42658 18506
rect 42600 18438 42612 18472
rect 42646 18438 42658 18472
rect 42600 18404 42658 18438
rect 42600 18370 42612 18404
rect 42646 18370 42658 18404
rect 42600 18336 42658 18370
rect 42600 18302 42612 18336
rect 42646 18302 42658 18336
rect 42600 18268 42658 18302
rect 42600 18234 42612 18268
rect 42646 18234 42658 18268
rect 42600 18200 42658 18234
rect 42600 18166 42612 18200
rect 42646 18166 42658 18200
rect 42600 18132 42658 18166
rect 42600 18098 42612 18132
rect 42646 18098 42658 18132
rect 42600 18064 42658 18098
rect 42600 18030 42612 18064
rect 42646 18030 42658 18064
rect 42600 17996 42658 18030
rect 42600 17962 42612 17996
rect 42646 17962 42658 17996
rect 42600 17928 42658 17962
rect 42600 17894 42612 17928
rect 42646 17894 42658 17928
rect 42600 17860 42658 17894
rect 42600 17826 42612 17860
rect 42646 17826 42658 17860
rect 42600 17792 42658 17826
rect 42600 17758 42612 17792
rect 42646 17758 42658 17792
rect 42600 17724 42658 17758
rect 42600 17690 42612 17724
rect 42646 17690 42658 17724
rect 42600 17656 42658 17690
rect 42600 17622 42612 17656
rect 42646 17622 42658 17656
rect 42600 17588 42658 17622
rect 42600 17554 42612 17588
rect 42646 17554 42658 17588
rect 42600 17520 42658 17554
rect 42600 17486 42612 17520
rect 42646 17486 42658 17520
rect 42600 17452 42658 17486
rect 42600 17418 42612 17452
rect 42646 17418 42658 17452
rect 42600 17384 42658 17418
rect 42600 17350 42612 17384
rect 42646 17350 42658 17384
rect 42600 17316 42658 17350
rect 42600 17282 42612 17316
rect 42646 17282 42658 17316
rect 42600 17248 42658 17282
rect 42600 17214 42612 17248
rect 42646 17214 42658 17248
rect 42600 17180 42658 17214
rect 42600 17146 42612 17180
rect 42646 17146 42658 17180
rect 42600 17112 42658 17146
rect 42600 17078 42612 17112
rect 42646 17078 42658 17112
rect 42600 17044 42658 17078
rect 42600 17010 42612 17044
rect 42646 17010 42658 17044
rect 42600 16976 42658 17010
rect 42600 16942 42612 16976
rect 42646 16942 42658 16976
rect 42600 16908 42658 16942
rect 42600 16874 42612 16908
rect 42646 16874 42658 16908
rect 42600 16843 42658 16874
rect 42858 18812 42916 18843
rect 42858 18778 42870 18812
rect 42904 18778 42916 18812
rect 42858 18744 42916 18778
rect 42858 18710 42870 18744
rect 42904 18710 42916 18744
rect 42858 18676 42916 18710
rect 42858 18642 42870 18676
rect 42904 18642 42916 18676
rect 42858 18608 42916 18642
rect 42858 18574 42870 18608
rect 42904 18574 42916 18608
rect 42858 18540 42916 18574
rect 42858 18506 42870 18540
rect 42904 18506 42916 18540
rect 42858 18472 42916 18506
rect 42858 18438 42870 18472
rect 42904 18438 42916 18472
rect 42858 18404 42916 18438
rect 42858 18370 42870 18404
rect 42904 18370 42916 18404
rect 42858 18336 42916 18370
rect 42858 18302 42870 18336
rect 42904 18302 42916 18336
rect 42858 18268 42916 18302
rect 42858 18234 42870 18268
rect 42904 18234 42916 18268
rect 42858 18200 42916 18234
rect 42858 18166 42870 18200
rect 42904 18166 42916 18200
rect 42858 18132 42916 18166
rect 42858 18098 42870 18132
rect 42904 18098 42916 18132
rect 42858 18064 42916 18098
rect 42858 18030 42870 18064
rect 42904 18030 42916 18064
rect 42858 17996 42916 18030
rect 42858 17962 42870 17996
rect 42904 17962 42916 17996
rect 42858 17928 42916 17962
rect 42858 17894 42870 17928
rect 42904 17894 42916 17928
rect 42858 17860 42916 17894
rect 42858 17826 42870 17860
rect 42904 17826 42916 17860
rect 42858 17792 42916 17826
rect 42858 17758 42870 17792
rect 42904 17758 42916 17792
rect 42858 17724 42916 17758
rect 42858 17690 42870 17724
rect 42904 17690 42916 17724
rect 42858 17656 42916 17690
rect 42858 17622 42870 17656
rect 42904 17622 42916 17656
rect 42858 17588 42916 17622
rect 42858 17554 42870 17588
rect 42904 17554 42916 17588
rect 42858 17520 42916 17554
rect 42858 17486 42870 17520
rect 42904 17486 42916 17520
rect 42858 17452 42916 17486
rect 42858 17418 42870 17452
rect 42904 17418 42916 17452
rect 42858 17384 42916 17418
rect 42858 17350 42870 17384
rect 42904 17350 42916 17384
rect 42858 17316 42916 17350
rect 42858 17282 42870 17316
rect 42904 17282 42916 17316
rect 42858 17248 42916 17282
rect 42858 17214 42870 17248
rect 42904 17214 42916 17248
rect 42858 17180 42916 17214
rect 42858 17146 42870 17180
rect 42904 17146 42916 17180
rect 42858 17112 42916 17146
rect 42858 17078 42870 17112
rect 42904 17078 42916 17112
rect 42858 17044 42916 17078
rect 42858 17010 42870 17044
rect 42904 17010 42916 17044
rect 42858 16976 42916 17010
rect 42858 16942 42870 16976
rect 42904 16942 42916 16976
rect 42858 16908 42916 16942
rect 42858 16874 42870 16908
rect 42904 16874 42916 16908
rect 42858 16843 42916 16874
rect 43116 18812 43174 18843
rect 43116 18778 43128 18812
rect 43162 18778 43174 18812
rect 43116 18744 43174 18778
rect 43116 18710 43128 18744
rect 43162 18710 43174 18744
rect 43116 18676 43174 18710
rect 43116 18642 43128 18676
rect 43162 18642 43174 18676
rect 43116 18608 43174 18642
rect 43116 18574 43128 18608
rect 43162 18574 43174 18608
rect 43116 18540 43174 18574
rect 43116 18506 43128 18540
rect 43162 18506 43174 18540
rect 43116 18472 43174 18506
rect 43116 18438 43128 18472
rect 43162 18438 43174 18472
rect 43116 18404 43174 18438
rect 43116 18370 43128 18404
rect 43162 18370 43174 18404
rect 43116 18336 43174 18370
rect 43116 18302 43128 18336
rect 43162 18302 43174 18336
rect 43116 18268 43174 18302
rect 43116 18234 43128 18268
rect 43162 18234 43174 18268
rect 43116 18200 43174 18234
rect 43116 18166 43128 18200
rect 43162 18166 43174 18200
rect 43116 18132 43174 18166
rect 43116 18098 43128 18132
rect 43162 18098 43174 18132
rect 43116 18064 43174 18098
rect 43116 18030 43128 18064
rect 43162 18030 43174 18064
rect 43116 17996 43174 18030
rect 43116 17962 43128 17996
rect 43162 17962 43174 17996
rect 43116 17928 43174 17962
rect 43116 17894 43128 17928
rect 43162 17894 43174 17928
rect 43116 17860 43174 17894
rect 43116 17826 43128 17860
rect 43162 17826 43174 17860
rect 43116 17792 43174 17826
rect 43116 17758 43128 17792
rect 43162 17758 43174 17792
rect 43116 17724 43174 17758
rect 43116 17690 43128 17724
rect 43162 17690 43174 17724
rect 43116 17656 43174 17690
rect 43116 17622 43128 17656
rect 43162 17622 43174 17656
rect 43116 17588 43174 17622
rect 43116 17554 43128 17588
rect 43162 17554 43174 17588
rect 43116 17520 43174 17554
rect 43116 17486 43128 17520
rect 43162 17486 43174 17520
rect 43116 17452 43174 17486
rect 43116 17418 43128 17452
rect 43162 17418 43174 17452
rect 43116 17384 43174 17418
rect 43116 17350 43128 17384
rect 43162 17350 43174 17384
rect 43116 17316 43174 17350
rect 43116 17282 43128 17316
rect 43162 17282 43174 17316
rect 43116 17248 43174 17282
rect 43116 17214 43128 17248
rect 43162 17214 43174 17248
rect 43116 17180 43174 17214
rect 43116 17146 43128 17180
rect 43162 17146 43174 17180
rect 43116 17112 43174 17146
rect 43116 17078 43128 17112
rect 43162 17078 43174 17112
rect 43116 17044 43174 17078
rect 43116 17010 43128 17044
rect 43162 17010 43174 17044
rect 43116 16976 43174 17010
rect 43116 16942 43128 16976
rect 43162 16942 43174 16976
rect 43116 16908 43174 16942
rect 43116 16874 43128 16908
rect 43162 16874 43174 16908
rect 43116 16843 43174 16874
rect 43374 18812 43432 18843
rect 43374 18778 43386 18812
rect 43420 18778 43432 18812
rect 43374 18744 43432 18778
rect 43374 18710 43386 18744
rect 43420 18710 43432 18744
rect 43374 18676 43432 18710
rect 43374 18642 43386 18676
rect 43420 18642 43432 18676
rect 43374 18608 43432 18642
rect 43374 18574 43386 18608
rect 43420 18574 43432 18608
rect 43374 18540 43432 18574
rect 43374 18506 43386 18540
rect 43420 18506 43432 18540
rect 43374 18472 43432 18506
rect 43374 18438 43386 18472
rect 43420 18438 43432 18472
rect 43374 18404 43432 18438
rect 43374 18370 43386 18404
rect 43420 18370 43432 18404
rect 43374 18336 43432 18370
rect 43374 18302 43386 18336
rect 43420 18302 43432 18336
rect 43374 18268 43432 18302
rect 43374 18234 43386 18268
rect 43420 18234 43432 18268
rect 43374 18200 43432 18234
rect 43374 18166 43386 18200
rect 43420 18166 43432 18200
rect 43374 18132 43432 18166
rect 43374 18098 43386 18132
rect 43420 18098 43432 18132
rect 43374 18064 43432 18098
rect 43374 18030 43386 18064
rect 43420 18030 43432 18064
rect 43374 17996 43432 18030
rect 43374 17962 43386 17996
rect 43420 17962 43432 17996
rect 43374 17928 43432 17962
rect 43374 17894 43386 17928
rect 43420 17894 43432 17928
rect 43374 17860 43432 17894
rect 43374 17826 43386 17860
rect 43420 17826 43432 17860
rect 43374 17792 43432 17826
rect 43374 17758 43386 17792
rect 43420 17758 43432 17792
rect 43374 17724 43432 17758
rect 43374 17690 43386 17724
rect 43420 17690 43432 17724
rect 43374 17656 43432 17690
rect 43374 17622 43386 17656
rect 43420 17622 43432 17656
rect 43374 17588 43432 17622
rect 43374 17554 43386 17588
rect 43420 17554 43432 17588
rect 43374 17520 43432 17554
rect 43374 17486 43386 17520
rect 43420 17486 43432 17520
rect 43374 17452 43432 17486
rect 43374 17418 43386 17452
rect 43420 17418 43432 17452
rect 43374 17384 43432 17418
rect 43374 17350 43386 17384
rect 43420 17350 43432 17384
rect 43374 17316 43432 17350
rect 43374 17282 43386 17316
rect 43420 17282 43432 17316
rect 43374 17248 43432 17282
rect 43374 17214 43386 17248
rect 43420 17214 43432 17248
rect 43374 17180 43432 17214
rect 43374 17146 43386 17180
rect 43420 17146 43432 17180
rect 43374 17112 43432 17146
rect 43374 17078 43386 17112
rect 43420 17078 43432 17112
rect 43374 17044 43432 17078
rect 43374 17010 43386 17044
rect 43420 17010 43432 17044
rect 43374 16976 43432 17010
rect 43374 16942 43386 16976
rect 43420 16942 43432 16976
rect 43374 16908 43432 16942
rect 43374 16874 43386 16908
rect 43420 16874 43432 16908
rect 43374 16843 43432 16874
rect 43632 18812 43690 18843
rect 43632 18778 43644 18812
rect 43678 18778 43690 18812
rect 43632 18744 43690 18778
rect 43632 18710 43644 18744
rect 43678 18710 43690 18744
rect 43632 18676 43690 18710
rect 43632 18642 43644 18676
rect 43678 18642 43690 18676
rect 43632 18608 43690 18642
rect 43632 18574 43644 18608
rect 43678 18574 43690 18608
rect 43632 18540 43690 18574
rect 43632 18506 43644 18540
rect 43678 18506 43690 18540
rect 43632 18472 43690 18506
rect 43632 18438 43644 18472
rect 43678 18438 43690 18472
rect 43632 18404 43690 18438
rect 43632 18370 43644 18404
rect 43678 18370 43690 18404
rect 43632 18336 43690 18370
rect 43632 18302 43644 18336
rect 43678 18302 43690 18336
rect 43632 18268 43690 18302
rect 43632 18234 43644 18268
rect 43678 18234 43690 18268
rect 43632 18200 43690 18234
rect 43632 18166 43644 18200
rect 43678 18166 43690 18200
rect 43632 18132 43690 18166
rect 43632 18098 43644 18132
rect 43678 18098 43690 18132
rect 43632 18064 43690 18098
rect 43632 18030 43644 18064
rect 43678 18030 43690 18064
rect 43632 17996 43690 18030
rect 43632 17962 43644 17996
rect 43678 17962 43690 17996
rect 43632 17928 43690 17962
rect 43632 17894 43644 17928
rect 43678 17894 43690 17928
rect 43632 17860 43690 17894
rect 43632 17826 43644 17860
rect 43678 17826 43690 17860
rect 43632 17792 43690 17826
rect 43632 17758 43644 17792
rect 43678 17758 43690 17792
rect 43632 17724 43690 17758
rect 43632 17690 43644 17724
rect 43678 17690 43690 17724
rect 43632 17656 43690 17690
rect 43632 17622 43644 17656
rect 43678 17622 43690 17656
rect 43632 17588 43690 17622
rect 43632 17554 43644 17588
rect 43678 17554 43690 17588
rect 43632 17520 43690 17554
rect 43632 17486 43644 17520
rect 43678 17486 43690 17520
rect 43632 17452 43690 17486
rect 43632 17418 43644 17452
rect 43678 17418 43690 17452
rect 43632 17384 43690 17418
rect 43632 17350 43644 17384
rect 43678 17350 43690 17384
rect 43632 17316 43690 17350
rect 43632 17282 43644 17316
rect 43678 17282 43690 17316
rect 43632 17248 43690 17282
rect 43632 17214 43644 17248
rect 43678 17214 43690 17248
rect 43632 17180 43690 17214
rect 43632 17146 43644 17180
rect 43678 17146 43690 17180
rect 43632 17112 43690 17146
rect 43632 17078 43644 17112
rect 43678 17078 43690 17112
rect 43632 17044 43690 17078
rect 43632 17010 43644 17044
rect 43678 17010 43690 17044
rect 43632 16976 43690 17010
rect 43632 16942 43644 16976
rect 43678 16942 43690 16976
rect 43632 16908 43690 16942
rect 43632 16874 43644 16908
rect 43678 16874 43690 16908
rect 43632 16843 43690 16874
rect 43890 18812 43948 18843
rect 43890 18778 43902 18812
rect 43936 18778 43948 18812
rect 43890 18744 43948 18778
rect 43890 18710 43902 18744
rect 43936 18710 43948 18744
rect 43890 18676 43948 18710
rect 43890 18642 43902 18676
rect 43936 18642 43948 18676
rect 43890 18608 43948 18642
rect 43890 18574 43902 18608
rect 43936 18574 43948 18608
rect 43890 18540 43948 18574
rect 43890 18506 43902 18540
rect 43936 18506 43948 18540
rect 43890 18472 43948 18506
rect 43890 18438 43902 18472
rect 43936 18438 43948 18472
rect 43890 18404 43948 18438
rect 43890 18370 43902 18404
rect 43936 18370 43948 18404
rect 43890 18336 43948 18370
rect 43890 18302 43902 18336
rect 43936 18302 43948 18336
rect 43890 18268 43948 18302
rect 43890 18234 43902 18268
rect 43936 18234 43948 18268
rect 43890 18200 43948 18234
rect 43890 18166 43902 18200
rect 43936 18166 43948 18200
rect 43890 18132 43948 18166
rect 43890 18098 43902 18132
rect 43936 18098 43948 18132
rect 43890 18064 43948 18098
rect 43890 18030 43902 18064
rect 43936 18030 43948 18064
rect 43890 17996 43948 18030
rect 43890 17962 43902 17996
rect 43936 17962 43948 17996
rect 43890 17928 43948 17962
rect 43890 17894 43902 17928
rect 43936 17894 43948 17928
rect 43890 17860 43948 17894
rect 43890 17826 43902 17860
rect 43936 17826 43948 17860
rect 43890 17792 43948 17826
rect 43890 17758 43902 17792
rect 43936 17758 43948 17792
rect 43890 17724 43948 17758
rect 43890 17690 43902 17724
rect 43936 17690 43948 17724
rect 43890 17656 43948 17690
rect 43890 17622 43902 17656
rect 43936 17622 43948 17656
rect 43890 17588 43948 17622
rect 43890 17554 43902 17588
rect 43936 17554 43948 17588
rect 43890 17520 43948 17554
rect 43890 17486 43902 17520
rect 43936 17486 43948 17520
rect 43890 17452 43948 17486
rect 43890 17418 43902 17452
rect 43936 17418 43948 17452
rect 43890 17384 43948 17418
rect 43890 17350 43902 17384
rect 43936 17350 43948 17384
rect 43890 17316 43948 17350
rect 43890 17282 43902 17316
rect 43936 17282 43948 17316
rect 43890 17248 43948 17282
rect 43890 17214 43902 17248
rect 43936 17214 43948 17248
rect 43890 17180 43948 17214
rect 43890 17146 43902 17180
rect 43936 17146 43948 17180
rect 43890 17112 43948 17146
rect 43890 17078 43902 17112
rect 43936 17078 43948 17112
rect 43890 17044 43948 17078
rect 43890 17010 43902 17044
rect 43936 17010 43948 17044
rect 43890 16976 43948 17010
rect 43890 16942 43902 16976
rect 43936 16942 43948 16976
rect 43890 16908 43948 16942
rect 43890 16874 43902 16908
rect 43936 16874 43948 16908
rect 43890 16843 43948 16874
rect 44148 18812 44206 18843
rect 44148 18778 44160 18812
rect 44194 18778 44206 18812
rect 44148 18744 44206 18778
rect 44148 18710 44160 18744
rect 44194 18710 44206 18744
rect 44148 18676 44206 18710
rect 44148 18642 44160 18676
rect 44194 18642 44206 18676
rect 44148 18608 44206 18642
rect 44148 18574 44160 18608
rect 44194 18574 44206 18608
rect 44148 18540 44206 18574
rect 44148 18506 44160 18540
rect 44194 18506 44206 18540
rect 44148 18472 44206 18506
rect 44148 18438 44160 18472
rect 44194 18438 44206 18472
rect 44148 18404 44206 18438
rect 44148 18370 44160 18404
rect 44194 18370 44206 18404
rect 44148 18336 44206 18370
rect 44148 18302 44160 18336
rect 44194 18302 44206 18336
rect 44148 18268 44206 18302
rect 44148 18234 44160 18268
rect 44194 18234 44206 18268
rect 44148 18200 44206 18234
rect 44148 18166 44160 18200
rect 44194 18166 44206 18200
rect 44148 18132 44206 18166
rect 44148 18098 44160 18132
rect 44194 18098 44206 18132
rect 44148 18064 44206 18098
rect 44148 18030 44160 18064
rect 44194 18030 44206 18064
rect 44148 17996 44206 18030
rect 44148 17962 44160 17996
rect 44194 17962 44206 17996
rect 44148 17928 44206 17962
rect 44148 17894 44160 17928
rect 44194 17894 44206 17928
rect 44148 17860 44206 17894
rect 44148 17826 44160 17860
rect 44194 17826 44206 17860
rect 44148 17792 44206 17826
rect 44148 17758 44160 17792
rect 44194 17758 44206 17792
rect 44148 17724 44206 17758
rect 44148 17690 44160 17724
rect 44194 17690 44206 17724
rect 44148 17656 44206 17690
rect 44148 17622 44160 17656
rect 44194 17622 44206 17656
rect 44148 17588 44206 17622
rect 44148 17554 44160 17588
rect 44194 17554 44206 17588
rect 44148 17520 44206 17554
rect 44148 17486 44160 17520
rect 44194 17486 44206 17520
rect 44148 17452 44206 17486
rect 44148 17418 44160 17452
rect 44194 17418 44206 17452
rect 44148 17384 44206 17418
rect 44148 17350 44160 17384
rect 44194 17350 44206 17384
rect 44148 17316 44206 17350
rect 44148 17282 44160 17316
rect 44194 17282 44206 17316
rect 44148 17248 44206 17282
rect 44148 17214 44160 17248
rect 44194 17214 44206 17248
rect 44148 17180 44206 17214
rect 44148 17146 44160 17180
rect 44194 17146 44206 17180
rect 44148 17112 44206 17146
rect 44148 17078 44160 17112
rect 44194 17078 44206 17112
rect 44148 17044 44206 17078
rect 44148 17010 44160 17044
rect 44194 17010 44206 17044
rect 44148 16976 44206 17010
rect 44148 16942 44160 16976
rect 44194 16942 44206 16976
rect 44148 16908 44206 16942
rect 44148 16874 44160 16908
rect 44194 16874 44206 16908
rect 44148 16843 44206 16874
rect 44406 18812 44464 18843
rect 44406 18778 44418 18812
rect 44452 18778 44464 18812
rect 44406 18744 44464 18778
rect 44406 18710 44418 18744
rect 44452 18710 44464 18744
rect 44406 18676 44464 18710
rect 44406 18642 44418 18676
rect 44452 18642 44464 18676
rect 44406 18608 44464 18642
rect 44406 18574 44418 18608
rect 44452 18574 44464 18608
rect 44406 18540 44464 18574
rect 44406 18506 44418 18540
rect 44452 18506 44464 18540
rect 44406 18472 44464 18506
rect 44406 18438 44418 18472
rect 44452 18438 44464 18472
rect 44406 18404 44464 18438
rect 44406 18370 44418 18404
rect 44452 18370 44464 18404
rect 44406 18336 44464 18370
rect 44406 18302 44418 18336
rect 44452 18302 44464 18336
rect 44406 18268 44464 18302
rect 44406 18234 44418 18268
rect 44452 18234 44464 18268
rect 44406 18200 44464 18234
rect 44406 18166 44418 18200
rect 44452 18166 44464 18200
rect 44406 18132 44464 18166
rect 44406 18098 44418 18132
rect 44452 18098 44464 18132
rect 44406 18064 44464 18098
rect 44406 18030 44418 18064
rect 44452 18030 44464 18064
rect 44406 17996 44464 18030
rect 44406 17962 44418 17996
rect 44452 17962 44464 17996
rect 44406 17928 44464 17962
rect 44406 17894 44418 17928
rect 44452 17894 44464 17928
rect 44406 17860 44464 17894
rect 44406 17826 44418 17860
rect 44452 17826 44464 17860
rect 44406 17792 44464 17826
rect 44406 17758 44418 17792
rect 44452 17758 44464 17792
rect 44406 17724 44464 17758
rect 44406 17690 44418 17724
rect 44452 17690 44464 17724
rect 44406 17656 44464 17690
rect 44406 17622 44418 17656
rect 44452 17622 44464 17656
rect 44406 17588 44464 17622
rect 44406 17554 44418 17588
rect 44452 17554 44464 17588
rect 44406 17520 44464 17554
rect 44406 17486 44418 17520
rect 44452 17486 44464 17520
rect 44406 17452 44464 17486
rect 44406 17418 44418 17452
rect 44452 17418 44464 17452
rect 44406 17384 44464 17418
rect 44406 17350 44418 17384
rect 44452 17350 44464 17384
rect 44406 17316 44464 17350
rect 44406 17282 44418 17316
rect 44452 17282 44464 17316
rect 44406 17248 44464 17282
rect 44406 17214 44418 17248
rect 44452 17214 44464 17248
rect 44406 17180 44464 17214
rect 44406 17146 44418 17180
rect 44452 17146 44464 17180
rect 44406 17112 44464 17146
rect 44406 17078 44418 17112
rect 44452 17078 44464 17112
rect 44406 17044 44464 17078
rect 44406 17010 44418 17044
rect 44452 17010 44464 17044
rect 44406 16976 44464 17010
rect 44406 16942 44418 16976
rect 44452 16942 44464 16976
rect 44406 16908 44464 16942
rect 44406 16874 44418 16908
rect 44452 16874 44464 16908
rect 44406 16843 44464 16874
rect 44664 18812 44722 18843
rect 44664 18778 44676 18812
rect 44710 18778 44722 18812
rect 44664 18744 44722 18778
rect 44664 18710 44676 18744
rect 44710 18710 44722 18744
rect 44664 18676 44722 18710
rect 44664 18642 44676 18676
rect 44710 18642 44722 18676
rect 44664 18608 44722 18642
rect 44664 18574 44676 18608
rect 44710 18574 44722 18608
rect 44664 18540 44722 18574
rect 44664 18506 44676 18540
rect 44710 18506 44722 18540
rect 44664 18472 44722 18506
rect 44664 18438 44676 18472
rect 44710 18438 44722 18472
rect 44664 18404 44722 18438
rect 44664 18370 44676 18404
rect 44710 18370 44722 18404
rect 44664 18336 44722 18370
rect 44664 18302 44676 18336
rect 44710 18302 44722 18336
rect 44664 18268 44722 18302
rect 44664 18234 44676 18268
rect 44710 18234 44722 18268
rect 44664 18200 44722 18234
rect 44664 18166 44676 18200
rect 44710 18166 44722 18200
rect 44664 18132 44722 18166
rect 44664 18098 44676 18132
rect 44710 18098 44722 18132
rect 44664 18064 44722 18098
rect 44664 18030 44676 18064
rect 44710 18030 44722 18064
rect 44664 17996 44722 18030
rect 44664 17962 44676 17996
rect 44710 17962 44722 17996
rect 44664 17928 44722 17962
rect 44664 17894 44676 17928
rect 44710 17894 44722 17928
rect 44664 17860 44722 17894
rect 44664 17826 44676 17860
rect 44710 17826 44722 17860
rect 44664 17792 44722 17826
rect 44664 17758 44676 17792
rect 44710 17758 44722 17792
rect 44664 17724 44722 17758
rect 44664 17690 44676 17724
rect 44710 17690 44722 17724
rect 44664 17656 44722 17690
rect 44664 17622 44676 17656
rect 44710 17622 44722 17656
rect 44664 17588 44722 17622
rect 44664 17554 44676 17588
rect 44710 17554 44722 17588
rect 44664 17520 44722 17554
rect 44664 17486 44676 17520
rect 44710 17486 44722 17520
rect 44664 17452 44722 17486
rect 44664 17418 44676 17452
rect 44710 17418 44722 17452
rect 44664 17384 44722 17418
rect 44664 17350 44676 17384
rect 44710 17350 44722 17384
rect 44664 17316 44722 17350
rect 44664 17282 44676 17316
rect 44710 17282 44722 17316
rect 44664 17248 44722 17282
rect 44664 17214 44676 17248
rect 44710 17214 44722 17248
rect 44664 17180 44722 17214
rect 44664 17146 44676 17180
rect 44710 17146 44722 17180
rect 44664 17112 44722 17146
rect 44664 17078 44676 17112
rect 44710 17078 44722 17112
rect 44664 17044 44722 17078
rect 44664 17010 44676 17044
rect 44710 17010 44722 17044
rect 44664 16976 44722 17010
rect 44664 16942 44676 16976
rect 44710 16942 44722 16976
rect 44664 16908 44722 16942
rect 44664 16874 44676 16908
rect 44710 16874 44722 16908
rect 44664 16843 44722 16874
rect 44922 18812 44980 18843
rect 44922 18778 44934 18812
rect 44968 18778 44980 18812
rect 44922 18744 44980 18778
rect 44922 18710 44934 18744
rect 44968 18710 44980 18744
rect 44922 18676 44980 18710
rect 44922 18642 44934 18676
rect 44968 18642 44980 18676
rect 44922 18608 44980 18642
rect 44922 18574 44934 18608
rect 44968 18574 44980 18608
rect 44922 18540 44980 18574
rect 44922 18506 44934 18540
rect 44968 18506 44980 18540
rect 44922 18472 44980 18506
rect 44922 18438 44934 18472
rect 44968 18438 44980 18472
rect 44922 18404 44980 18438
rect 44922 18370 44934 18404
rect 44968 18370 44980 18404
rect 44922 18336 44980 18370
rect 44922 18302 44934 18336
rect 44968 18302 44980 18336
rect 44922 18268 44980 18302
rect 44922 18234 44934 18268
rect 44968 18234 44980 18268
rect 44922 18200 44980 18234
rect 44922 18166 44934 18200
rect 44968 18166 44980 18200
rect 44922 18132 44980 18166
rect 44922 18098 44934 18132
rect 44968 18098 44980 18132
rect 44922 18064 44980 18098
rect 44922 18030 44934 18064
rect 44968 18030 44980 18064
rect 44922 17996 44980 18030
rect 44922 17962 44934 17996
rect 44968 17962 44980 17996
rect 44922 17928 44980 17962
rect 44922 17894 44934 17928
rect 44968 17894 44980 17928
rect 44922 17860 44980 17894
rect 44922 17826 44934 17860
rect 44968 17826 44980 17860
rect 44922 17792 44980 17826
rect 44922 17758 44934 17792
rect 44968 17758 44980 17792
rect 44922 17724 44980 17758
rect 44922 17690 44934 17724
rect 44968 17690 44980 17724
rect 44922 17656 44980 17690
rect 44922 17622 44934 17656
rect 44968 17622 44980 17656
rect 44922 17588 44980 17622
rect 44922 17554 44934 17588
rect 44968 17554 44980 17588
rect 44922 17520 44980 17554
rect 44922 17486 44934 17520
rect 44968 17486 44980 17520
rect 44922 17452 44980 17486
rect 44922 17418 44934 17452
rect 44968 17418 44980 17452
rect 44922 17384 44980 17418
rect 44922 17350 44934 17384
rect 44968 17350 44980 17384
rect 44922 17316 44980 17350
rect 44922 17282 44934 17316
rect 44968 17282 44980 17316
rect 44922 17248 44980 17282
rect 44922 17214 44934 17248
rect 44968 17214 44980 17248
rect 44922 17180 44980 17214
rect 44922 17146 44934 17180
rect 44968 17146 44980 17180
rect 44922 17112 44980 17146
rect 44922 17078 44934 17112
rect 44968 17078 44980 17112
rect 44922 17044 44980 17078
rect 44922 17010 44934 17044
rect 44968 17010 44980 17044
rect 44922 16976 44980 17010
rect 44922 16942 44934 16976
rect 44968 16942 44980 16976
rect 44922 16908 44980 16942
rect 44922 16874 44934 16908
rect 44968 16874 44980 16908
rect 44922 16843 44980 16874
rect 45180 18812 45238 18843
rect 45180 18778 45192 18812
rect 45226 18778 45238 18812
rect 45180 18744 45238 18778
rect 45180 18710 45192 18744
rect 45226 18710 45238 18744
rect 45180 18676 45238 18710
rect 45180 18642 45192 18676
rect 45226 18642 45238 18676
rect 45180 18608 45238 18642
rect 45180 18574 45192 18608
rect 45226 18574 45238 18608
rect 45180 18540 45238 18574
rect 45180 18506 45192 18540
rect 45226 18506 45238 18540
rect 45180 18472 45238 18506
rect 45180 18438 45192 18472
rect 45226 18438 45238 18472
rect 45180 18404 45238 18438
rect 45180 18370 45192 18404
rect 45226 18370 45238 18404
rect 45180 18336 45238 18370
rect 45180 18302 45192 18336
rect 45226 18302 45238 18336
rect 45180 18268 45238 18302
rect 45180 18234 45192 18268
rect 45226 18234 45238 18268
rect 45180 18200 45238 18234
rect 45180 18166 45192 18200
rect 45226 18166 45238 18200
rect 45180 18132 45238 18166
rect 45180 18098 45192 18132
rect 45226 18098 45238 18132
rect 45180 18064 45238 18098
rect 45180 18030 45192 18064
rect 45226 18030 45238 18064
rect 45180 17996 45238 18030
rect 45180 17962 45192 17996
rect 45226 17962 45238 17996
rect 45180 17928 45238 17962
rect 45180 17894 45192 17928
rect 45226 17894 45238 17928
rect 45180 17860 45238 17894
rect 45180 17826 45192 17860
rect 45226 17826 45238 17860
rect 45180 17792 45238 17826
rect 45180 17758 45192 17792
rect 45226 17758 45238 17792
rect 45180 17724 45238 17758
rect 45180 17690 45192 17724
rect 45226 17690 45238 17724
rect 45180 17656 45238 17690
rect 45180 17622 45192 17656
rect 45226 17622 45238 17656
rect 45180 17588 45238 17622
rect 45180 17554 45192 17588
rect 45226 17554 45238 17588
rect 45180 17520 45238 17554
rect 45180 17486 45192 17520
rect 45226 17486 45238 17520
rect 45180 17452 45238 17486
rect 45180 17418 45192 17452
rect 45226 17418 45238 17452
rect 45180 17384 45238 17418
rect 45180 17350 45192 17384
rect 45226 17350 45238 17384
rect 45180 17316 45238 17350
rect 45180 17282 45192 17316
rect 45226 17282 45238 17316
rect 45180 17248 45238 17282
rect 45180 17214 45192 17248
rect 45226 17214 45238 17248
rect 45180 17180 45238 17214
rect 45180 17146 45192 17180
rect 45226 17146 45238 17180
rect 45180 17112 45238 17146
rect 45180 17078 45192 17112
rect 45226 17078 45238 17112
rect 45180 17044 45238 17078
rect 45180 17010 45192 17044
rect 45226 17010 45238 17044
rect 45180 16976 45238 17010
rect 45180 16942 45192 16976
rect 45226 16942 45238 16976
rect 45180 16908 45238 16942
rect 45180 16874 45192 16908
rect 45226 16874 45238 16908
rect 45180 16843 45238 16874
rect 12982 14746 13040 14767
rect 12982 14712 12994 14746
rect 13028 14712 13040 14746
rect 12982 14678 13040 14712
rect 12982 14644 12994 14678
rect 13028 14644 13040 14678
rect 12982 14610 13040 14644
rect 12982 14576 12994 14610
rect 13028 14576 13040 14610
rect 12982 14542 13040 14576
rect 12982 14508 12994 14542
rect 13028 14508 13040 14542
rect 12982 14474 13040 14508
rect 12982 14440 12994 14474
rect 13028 14440 13040 14474
rect 12982 14406 13040 14440
rect 12982 14372 12994 14406
rect 13028 14372 13040 14406
rect 12982 14338 13040 14372
rect 12982 14304 12994 14338
rect 13028 14304 13040 14338
rect 12982 14270 13040 14304
rect 12982 14236 12994 14270
rect 13028 14236 13040 14270
rect 12982 14202 13040 14236
rect 12982 14168 12994 14202
rect 13028 14168 13040 14202
rect 12982 14134 13040 14168
rect 12982 14100 12994 14134
rect 13028 14100 13040 14134
rect 12982 14066 13040 14100
rect 12982 14032 12994 14066
rect 13028 14032 13040 14066
rect 12982 13998 13040 14032
rect 12982 13964 12994 13998
rect 13028 13964 13040 13998
rect 12982 13930 13040 13964
rect 12982 13896 12994 13930
rect 13028 13896 13040 13930
rect 12982 13862 13040 13896
rect 12982 13828 12994 13862
rect 13028 13828 13040 13862
rect 12982 13794 13040 13828
rect 12982 13760 12994 13794
rect 13028 13760 13040 13794
rect 12982 13726 13040 13760
rect 12982 13692 12994 13726
rect 13028 13692 13040 13726
rect 12982 13658 13040 13692
rect 12982 13624 12994 13658
rect 13028 13624 13040 13658
rect 12982 13590 13040 13624
rect 12982 13556 12994 13590
rect 13028 13556 13040 13590
rect 12982 13522 13040 13556
rect 12982 13488 12994 13522
rect 13028 13488 13040 13522
rect 12982 13454 13040 13488
rect 12982 13420 12994 13454
rect 13028 13420 13040 13454
rect 12982 13386 13040 13420
rect 12982 13352 12994 13386
rect 13028 13352 13040 13386
rect 12982 13318 13040 13352
rect 12982 13284 12994 13318
rect 13028 13284 13040 13318
rect 12982 13250 13040 13284
rect 12982 13216 12994 13250
rect 13028 13216 13040 13250
rect 12982 13182 13040 13216
rect 12982 13148 12994 13182
rect 13028 13148 13040 13182
rect 12982 13114 13040 13148
rect 12982 13080 12994 13114
rect 13028 13080 13040 13114
rect 12982 13046 13040 13080
rect 12982 13012 12994 13046
rect 13028 13012 13040 13046
rect 12982 12978 13040 13012
rect 12982 12944 12994 12978
rect 13028 12944 13040 12978
rect 12982 12910 13040 12944
rect 12982 12876 12994 12910
rect 13028 12876 13040 12910
rect 12982 12842 13040 12876
rect 12982 12808 12994 12842
rect 13028 12808 13040 12842
rect 12982 12774 13040 12808
rect 12982 12740 12994 12774
rect 13028 12740 13040 12774
rect 12982 12706 13040 12740
rect 12982 12672 12994 12706
rect 13028 12672 13040 12706
rect 12982 12638 13040 12672
rect 12982 12604 12994 12638
rect 13028 12604 13040 12638
rect 12982 12570 13040 12604
rect 12982 12536 12994 12570
rect 13028 12536 13040 12570
rect 12982 12502 13040 12536
rect 12982 12468 12994 12502
rect 13028 12468 13040 12502
rect 12982 12434 13040 12468
rect 12982 12400 12994 12434
rect 13028 12400 13040 12434
rect 12982 12366 13040 12400
rect 12982 12332 12994 12366
rect 13028 12332 13040 12366
rect 12982 12298 13040 12332
rect 12982 12264 12994 12298
rect 13028 12264 13040 12298
rect 12982 12230 13040 12264
rect 12982 12196 12994 12230
rect 13028 12196 13040 12230
rect 12982 12162 13040 12196
rect 12982 12128 12994 12162
rect 13028 12128 13040 12162
rect 12982 12094 13040 12128
rect 12982 12060 12994 12094
rect 13028 12060 13040 12094
rect 12982 12026 13040 12060
rect 12982 11992 12994 12026
rect 13028 11992 13040 12026
rect 12982 11958 13040 11992
rect 12982 11924 12994 11958
rect 13028 11924 13040 11958
rect 12982 11890 13040 11924
rect 12982 11856 12994 11890
rect 13028 11856 13040 11890
rect 12982 11822 13040 11856
rect 12982 11788 12994 11822
rect 13028 11788 13040 11822
rect 12982 11767 13040 11788
rect 14040 14746 14098 14767
rect 14040 14712 14052 14746
rect 14086 14712 14098 14746
rect 14040 14678 14098 14712
rect 14040 14644 14052 14678
rect 14086 14644 14098 14678
rect 14040 14610 14098 14644
rect 14040 14576 14052 14610
rect 14086 14576 14098 14610
rect 14040 14542 14098 14576
rect 14040 14508 14052 14542
rect 14086 14508 14098 14542
rect 14040 14474 14098 14508
rect 14040 14440 14052 14474
rect 14086 14440 14098 14474
rect 14040 14406 14098 14440
rect 14040 14372 14052 14406
rect 14086 14372 14098 14406
rect 14040 14338 14098 14372
rect 14040 14304 14052 14338
rect 14086 14304 14098 14338
rect 14040 14270 14098 14304
rect 14040 14236 14052 14270
rect 14086 14236 14098 14270
rect 14040 14202 14098 14236
rect 14040 14168 14052 14202
rect 14086 14168 14098 14202
rect 14040 14134 14098 14168
rect 14040 14100 14052 14134
rect 14086 14100 14098 14134
rect 14040 14066 14098 14100
rect 14040 14032 14052 14066
rect 14086 14032 14098 14066
rect 14040 13998 14098 14032
rect 14040 13964 14052 13998
rect 14086 13964 14098 13998
rect 14040 13930 14098 13964
rect 14040 13896 14052 13930
rect 14086 13896 14098 13930
rect 14040 13862 14098 13896
rect 14040 13828 14052 13862
rect 14086 13828 14098 13862
rect 14040 13794 14098 13828
rect 14040 13760 14052 13794
rect 14086 13760 14098 13794
rect 14040 13726 14098 13760
rect 14040 13692 14052 13726
rect 14086 13692 14098 13726
rect 14040 13658 14098 13692
rect 14040 13624 14052 13658
rect 14086 13624 14098 13658
rect 14040 13590 14098 13624
rect 14040 13556 14052 13590
rect 14086 13556 14098 13590
rect 14040 13522 14098 13556
rect 14040 13488 14052 13522
rect 14086 13488 14098 13522
rect 14040 13454 14098 13488
rect 14040 13420 14052 13454
rect 14086 13420 14098 13454
rect 14040 13386 14098 13420
rect 14040 13352 14052 13386
rect 14086 13352 14098 13386
rect 14040 13318 14098 13352
rect 14040 13284 14052 13318
rect 14086 13284 14098 13318
rect 14040 13250 14098 13284
rect 14040 13216 14052 13250
rect 14086 13216 14098 13250
rect 14040 13182 14098 13216
rect 14040 13148 14052 13182
rect 14086 13148 14098 13182
rect 14040 13114 14098 13148
rect 14040 13080 14052 13114
rect 14086 13080 14098 13114
rect 14040 13046 14098 13080
rect 14040 13012 14052 13046
rect 14086 13012 14098 13046
rect 14040 12978 14098 13012
rect 14040 12944 14052 12978
rect 14086 12944 14098 12978
rect 14040 12910 14098 12944
rect 14040 12876 14052 12910
rect 14086 12876 14098 12910
rect 14040 12842 14098 12876
rect 14040 12808 14052 12842
rect 14086 12808 14098 12842
rect 14040 12774 14098 12808
rect 14040 12740 14052 12774
rect 14086 12740 14098 12774
rect 14040 12706 14098 12740
rect 14040 12672 14052 12706
rect 14086 12672 14098 12706
rect 14040 12638 14098 12672
rect 14040 12604 14052 12638
rect 14086 12604 14098 12638
rect 14040 12570 14098 12604
rect 14040 12536 14052 12570
rect 14086 12536 14098 12570
rect 14040 12502 14098 12536
rect 14040 12468 14052 12502
rect 14086 12468 14098 12502
rect 14040 12434 14098 12468
rect 14040 12400 14052 12434
rect 14086 12400 14098 12434
rect 14040 12366 14098 12400
rect 14040 12332 14052 12366
rect 14086 12332 14098 12366
rect 14040 12298 14098 12332
rect 14040 12264 14052 12298
rect 14086 12264 14098 12298
rect 14040 12230 14098 12264
rect 14040 12196 14052 12230
rect 14086 12196 14098 12230
rect 14040 12162 14098 12196
rect 14040 12128 14052 12162
rect 14086 12128 14098 12162
rect 14040 12094 14098 12128
rect 14040 12060 14052 12094
rect 14086 12060 14098 12094
rect 14040 12026 14098 12060
rect 14040 11992 14052 12026
rect 14086 11992 14098 12026
rect 14040 11958 14098 11992
rect 14040 11924 14052 11958
rect 14086 11924 14098 11958
rect 14040 11890 14098 11924
rect 14040 11856 14052 11890
rect 14086 11856 14098 11890
rect 14040 11822 14098 11856
rect 14040 11788 14052 11822
rect 14086 11788 14098 11822
rect 14040 11767 14098 11788
rect 15098 14746 15156 14767
rect 15098 14712 15110 14746
rect 15144 14712 15156 14746
rect 15098 14678 15156 14712
rect 15098 14644 15110 14678
rect 15144 14644 15156 14678
rect 15098 14610 15156 14644
rect 15098 14576 15110 14610
rect 15144 14576 15156 14610
rect 15098 14542 15156 14576
rect 15098 14508 15110 14542
rect 15144 14508 15156 14542
rect 15098 14474 15156 14508
rect 15098 14440 15110 14474
rect 15144 14440 15156 14474
rect 15098 14406 15156 14440
rect 15098 14372 15110 14406
rect 15144 14372 15156 14406
rect 15098 14338 15156 14372
rect 15098 14304 15110 14338
rect 15144 14304 15156 14338
rect 15098 14270 15156 14304
rect 15098 14236 15110 14270
rect 15144 14236 15156 14270
rect 15098 14202 15156 14236
rect 15098 14168 15110 14202
rect 15144 14168 15156 14202
rect 15098 14134 15156 14168
rect 15098 14100 15110 14134
rect 15144 14100 15156 14134
rect 15098 14066 15156 14100
rect 15098 14032 15110 14066
rect 15144 14032 15156 14066
rect 15098 13998 15156 14032
rect 15098 13964 15110 13998
rect 15144 13964 15156 13998
rect 15098 13930 15156 13964
rect 15098 13896 15110 13930
rect 15144 13896 15156 13930
rect 15098 13862 15156 13896
rect 15098 13828 15110 13862
rect 15144 13828 15156 13862
rect 15098 13794 15156 13828
rect 15098 13760 15110 13794
rect 15144 13760 15156 13794
rect 15098 13726 15156 13760
rect 15098 13692 15110 13726
rect 15144 13692 15156 13726
rect 15098 13658 15156 13692
rect 15098 13624 15110 13658
rect 15144 13624 15156 13658
rect 15098 13590 15156 13624
rect 15098 13556 15110 13590
rect 15144 13556 15156 13590
rect 15098 13522 15156 13556
rect 15098 13488 15110 13522
rect 15144 13488 15156 13522
rect 15098 13454 15156 13488
rect 15098 13420 15110 13454
rect 15144 13420 15156 13454
rect 15098 13386 15156 13420
rect 15098 13352 15110 13386
rect 15144 13352 15156 13386
rect 15098 13318 15156 13352
rect 15098 13284 15110 13318
rect 15144 13284 15156 13318
rect 15098 13250 15156 13284
rect 15098 13216 15110 13250
rect 15144 13216 15156 13250
rect 15098 13182 15156 13216
rect 15098 13148 15110 13182
rect 15144 13148 15156 13182
rect 15098 13114 15156 13148
rect 15098 13080 15110 13114
rect 15144 13080 15156 13114
rect 15098 13046 15156 13080
rect 15098 13012 15110 13046
rect 15144 13012 15156 13046
rect 15098 12978 15156 13012
rect 15098 12944 15110 12978
rect 15144 12944 15156 12978
rect 15098 12910 15156 12944
rect 15098 12876 15110 12910
rect 15144 12876 15156 12910
rect 15098 12842 15156 12876
rect 15098 12808 15110 12842
rect 15144 12808 15156 12842
rect 15098 12774 15156 12808
rect 15098 12740 15110 12774
rect 15144 12740 15156 12774
rect 15098 12706 15156 12740
rect 15098 12672 15110 12706
rect 15144 12672 15156 12706
rect 15098 12638 15156 12672
rect 15098 12604 15110 12638
rect 15144 12604 15156 12638
rect 15098 12570 15156 12604
rect 15098 12536 15110 12570
rect 15144 12536 15156 12570
rect 15098 12502 15156 12536
rect 15098 12468 15110 12502
rect 15144 12468 15156 12502
rect 15098 12434 15156 12468
rect 15098 12400 15110 12434
rect 15144 12400 15156 12434
rect 15098 12366 15156 12400
rect 15098 12332 15110 12366
rect 15144 12332 15156 12366
rect 15098 12298 15156 12332
rect 15098 12264 15110 12298
rect 15144 12264 15156 12298
rect 15098 12230 15156 12264
rect 15098 12196 15110 12230
rect 15144 12196 15156 12230
rect 15098 12162 15156 12196
rect 15098 12128 15110 12162
rect 15144 12128 15156 12162
rect 15098 12094 15156 12128
rect 15098 12060 15110 12094
rect 15144 12060 15156 12094
rect 15098 12026 15156 12060
rect 15098 11992 15110 12026
rect 15144 11992 15156 12026
rect 15098 11958 15156 11992
rect 15098 11924 15110 11958
rect 15144 11924 15156 11958
rect 15098 11890 15156 11924
rect 15098 11856 15110 11890
rect 15144 11856 15156 11890
rect 15098 11822 15156 11856
rect 15098 11788 15110 11822
rect 15144 11788 15156 11822
rect 15098 11767 15156 11788
rect 15552 14746 15610 14767
rect 15552 14712 15564 14746
rect 15598 14712 15610 14746
rect 15552 14678 15610 14712
rect 15552 14644 15564 14678
rect 15598 14644 15610 14678
rect 15552 14610 15610 14644
rect 15552 14576 15564 14610
rect 15598 14576 15610 14610
rect 15552 14542 15610 14576
rect 15552 14508 15564 14542
rect 15598 14508 15610 14542
rect 15552 14474 15610 14508
rect 15552 14440 15564 14474
rect 15598 14440 15610 14474
rect 15552 14406 15610 14440
rect 15552 14372 15564 14406
rect 15598 14372 15610 14406
rect 15552 14338 15610 14372
rect 15552 14304 15564 14338
rect 15598 14304 15610 14338
rect 15552 14270 15610 14304
rect 15552 14236 15564 14270
rect 15598 14236 15610 14270
rect 15552 14202 15610 14236
rect 15552 14168 15564 14202
rect 15598 14168 15610 14202
rect 15552 14134 15610 14168
rect 15552 14100 15564 14134
rect 15598 14100 15610 14134
rect 15552 14066 15610 14100
rect 15552 14032 15564 14066
rect 15598 14032 15610 14066
rect 15552 13998 15610 14032
rect 15552 13964 15564 13998
rect 15598 13964 15610 13998
rect 15552 13930 15610 13964
rect 15552 13896 15564 13930
rect 15598 13896 15610 13930
rect 15552 13862 15610 13896
rect 15552 13828 15564 13862
rect 15598 13828 15610 13862
rect 15552 13794 15610 13828
rect 15552 13760 15564 13794
rect 15598 13760 15610 13794
rect 15552 13726 15610 13760
rect 15552 13692 15564 13726
rect 15598 13692 15610 13726
rect 15552 13658 15610 13692
rect 15552 13624 15564 13658
rect 15598 13624 15610 13658
rect 15552 13590 15610 13624
rect 15552 13556 15564 13590
rect 15598 13556 15610 13590
rect 15552 13522 15610 13556
rect 15552 13488 15564 13522
rect 15598 13488 15610 13522
rect 15552 13454 15610 13488
rect 15552 13420 15564 13454
rect 15598 13420 15610 13454
rect 15552 13386 15610 13420
rect 15552 13352 15564 13386
rect 15598 13352 15610 13386
rect 15552 13318 15610 13352
rect 15552 13284 15564 13318
rect 15598 13284 15610 13318
rect 15552 13250 15610 13284
rect 15552 13216 15564 13250
rect 15598 13216 15610 13250
rect 15552 13182 15610 13216
rect 15552 13148 15564 13182
rect 15598 13148 15610 13182
rect 15552 13114 15610 13148
rect 15552 13080 15564 13114
rect 15598 13080 15610 13114
rect 15552 13046 15610 13080
rect 15552 13012 15564 13046
rect 15598 13012 15610 13046
rect 15552 12978 15610 13012
rect 15552 12944 15564 12978
rect 15598 12944 15610 12978
rect 15552 12910 15610 12944
rect 15552 12876 15564 12910
rect 15598 12876 15610 12910
rect 15552 12842 15610 12876
rect 15552 12808 15564 12842
rect 15598 12808 15610 12842
rect 15552 12774 15610 12808
rect 15552 12740 15564 12774
rect 15598 12740 15610 12774
rect 15552 12706 15610 12740
rect 15552 12672 15564 12706
rect 15598 12672 15610 12706
rect 15552 12638 15610 12672
rect 15552 12604 15564 12638
rect 15598 12604 15610 12638
rect 15552 12570 15610 12604
rect 15552 12536 15564 12570
rect 15598 12536 15610 12570
rect 15552 12502 15610 12536
rect 15552 12468 15564 12502
rect 15598 12468 15610 12502
rect 15552 12434 15610 12468
rect 15552 12400 15564 12434
rect 15598 12400 15610 12434
rect 15552 12366 15610 12400
rect 15552 12332 15564 12366
rect 15598 12332 15610 12366
rect 15552 12298 15610 12332
rect 15552 12264 15564 12298
rect 15598 12264 15610 12298
rect 15552 12230 15610 12264
rect 15552 12196 15564 12230
rect 15598 12196 15610 12230
rect 15552 12162 15610 12196
rect 15552 12128 15564 12162
rect 15598 12128 15610 12162
rect 15552 12094 15610 12128
rect 15552 12060 15564 12094
rect 15598 12060 15610 12094
rect 15552 12026 15610 12060
rect 15552 11992 15564 12026
rect 15598 11992 15610 12026
rect 15552 11958 15610 11992
rect 15552 11924 15564 11958
rect 15598 11924 15610 11958
rect 15552 11890 15610 11924
rect 15552 11856 15564 11890
rect 15598 11856 15610 11890
rect 15552 11822 15610 11856
rect 15552 11788 15564 11822
rect 15598 11788 15610 11822
rect 15552 11767 15610 11788
rect 16610 14746 16668 14767
rect 16610 14712 16622 14746
rect 16656 14712 16668 14746
rect 16610 14678 16668 14712
rect 16610 14644 16622 14678
rect 16656 14644 16668 14678
rect 16610 14610 16668 14644
rect 16610 14576 16622 14610
rect 16656 14576 16668 14610
rect 16610 14542 16668 14576
rect 16610 14508 16622 14542
rect 16656 14508 16668 14542
rect 16610 14474 16668 14508
rect 16610 14440 16622 14474
rect 16656 14440 16668 14474
rect 16610 14406 16668 14440
rect 16610 14372 16622 14406
rect 16656 14372 16668 14406
rect 16610 14338 16668 14372
rect 16610 14304 16622 14338
rect 16656 14304 16668 14338
rect 16610 14270 16668 14304
rect 16610 14236 16622 14270
rect 16656 14236 16668 14270
rect 16610 14202 16668 14236
rect 16610 14168 16622 14202
rect 16656 14168 16668 14202
rect 16610 14134 16668 14168
rect 16610 14100 16622 14134
rect 16656 14100 16668 14134
rect 16610 14066 16668 14100
rect 16610 14032 16622 14066
rect 16656 14032 16668 14066
rect 16610 13998 16668 14032
rect 16610 13964 16622 13998
rect 16656 13964 16668 13998
rect 16610 13930 16668 13964
rect 16610 13896 16622 13930
rect 16656 13896 16668 13930
rect 16610 13862 16668 13896
rect 16610 13828 16622 13862
rect 16656 13828 16668 13862
rect 16610 13794 16668 13828
rect 16610 13760 16622 13794
rect 16656 13760 16668 13794
rect 16610 13726 16668 13760
rect 16610 13692 16622 13726
rect 16656 13692 16668 13726
rect 16610 13658 16668 13692
rect 16610 13624 16622 13658
rect 16656 13624 16668 13658
rect 16610 13590 16668 13624
rect 16610 13556 16622 13590
rect 16656 13556 16668 13590
rect 16610 13522 16668 13556
rect 16610 13488 16622 13522
rect 16656 13488 16668 13522
rect 16610 13454 16668 13488
rect 16610 13420 16622 13454
rect 16656 13420 16668 13454
rect 16610 13386 16668 13420
rect 16610 13352 16622 13386
rect 16656 13352 16668 13386
rect 16610 13318 16668 13352
rect 16610 13284 16622 13318
rect 16656 13284 16668 13318
rect 16610 13250 16668 13284
rect 16610 13216 16622 13250
rect 16656 13216 16668 13250
rect 16610 13182 16668 13216
rect 16610 13148 16622 13182
rect 16656 13148 16668 13182
rect 16610 13114 16668 13148
rect 16610 13080 16622 13114
rect 16656 13080 16668 13114
rect 16610 13046 16668 13080
rect 16610 13012 16622 13046
rect 16656 13012 16668 13046
rect 16610 12978 16668 13012
rect 16610 12944 16622 12978
rect 16656 12944 16668 12978
rect 16610 12910 16668 12944
rect 16610 12876 16622 12910
rect 16656 12876 16668 12910
rect 16610 12842 16668 12876
rect 16610 12808 16622 12842
rect 16656 12808 16668 12842
rect 16610 12774 16668 12808
rect 16610 12740 16622 12774
rect 16656 12740 16668 12774
rect 16610 12706 16668 12740
rect 16610 12672 16622 12706
rect 16656 12672 16668 12706
rect 16610 12638 16668 12672
rect 16610 12604 16622 12638
rect 16656 12604 16668 12638
rect 16610 12570 16668 12604
rect 16610 12536 16622 12570
rect 16656 12536 16668 12570
rect 16610 12502 16668 12536
rect 16610 12468 16622 12502
rect 16656 12468 16668 12502
rect 16610 12434 16668 12468
rect 16610 12400 16622 12434
rect 16656 12400 16668 12434
rect 16610 12366 16668 12400
rect 16610 12332 16622 12366
rect 16656 12332 16668 12366
rect 16610 12298 16668 12332
rect 16610 12264 16622 12298
rect 16656 12264 16668 12298
rect 16610 12230 16668 12264
rect 16610 12196 16622 12230
rect 16656 12196 16668 12230
rect 16610 12162 16668 12196
rect 16610 12128 16622 12162
rect 16656 12128 16668 12162
rect 16610 12094 16668 12128
rect 16610 12060 16622 12094
rect 16656 12060 16668 12094
rect 16610 12026 16668 12060
rect 16610 11992 16622 12026
rect 16656 11992 16668 12026
rect 16610 11958 16668 11992
rect 16610 11924 16622 11958
rect 16656 11924 16668 11958
rect 16610 11890 16668 11924
rect 16610 11856 16622 11890
rect 16656 11856 16668 11890
rect 16610 11822 16668 11856
rect 16610 11788 16622 11822
rect 16656 11788 16668 11822
rect 16610 11767 16668 11788
rect 17062 14756 17120 14777
rect 17062 14722 17074 14756
rect 17108 14722 17120 14756
rect 17062 14688 17120 14722
rect 17062 14654 17074 14688
rect 17108 14654 17120 14688
rect 17062 14620 17120 14654
rect 17062 14586 17074 14620
rect 17108 14586 17120 14620
rect 17062 14552 17120 14586
rect 17062 14518 17074 14552
rect 17108 14518 17120 14552
rect 17062 14484 17120 14518
rect 17062 14450 17074 14484
rect 17108 14450 17120 14484
rect 17062 14416 17120 14450
rect 17062 14382 17074 14416
rect 17108 14382 17120 14416
rect 17062 14348 17120 14382
rect 17062 14314 17074 14348
rect 17108 14314 17120 14348
rect 17062 14280 17120 14314
rect 17062 14246 17074 14280
rect 17108 14246 17120 14280
rect 17062 14212 17120 14246
rect 17062 14178 17074 14212
rect 17108 14178 17120 14212
rect 17062 14144 17120 14178
rect 17062 14110 17074 14144
rect 17108 14110 17120 14144
rect 17062 14076 17120 14110
rect 17062 14042 17074 14076
rect 17108 14042 17120 14076
rect 17062 14008 17120 14042
rect 17062 13974 17074 14008
rect 17108 13974 17120 14008
rect 17062 13940 17120 13974
rect 17062 13906 17074 13940
rect 17108 13906 17120 13940
rect 17062 13872 17120 13906
rect 17062 13838 17074 13872
rect 17108 13838 17120 13872
rect 17062 13804 17120 13838
rect 17062 13770 17074 13804
rect 17108 13770 17120 13804
rect 17062 13736 17120 13770
rect 17062 13702 17074 13736
rect 17108 13702 17120 13736
rect 17062 13668 17120 13702
rect 17062 13634 17074 13668
rect 17108 13634 17120 13668
rect 17062 13600 17120 13634
rect 17062 13566 17074 13600
rect 17108 13566 17120 13600
rect 17062 13532 17120 13566
rect 17062 13498 17074 13532
rect 17108 13498 17120 13532
rect 17062 13464 17120 13498
rect 17062 13430 17074 13464
rect 17108 13430 17120 13464
rect 17062 13396 17120 13430
rect 17062 13362 17074 13396
rect 17108 13362 17120 13396
rect 17062 13328 17120 13362
rect 17062 13294 17074 13328
rect 17108 13294 17120 13328
rect 17062 13260 17120 13294
rect 17062 13226 17074 13260
rect 17108 13226 17120 13260
rect 17062 13192 17120 13226
rect 17062 13158 17074 13192
rect 17108 13158 17120 13192
rect 17062 13124 17120 13158
rect 17062 13090 17074 13124
rect 17108 13090 17120 13124
rect 17062 13056 17120 13090
rect 17062 13022 17074 13056
rect 17108 13022 17120 13056
rect 17062 12988 17120 13022
rect 17062 12954 17074 12988
rect 17108 12954 17120 12988
rect 17062 12920 17120 12954
rect 17062 12886 17074 12920
rect 17108 12886 17120 12920
rect 17062 12852 17120 12886
rect 17062 12818 17074 12852
rect 17108 12818 17120 12852
rect 17062 12784 17120 12818
rect 17062 12750 17074 12784
rect 17108 12750 17120 12784
rect 17062 12716 17120 12750
rect 17062 12682 17074 12716
rect 17108 12682 17120 12716
rect 17062 12648 17120 12682
rect 17062 12614 17074 12648
rect 17108 12614 17120 12648
rect 17062 12580 17120 12614
rect 17062 12546 17074 12580
rect 17108 12546 17120 12580
rect 17062 12512 17120 12546
rect 17062 12478 17074 12512
rect 17108 12478 17120 12512
rect 17062 12444 17120 12478
rect 17062 12410 17074 12444
rect 17108 12410 17120 12444
rect 17062 12376 17120 12410
rect 17062 12342 17074 12376
rect 17108 12342 17120 12376
rect 17062 12308 17120 12342
rect 17062 12274 17074 12308
rect 17108 12274 17120 12308
rect 17062 12240 17120 12274
rect 17062 12206 17074 12240
rect 17108 12206 17120 12240
rect 17062 12172 17120 12206
rect 17062 12138 17074 12172
rect 17108 12138 17120 12172
rect 17062 12104 17120 12138
rect 17062 12070 17074 12104
rect 17108 12070 17120 12104
rect 17062 12036 17120 12070
rect 17062 12002 17074 12036
rect 17108 12002 17120 12036
rect 17062 11968 17120 12002
rect 17062 11934 17074 11968
rect 17108 11934 17120 11968
rect 17062 11900 17120 11934
rect 17062 11866 17074 11900
rect 17108 11866 17120 11900
rect 17062 11832 17120 11866
rect 17062 11798 17074 11832
rect 17108 11798 17120 11832
rect 17062 11777 17120 11798
rect 18120 14756 18178 14777
rect 18120 14722 18132 14756
rect 18166 14722 18178 14756
rect 18120 14688 18178 14722
rect 18120 14654 18132 14688
rect 18166 14654 18178 14688
rect 18120 14620 18178 14654
rect 18120 14586 18132 14620
rect 18166 14586 18178 14620
rect 18120 14552 18178 14586
rect 18120 14518 18132 14552
rect 18166 14518 18178 14552
rect 18120 14484 18178 14518
rect 18120 14450 18132 14484
rect 18166 14450 18178 14484
rect 18120 14416 18178 14450
rect 18120 14382 18132 14416
rect 18166 14382 18178 14416
rect 18120 14348 18178 14382
rect 18120 14314 18132 14348
rect 18166 14314 18178 14348
rect 18120 14280 18178 14314
rect 18120 14246 18132 14280
rect 18166 14246 18178 14280
rect 18120 14212 18178 14246
rect 18120 14178 18132 14212
rect 18166 14178 18178 14212
rect 18120 14144 18178 14178
rect 18120 14110 18132 14144
rect 18166 14110 18178 14144
rect 18120 14076 18178 14110
rect 18120 14042 18132 14076
rect 18166 14042 18178 14076
rect 18120 14008 18178 14042
rect 18120 13974 18132 14008
rect 18166 13974 18178 14008
rect 18120 13940 18178 13974
rect 18120 13906 18132 13940
rect 18166 13906 18178 13940
rect 18120 13872 18178 13906
rect 18120 13838 18132 13872
rect 18166 13838 18178 13872
rect 18120 13804 18178 13838
rect 18120 13770 18132 13804
rect 18166 13770 18178 13804
rect 18120 13736 18178 13770
rect 18120 13702 18132 13736
rect 18166 13702 18178 13736
rect 18120 13668 18178 13702
rect 18120 13634 18132 13668
rect 18166 13634 18178 13668
rect 18120 13600 18178 13634
rect 18120 13566 18132 13600
rect 18166 13566 18178 13600
rect 18120 13532 18178 13566
rect 18120 13498 18132 13532
rect 18166 13498 18178 13532
rect 18120 13464 18178 13498
rect 18120 13430 18132 13464
rect 18166 13430 18178 13464
rect 18120 13396 18178 13430
rect 18120 13362 18132 13396
rect 18166 13362 18178 13396
rect 18120 13328 18178 13362
rect 18120 13294 18132 13328
rect 18166 13294 18178 13328
rect 18120 13260 18178 13294
rect 18120 13226 18132 13260
rect 18166 13226 18178 13260
rect 18120 13192 18178 13226
rect 18120 13158 18132 13192
rect 18166 13158 18178 13192
rect 18120 13124 18178 13158
rect 18120 13090 18132 13124
rect 18166 13090 18178 13124
rect 18120 13056 18178 13090
rect 18120 13022 18132 13056
rect 18166 13022 18178 13056
rect 18120 12988 18178 13022
rect 18120 12954 18132 12988
rect 18166 12954 18178 12988
rect 18120 12920 18178 12954
rect 18120 12886 18132 12920
rect 18166 12886 18178 12920
rect 18120 12852 18178 12886
rect 18120 12818 18132 12852
rect 18166 12818 18178 12852
rect 18120 12784 18178 12818
rect 18120 12750 18132 12784
rect 18166 12750 18178 12784
rect 18120 12716 18178 12750
rect 18120 12682 18132 12716
rect 18166 12682 18178 12716
rect 18120 12648 18178 12682
rect 18120 12614 18132 12648
rect 18166 12614 18178 12648
rect 18120 12580 18178 12614
rect 18120 12546 18132 12580
rect 18166 12546 18178 12580
rect 18120 12512 18178 12546
rect 18120 12478 18132 12512
rect 18166 12478 18178 12512
rect 18120 12444 18178 12478
rect 18120 12410 18132 12444
rect 18166 12410 18178 12444
rect 18120 12376 18178 12410
rect 18120 12342 18132 12376
rect 18166 12342 18178 12376
rect 18120 12308 18178 12342
rect 18120 12274 18132 12308
rect 18166 12274 18178 12308
rect 18120 12240 18178 12274
rect 18120 12206 18132 12240
rect 18166 12206 18178 12240
rect 18120 12172 18178 12206
rect 18120 12138 18132 12172
rect 18166 12138 18178 12172
rect 18120 12104 18178 12138
rect 18120 12070 18132 12104
rect 18166 12070 18178 12104
rect 18120 12036 18178 12070
rect 18120 12002 18132 12036
rect 18166 12002 18178 12036
rect 18120 11968 18178 12002
rect 18120 11934 18132 11968
rect 18166 11934 18178 11968
rect 18120 11900 18178 11934
rect 18120 11866 18132 11900
rect 18166 11866 18178 11900
rect 18120 11832 18178 11866
rect 18120 11798 18132 11832
rect 18166 11798 18178 11832
rect 18120 11777 18178 11798
rect 18526 14740 18584 14761
rect 18526 14706 18538 14740
rect 18572 14706 18584 14740
rect 18526 14672 18584 14706
rect 18526 14638 18538 14672
rect 18572 14638 18584 14672
rect 18526 14604 18584 14638
rect 18526 14570 18538 14604
rect 18572 14570 18584 14604
rect 18526 14536 18584 14570
rect 18526 14502 18538 14536
rect 18572 14502 18584 14536
rect 18526 14468 18584 14502
rect 18526 14434 18538 14468
rect 18572 14434 18584 14468
rect 18526 14400 18584 14434
rect 18526 14366 18538 14400
rect 18572 14366 18584 14400
rect 18526 14332 18584 14366
rect 18526 14298 18538 14332
rect 18572 14298 18584 14332
rect 18526 14264 18584 14298
rect 18526 14230 18538 14264
rect 18572 14230 18584 14264
rect 18526 14196 18584 14230
rect 18526 14162 18538 14196
rect 18572 14162 18584 14196
rect 18526 14128 18584 14162
rect 18526 14094 18538 14128
rect 18572 14094 18584 14128
rect 18526 14060 18584 14094
rect 18526 14026 18538 14060
rect 18572 14026 18584 14060
rect 18526 13992 18584 14026
rect 18526 13958 18538 13992
rect 18572 13958 18584 13992
rect 18526 13924 18584 13958
rect 18526 13890 18538 13924
rect 18572 13890 18584 13924
rect 18526 13856 18584 13890
rect 18526 13822 18538 13856
rect 18572 13822 18584 13856
rect 18526 13788 18584 13822
rect 18526 13754 18538 13788
rect 18572 13754 18584 13788
rect 18526 13720 18584 13754
rect 18526 13686 18538 13720
rect 18572 13686 18584 13720
rect 18526 13652 18584 13686
rect 18526 13618 18538 13652
rect 18572 13618 18584 13652
rect 18526 13584 18584 13618
rect 18526 13550 18538 13584
rect 18572 13550 18584 13584
rect 18526 13516 18584 13550
rect 18526 13482 18538 13516
rect 18572 13482 18584 13516
rect 18526 13448 18584 13482
rect 18526 13414 18538 13448
rect 18572 13414 18584 13448
rect 18526 13380 18584 13414
rect 18526 13346 18538 13380
rect 18572 13346 18584 13380
rect 18526 13312 18584 13346
rect 18526 13278 18538 13312
rect 18572 13278 18584 13312
rect 18526 13244 18584 13278
rect 18526 13210 18538 13244
rect 18572 13210 18584 13244
rect 18526 13176 18584 13210
rect 18526 13142 18538 13176
rect 18572 13142 18584 13176
rect 18526 13108 18584 13142
rect 18526 13074 18538 13108
rect 18572 13074 18584 13108
rect 18526 13040 18584 13074
rect 18526 13006 18538 13040
rect 18572 13006 18584 13040
rect 18526 12972 18584 13006
rect 18526 12938 18538 12972
rect 18572 12938 18584 12972
rect 18526 12904 18584 12938
rect 18526 12870 18538 12904
rect 18572 12870 18584 12904
rect 18526 12836 18584 12870
rect 18526 12802 18538 12836
rect 18572 12802 18584 12836
rect 18526 12768 18584 12802
rect 18526 12734 18538 12768
rect 18572 12734 18584 12768
rect 18526 12700 18584 12734
rect 18526 12666 18538 12700
rect 18572 12666 18584 12700
rect 18526 12632 18584 12666
rect 18526 12598 18538 12632
rect 18572 12598 18584 12632
rect 18526 12564 18584 12598
rect 18526 12530 18538 12564
rect 18572 12530 18584 12564
rect 18526 12496 18584 12530
rect 18526 12462 18538 12496
rect 18572 12462 18584 12496
rect 18526 12428 18584 12462
rect 18526 12394 18538 12428
rect 18572 12394 18584 12428
rect 18526 12360 18584 12394
rect 18526 12326 18538 12360
rect 18572 12326 18584 12360
rect 18526 12292 18584 12326
rect 18526 12258 18538 12292
rect 18572 12258 18584 12292
rect 18526 12224 18584 12258
rect 18526 12190 18538 12224
rect 18572 12190 18584 12224
rect 18526 12156 18584 12190
rect 18526 12122 18538 12156
rect 18572 12122 18584 12156
rect 18526 12088 18584 12122
rect 18526 12054 18538 12088
rect 18572 12054 18584 12088
rect 18526 12020 18584 12054
rect 18526 11986 18538 12020
rect 18572 11986 18584 12020
rect 18526 11952 18584 11986
rect 18526 11918 18538 11952
rect 18572 11918 18584 11952
rect 18526 11884 18584 11918
rect 18526 11850 18538 11884
rect 18572 11850 18584 11884
rect 18526 11816 18584 11850
rect 18526 11782 18538 11816
rect 18572 11782 18584 11816
rect 18526 11761 18584 11782
rect 19584 14740 19642 14761
rect 19584 14706 19596 14740
rect 19630 14706 19642 14740
rect 19584 14672 19642 14706
rect 19584 14638 19596 14672
rect 19630 14638 19642 14672
rect 19584 14604 19642 14638
rect 19584 14570 19596 14604
rect 19630 14570 19642 14604
rect 19584 14536 19642 14570
rect 19584 14502 19596 14536
rect 19630 14502 19642 14536
rect 19584 14468 19642 14502
rect 19584 14434 19596 14468
rect 19630 14434 19642 14468
rect 19584 14400 19642 14434
rect 19584 14366 19596 14400
rect 19630 14366 19642 14400
rect 19584 14332 19642 14366
rect 19584 14298 19596 14332
rect 19630 14298 19642 14332
rect 19584 14264 19642 14298
rect 19584 14230 19596 14264
rect 19630 14230 19642 14264
rect 19584 14196 19642 14230
rect 19584 14162 19596 14196
rect 19630 14162 19642 14196
rect 19584 14128 19642 14162
rect 19584 14094 19596 14128
rect 19630 14094 19642 14128
rect 19584 14060 19642 14094
rect 19584 14026 19596 14060
rect 19630 14026 19642 14060
rect 19584 13992 19642 14026
rect 19584 13958 19596 13992
rect 19630 13958 19642 13992
rect 19584 13924 19642 13958
rect 19584 13890 19596 13924
rect 19630 13890 19642 13924
rect 19584 13856 19642 13890
rect 19584 13822 19596 13856
rect 19630 13822 19642 13856
rect 19584 13788 19642 13822
rect 19584 13754 19596 13788
rect 19630 13754 19642 13788
rect 19584 13720 19642 13754
rect 19584 13686 19596 13720
rect 19630 13686 19642 13720
rect 19584 13652 19642 13686
rect 19584 13618 19596 13652
rect 19630 13618 19642 13652
rect 19584 13584 19642 13618
rect 19584 13550 19596 13584
rect 19630 13550 19642 13584
rect 19584 13516 19642 13550
rect 19584 13482 19596 13516
rect 19630 13482 19642 13516
rect 19584 13448 19642 13482
rect 19584 13414 19596 13448
rect 19630 13414 19642 13448
rect 19584 13380 19642 13414
rect 19584 13346 19596 13380
rect 19630 13346 19642 13380
rect 19584 13312 19642 13346
rect 19584 13278 19596 13312
rect 19630 13278 19642 13312
rect 19584 13244 19642 13278
rect 19584 13210 19596 13244
rect 19630 13210 19642 13244
rect 19584 13176 19642 13210
rect 19584 13142 19596 13176
rect 19630 13142 19642 13176
rect 19584 13108 19642 13142
rect 19584 13074 19596 13108
rect 19630 13074 19642 13108
rect 19584 13040 19642 13074
rect 19584 13006 19596 13040
rect 19630 13006 19642 13040
rect 19584 12972 19642 13006
rect 19584 12938 19596 12972
rect 19630 12938 19642 12972
rect 19584 12904 19642 12938
rect 19584 12870 19596 12904
rect 19630 12870 19642 12904
rect 19584 12836 19642 12870
rect 19584 12802 19596 12836
rect 19630 12802 19642 12836
rect 19584 12768 19642 12802
rect 19584 12734 19596 12768
rect 19630 12734 19642 12768
rect 19584 12700 19642 12734
rect 19584 12666 19596 12700
rect 19630 12666 19642 12700
rect 19584 12632 19642 12666
rect 19584 12598 19596 12632
rect 19630 12598 19642 12632
rect 19584 12564 19642 12598
rect 19584 12530 19596 12564
rect 19630 12530 19642 12564
rect 19584 12496 19642 12530
rect 19584 12462 19596 12496
rect 19630 12462 19642 12496
rect 19584 12428 19642 12462
rect 19584 12394 19596 12428
rect 19630 12394 19642 12428
rect 19584 12360 19642 12394
rect 19584 12326 19596 12360
rect 19630 12326 19642 12360
rect 19584 12292 19642 12326
rect 19584 12258 19596 12292
rect 19630 12258 19642 12292
rect 19584 12224 19642 12258
rect 19584 12190 19596 12224
rect 19630 12190 19642 12224
rect 19584 12156 19642 12190
rect 19584 12122 19596 12156
rect 19630 12122 19642 12156
rect 19584 12088 19642 12122
rect 19584 12054 19596 12088
rect 19630 12054 19642 12088
rect 19584 12020 19642 12054
rect 19584 11986 19596 12020
rect 19630 11986 19642 12020
rect 19584 11952 19642 11986
rect 19584 11918 19596 11952
rect 19630 11918 19642 11952
rect 19584 11884 19642 11918
rect 19584 11850 19596 11884
rect 19630 11850 19642 11884
rect 19584 11816 19642 11850
rect 19584 11782 19596 11816
rect 19630 11782 19642 11816
rect 19584 11761 19642 11782
rect 14942 11226 15000 11247
rect 14942 11192 14954 11226
rect 14988 11192 15000 11226
rect 14942 11158 15000 11192
rect 14942 11124 14954 11158
rect 14988 11124 15000 11158
rect 14942 11090 15000 11124
rect 14942 11056 14954 11090
rect 14988 11056 15000 11090
rect 14942 11022 15000 11056
rect 14942 10988 14954 11022
rect 14988 10988 15000 11022
rect 14942 10954 15000 10988
rect 14942 10920 14954 10954
rect 14988 10920 15000 10954
rect 14942 10886 15000 10920
rect 14942 10852 14954 10886
rect 14988 10852 15000 10886
rect 14942 10818 15000 10852
rect 14942 10784 14954 10818
rect 14988 10784 15000 10818
rect 14942 10750 15000 10784
rect 14942 10716 14954 10750
rect 14988 10716 15000 10750
rect 14942 10682 15000 10716
rect 14942 10648 14954 10682
rect 14988 10648 15000 10682
rect 14942 10614 15000 10648
rect 14942 10580 14954 10614
rect 14988 10580 15000 10614
rect 14942 10546 15000 10580
rect 14942 10512 14954 10546
rect 14988 10512 15000 10546
rect 14942 10478 15000 10512
rect 14942 10444 14954 10478
rect 14988 10444 15000 10478
rect 14942 10410 15000 10444
rect 14942 10376 14954 10410
rect 14988 10376 15000 10410
rect 14942 10342 15000 10376
rect 14942 10308 14954 10342
rect 14988 10308 15000 10342
rect 14942 10274 15000 10308
rect 14942 10240 14954 10274
rect 14988 10240 15000 10274
rect 14942 10206 15000 10240
rect 14942 10172 14954 10206
rect 14988 10172 15000 10206
rect 14942 10138 15000 10172
rect 14942 10104 14954 10138
rect 14988 10104 15000 10138
rect 14942 10070 15000 10104
rect 14942 10036 14954 10070
rect 14988 10036 15000 10070
rect 14942 10002 15000 10036
rect 14942 9968 14954 10002
rect 14988 9968 15000 10002
rect 14942 9934 15000 9968
rect 14942 9900 14954 9934
rect 14988 9900 15000 9934
rect 14942 9866 15000 9900
rect 14942 9832 14954 9866
rect 14988 9832 15000 9866
rect 14942 9798 15000 9832
rect 14942 9764 14954 9798
rect 14988 9764 15000 9798
rect 14942 9730 15000 9764
rect 14942 9696 14954 9730
rect 14988 9696 15000 9730
rect 14942 9662 15000 9696
rect 14942 9628 14954 9662
rect 14988 9628 15000 9662
rect 14942 9594 15000 9628
rect 14942 9560 14954 9594
rect 14988 9560 15000 9594
rect 14942 9526 15000 9560
rect 14942 9492 14954 9526
rect 14988 9492 15000 9526
rect 14942 9458 15000 9492
rect 14942 9424 14954 9458
rect 14988 9424 15000 9458
rect 14942 9390 15000 9424
rect 14942 9356 14954 9390
rect 14988 9356 15000 9390
rect 14942 9322 15000 9356
rect 14942 9288 14954 9322
rect 14988 9288 15000 9322
rect 14942 9254 15000 9288
rect 14942 9220 14954 9254
rect 14988 9220 15000 9254
rect 14942 9186 15000 9220
rect 14942 9152 14954 9186
rect 14988 9152 15000 9186
rect 14942 9118 15000 9152
rect 14942 9084 14954 9118
rect 14988 9084 15000 9118
rect 14942 9050 15000 9084
rect 14942 9016 14954 9050
rect 14988 9016 15000 9050
rect 14942 8982 15000 9016
rect 14942 8948 14954 8982
rect 14988 8948 15000 8982
rect 14942 8914 15000 8948
rect 14942 8880 14954 8914
rect 14988 8880 15000 8914
rect 14942 8846 15000 8880
rect 14942 8812 14954 8846
rect 14988 8812 15000 8846
rect 14942 8778 15000 8812
rect 14942 8744 14954 8778
rect 14988 8744 15000 8778
rect 14942 8710 15000 8744
rect 14942 8676 14954 8710
rect 14988 8676 15000 8710
rect 14942 8642 15000 8676
rect 14942 8608 14954 8642
rect 14988 8608 15000 8642
rect 14942 8574 15000 8608
rect 14942 8540 14954 8574
rect 14988 8540 15000 8574
rect 14942 8506 15000 8540
rect 14942 8472 14954 8506
rect 14988 8472 15000 8506
rect 14942 8438 15000 8472
rect 14942 8404 14954 8438
rect 14988 8404 15000 8438
rect 14942 8370 15000 8404
rect 14942 8336 14954 8370
rect 14988 8336 15000 8370
rect 14942 8302 15000 8336
rect 14942 8268 14954 8302
rect 14988 8268 15000 8302
rect 14942 8247 15000 8268
rect 16000 11226 16058 11247
rect 16000 11192 16012 11226
rect 16046 11192 16058 11226
rect 16000 11158 16058 11192
rect 16000 11124 16012 11158
rect 16046 11124 16058 11158
rect 16000 11090 16058 11124
rect 16000 11056 16012 11090
rect 16046 11056 16058 11090
rect 16000 11022 16058 11056
rect 16000 10988 16012 11022
rect 16046 10988 16058 11022
rect 16000 10954 16058 10988
rect 16000 10920 16012 10954
rect 16046 10920 16058 10954
rect 16000 10886 16058 10920
rect 16000 10852 16012 10886
rect 16046 10852 16058 10886
rect 16000 10818 16058 10852
rect 16000 10784 16012 10818
rect 16046 10784 16058 10818
rect 16000 10750 16058 10784
rect 16000 10716 16012 10750
rect 16046 10716 16058 10750
rect 16000 10682 16058 10716
rect 16000 10648 16012 10682
rect 16046 10648 16058 10682
rect 16000 10614 16058 10648
rect 16000 10580 16012 10614
rect 16046 10580 16058 10614
rect 16000 10546 16058 10580
rect 16000 10512 16012 10546
rect 16046 10512 16058 10546
rect 16000 10478 16058 10512
rect 16000 10444 16012 10478
rect 16046 10444 16058 10478
rect 16000 10410 16058 10444
rect 16000 10376 16012 10410
rect 16046 10376 16058 10410
rect 16000 10342 16058 10376
rect 16000 10308 16012 10342
rect 16046 10308 16058 10342
rect 16000 10274 16058 10308
rect 16000 10240 16012 10274
rect 16046 10240 16058 10274
rect 16000 10206 16058 10240
rect 16000 10172 16012 10206
rect 16046 10172 16058 10206
rect 16000 10138 16058 10172
rect 16000 10104 16012 10138
rect 16046 10104 16058 10138
rect 16000 10070 16058 10104
rect 16000 10036 16012 10070
rect 16046 10036 16058 10070
rect 16000 10002 16058 10036
rect 16000 9968 16012 10002
rect 16046 9968 16058 10002
rect 16000 9934 16058 9968
rect 16000 9900 16012 9934
rect 16046 9900 16058 9934
rect 16000 9866 16058 9900
rect 16000 9832 16012 9866
rect 16046 9832 16058 9866
rect 16000 9798 16058 9832
rect 16000 9764 16012 9798
rect 16046 9764 16058 9798
rect 16000 9730 16058 9764
rect 16000 9696 16012 9730
rect 16046 9696 16058 9730
rect 16000 9662 16058 9696
rect 16000 9628 16012 9662
rect 16046 9628 16058 9662
rect 16000 9594 16058 9628
rect 16000 9560 16012 9594
rect 16046 9560 16058 9594
rect 16000 9526 16058 9560
rect 16000 9492 16012 9526
rect 16046 9492 16058 9526
rect 16000 9458 16058 9492
rect 16000 9424 16012 9458
rect 16046 9424 16058 9458
rect 16000 9390 16058 9424
rect 16000 9356 16012 9390
rect 16046 9356 16058 9390
rect 16000 9322 16058 9356
rect 16000 9288 16012 9322
rect 16046 9288 16058 9322
rect 16000 9254 16058 9288
rect 16000 9220 16012 9254
rect 16046 9220 16058 9254
rect 16000 9186 16058 9220
rect 16000 9152 16012 9186
rect 16046 9152 16058 9186
rect 16000 9118 16058 9152
rect 16000 9084 16012 9118
rect 16046 9084 16058 9118
rect 16000 9050 16058 9084
rect 16000 9016 16012 9050
rect 16046 9016 16058 9050
rect 16000 8982 16058 9016
rect 16000 8948 16012 8982
rect 16046 8948 16058 8982
rect 16000 8914 16058 8948
rect 16000 8880 16012 8914
rect 16046 8880 16058 8914
rect 16000 8846 16058 8880
rect 16000 8812 16012 8846
rect 16046 8812 16058 8846
rect 16000 8778 16058 8812
rect 16000 8744 16012 8778
rect 16046 8744 16058 8778
rect 16000 8710 16058 8744
rect 16000 8676 16012 8710
rect 16046 8676 16058 8710
rect 16000 8642 16058 8676
rect 16000 8608 16012 8642
rect 16046 8608 16058 8642
rect 16000 8574 16058 8608
rect 16000 8540 16012 8574
rect 16046 8540 16058 8574
rect 16000 8506 16058 8540
rect 16000 8472 16012 8506
rect 16046 8472 16058 8506
rect 16000 8438 16058 8472
rect 16000 8404 16012 8438
rect 16046 8404 16058 8438
rect 16000 8370 16058 8404
rect 16000 8336 16012 8370
rect 16046 8336 16058 8370
rect 16000 8302 16058 8336
rect 16000 8268 16012 8302
rect 16046 8268 16058 8302
rect 16000 8247 16058 8268
rect 17058 11226 17116 11247
rect 17058 11192 17070 11226
rect 17104 11192 17116 11226
rect 17058 11158 17116 11192
rect 17058 11124 17070 11158
rect 17104 11124 17116 11158
rect 17058 11090 17116 11124
rect 17058 11056 17070 11090
rect 17104 11056 17116 11090
rect 17058 11022 17116 11056
rect 17058 10988 17070 11022
rect 17104 10988 17116 11022
rect 17058 10954 17116 10988
rect 17058 10920 17070 10954
rect 17104 10920 17116 10954
rect 17058 10886 17116 10920
rect 17058 10852 17070 10886
rect 17104 10852 17116 10886
rect 17058 10818 17116 10852
rect 17058 10784 17070 10818
rect 17104 10784 17116 10818
rect 17058 10750 17116 10784
rect 17058 10716 17070 10750
rect 17104 10716 17116 10750
rect 17058 10682 17116 10716
rect 17058 10648 17070 10682
rect 17104 10648 17116 10682
rect 17058 10614 17116 10648
rect 17058 10580 17070 10614
rect 17104 10580 17116 10614
rect 17058 10546 17116 10580
rect 17058 10512 17070 10546
rect 17104 10512 17116 10546
rect 17058 10478 17116 10512
rect 17058 10444 17070 10478
rect 17104 10444 17116 10478
rect 17058 10410 17116 10444
rect 17058 10376 17070 10410
rect 17104 10376 17116 10410
rect 17058 10342 17116 10376
rect 17058 10308 17070 10342
rect 17104 10308 17116 10342
rect 17058 10274 17116 10308
rect 17058 10240 17070 10274
rect 17104 10240 17116 10274
rect 17058 10206 17116 10240
rect 17058 10172 17070 10206
rect 17104 10172 17116 10206
rect 17058 10138 17116 10172
rect 17058 10104 17070 10138
rect 17104 10104 17116 10138
rect 17058 10070 17116 10104
rect 17058 10036 17070 10070
rect 17104 10036 17116 10070
rect 17058 10002 17116 10036
rect 17058 9968 17070 10002
rect 17104 9968 17116 10002
rect 17058 9934 17116 9968
rect 17058 9900 17070 9934
rect 17104 9900 17116 9934
rect 17058 9866 17116 9900
rect 17058 9832 17070 9866
rect 17104 9832 17116 9866
rect 17058 9798 17116 9832
rect 17058 9764 17070 9798
rect 17104 9764 17116 9798
rect 17058 9730 17116 9764
rect 17058 9696 17070 9730
rect 17104 9696 17116 9730
rect 17058 9662 17116 9696
rect 17058 9628 17070 9662
rect 17104 9628 17116 9662
rect 17058 9594 17116 9628
rect 17058 9560 17070 9594
rect 17104 9560 17116 9594
rect 17058 9526 17116 9560
rect 17058 9492 17070 9526
rect 17104 9492 17116 9526
rect 17058 9458 17116 9492
rect 17058 9424 17070 9458
rect 17104 9424 17116 9458
rect 17058 9390 17116 9424
rect 17058 9356 17070 9390
rect 17104 9356 17116 9390
rect 17058 9322 17116 9356
rect 17058 9288 17070 9322
rect 17104 9288 17116 9322
rect 17058 9254 17116 9288
rect 17058 9220 17070 9254
rect 17104 9220 17116 9254
rect 17058 9186 17116 9220
rect 17058 9152 17070 9186
rect 17104 9152 17116 9186
rect 17058 9118 17116 9152
rect 17058 9084 17070 9118
rect 17104 9084 17116 9118
rect 17058 9050 17116 9084
rect 17058 9016 17070 9050
rect 17104 9016 17116 9050
rect 17058 8982 17116 9016
rect 17058 8948 17070 8982
rect 17104 8948 17116 8982
rect 17058 8914 17116 8948
rect 17058 8880 17070 8914
rect 17104 8880 17116 8914
rect 17058 8846 17116 8880
rect 17058 8812 17070 8846
rect 17104 8812 17116 8846
rect 17058 8778 17116 8812
rect 17058 8744 17070 8778
rect 17104 8744 17116 8778
rect 17058 8710 17116 8744
rect 17058 8676 17070 8710
rect 17104 8676 17116 8710
rect 17058 8642 17116 8676
rect 17058 8608 17070 8642
rect 17104 8608 17116 8642
rect 17058 8574 17116 8608
rect 17058 8540 17070 8574
rect 17104 8540 17116 8574
rect 17058 8506 17116 8540
rect 17058 8472 17070 8506
rect 17104 8472 17116 8506
rect 17058 8438 17116 8472
rect 17058 8404 17070 8438
rect 17104 8404 17116 8438
rect 17058 8370 17116 8404
rect 17058 8336 17070 8370
rect 17104 8336 17116 8370
rect 17058 8302 17116 8336
rect 17058 8268 17070 8302
rect 17104 8268 17116 8302
rect 17058 8247 17116 8268
rect 17466 11200 17524 11221
rect 17466 11166 17478 11200
rect 17512 11166 17524 11200
rect 17466 11132 17524 11166
rect 17466 11098 17478 11132
rect 17512 11098 17524 11132
rect 17466 11064 17524 11098
rect 17466 11030 17478 11064
rect 17512 11030 17524 11064
rect 17466 10996 17524 11030
rect 17466 10962 17478 10996
rect 17512 10962 17524 10996
rect 17466 10928 17524 10962
rect 17466 10894 17478 10928
rect 17512 10894 17524 10928
rect 17466 10860 17524 10894
rect 17466 10826 17478 10860
rect 17512 10826 17524 10860
rect 17466 10792 17524 10826
rect 17466 10758 17478 10792
rect 17512 10758 17524 10792
rect 17466 10724 17524 10758
rect 17466 10690 17478 10724
rect 17512 10690 17524 10724
rect 17466 10656 17524 10690
rect 17466 10622 17478 10656
rect 17512 10622 17524 10656
rect 17466 10588 17524 10622
rect 17466 10554 17478 10588
rect 17512 10554 17524 10588
rect 17466 10520 17524 10554
rect 17466 10486 17478 10520
rect 17512 10486 17524 10520
rect 17466 10452 17524 10486
rect 17466 10418 17478 10452
rect 17512 10418 17524 10452
rect 17466 10384 17524 10418
rect 17466 10350 17478 10384
rect 17512 10350 17524 10384
rect 17466 10316 17524 10350
rect 17466 10282 17478 10316
rect 17512 10282 17524 10316
rect 17466 10248 17524 10282
rect 17466 10214 17478 10248
rect 17512 10214 17524 10248
rect 17466 10180 17524 10214
rect 17466 10146 17478 10180
rect 17512 10146 17524 10180
rect 17466 10112 17524 10146
rect 17466 10078 17478 10112
rect 17512 10078 17524 10112
rect 17466 10044 17524 10078
rect 17466 10010 17478 10044
rect 17512 10010 17524 10044
rect 17466 9976 17524 10010
rect 17466 9942 17478 9976
rect 17512 9942 17524 9976
rect 17466 9908 17524 9942
rect 17466 9874 17478 9908
rect 17512 9874 17524 9908
rect 17466 9840 17524 9874
rect 17466 9806 17478 9840
rect 17512 9806 17524 9840
rect 17466 9772 17524 9806
rect 17466 9738 17478 9772
rect 17512 9738 17524 9772
rect 17466 9704 17524 9738
rect 17466 9670 17478 9704
rect 17512 9670 17524 9704
rect 17466 9636 17524 9670
rect 17466 9602 17478 9636
rect 17512 9602 17524 9636
rect 17466 9568 17524 9602
rect 17466 9534 17478 9568
rect 17512 9534 17524 9568
rect 17466 9500 17524 9534
rect 17466 9466 17478 9500
rect 17512 9466 17524 9500
rect 17466 9432 17524 9466
rect 17466 9398 17478 9432
rect 17512 9398 17524 9432
rect 17466 9364 17524 9398
rect 17466 9330 17478 9364
rect 17512 9330 17524 9364
rect 17466 9296 17524 9330
rect 17466 9262 17478 9296
rect 17512 9262 17524 9296
rect 17466 9228 17524 9262
rect 17466 9194 17478 9228
rect 17512 9194 17524 9228
rect 17466 9160 17524 9194
rect 17466 9126 17478 9160
rect 17512 9126 17524 9160
rect 17466 9092 17524 9126
rect 17466 9058 17478 9092
rect 17512 9058 17524 9092
rect 17466 9024 17524 9058
rect 17466 8990 17478 9024
rect 17512 8990 17524 9024
rect 17466 8956 17524 8990
rect 17466 8922 17478 8956
rect 17512 8922 17524 8956
rect 17466 8888 17524 8922
rect 17466 8854 17478 8888
rect 17512 8854 17524 8888
rect 17466 8820 17524 8854
rect 17466 8786 17478 8820
rect 17512 8786 17524 8820
rect 17466 8752 17524 8786
rect 17466 8718 17478 8752
rect 17512 8718 17524 8752
rect 17466 8684 17524 8718
rect 17466 8650 17478 8684
rect 17512 8650 17524 8684
rect 17466 8616 17524 8650
rect 17466 8582 17478 8616
rect 17512 8582 17524 8616
rect 17466 8548 17524 8582
rect 17466 8514 17478 8548
rect 17512 8514 17524 8548
rect 17466 8480 17524 8514
rect 17466 8446 17478 8480
rect 17512 8446 17524 8480
rect 17466 8412 17524 8446
rect 17466 8378 17478 8412
rect 17512 8378 17524 8412
rect 17466 8344 17524 8378
rect 17466 8310 17478 8344
rect 17512 8310 17524 8344
rect 17466 8276 17524 8310
rect 17466 8242 17478 8276
rect 17512 8242 17524 8276
rect 17466 8221 17524 8242
rect 18524 11200 18582 11221
rect 18524 11166 18536 11200
rect 18570 11166 18582 11200
rect 18524 11132 18582 11166
rect 18524 11098 18536 11132
rect 18570 11098 18582 11132
rect 18524 11064 18582 11098
rect 18524 11030 18536 11064
rect 18570 11030 18582 11064
rect 18524 10996 18582 11030
rect 18524 10962 18536 10996
rect 18570 10962 18582 10996
rect 18524 10928 18582 10962
rect 18524 10894 18536 10928
rect 18570 10894 18582 10928
rect 18524 10860 18582 10894
rect 18524 10826 18536 10860
rect 18570 10826 18582 10860
rect 18524 10792 18582 10826
rect 18524 10758 18536 10792
rect 18570 10758 18582 10792
rect 18524 10724 18582 10758
rect 18524 10690 18536 10724
rect 18570 10690 18582 10724
rect 18524 10656 18582 10690
rect 18524 10622 18536 10656
rect 18570 10622 18582 10656
rect 18524 10588 18582 10622
rect 18524 10554 18536 10588
rect 18570 10554 18582 10588
rect 18524 10520 18582 10554
rect 18524 10486 18536 10520
rect 18570 10486 18582 10520
rect 18524 10452 18582 10486
rect 18524 10418 18536 10452
rect 18570 10418 18582 10452
rect 18524 10384 18582 10418
rect 18524 10350 18536 10384
rect 18570 10350 18582 10384
rect 18524 10316 18582 10350
rect 18524 10282 18536 10316
rect 18570 10282 18582 10316
rect 18524 10248 18582 10282
rect 18524 10214 18536 10248
rect 18570 10214 18582 10248
rect 18524 10180 18582 10214
rect 18524 10146 18536 10180
rect 18570 10146 18582 10180
rect 18524 10112 18582 10146
rect 18524 10078 18536 10112
rect 18570 10078 18582 10112
rect 18524 10044 18582 10078
rect 18524 10010 18536 10044
rect 18570 10010 18582 10044
rect 18524 9976 18582 10010
rect 18524 9942 18536 9976
rect 18570 9942 18582 9976
rect 18524 9908 18582 9942
rect 18524 9874 18536 9908
rect 18570 9874 18582 9908
rect 18524 9840 18582 9874
rect 18524 9806 18536 9840
rect 18570 9806 18582 9840
rect 18524 9772 18582 9806
rect 18524 9738 18536 9772
rect 18570 9738 18582 9772
rect 18524 9704 18582 9738
rect 18524 9670 18536 9704
rect 18570 9670 18582 9704
rect 18524 9636 18582 9670
rect 18524 9602 18536 9636
rect 18570 9602 18582 9636
rect 18524 9568 18582 9602
rect 18524 9534 18536 9568
rect 18570 9534 18582 9568
rect 18524 9500 18582 9534
rect 18524 9466 18536 9500
rect 18570 9466 18582 9500
rect 18524 9432 18582 9466
rect 18524 9398 18536 9432
rect 18570 9398 18582 9432
rect 18524 9364 18582 9398
rect 18524 9330 18536 9364
rect 18570 9330 18582 9364
rect 18524 9296 18582 9330
rect 18524 9262 18536 9296
rect 18570 9262 18582 9296
rect 18524 9228 18582 9262
rect 18524 9194 18536 9228
rect 18570 9194 18582 9228
rect 18524 9160 18582 9194
rect 18524 9126 18536 9160
rect 18570 9126 18582 9160
rect 18524 9092 18582 9126
rect 18524 9058 18536 9092
rect 18570 9058 18582 9092
rect 18524 9024 18582 9058
rect 18524 8990 18536 9024
rect 18570 8990 18582 9024
rect 18524 8956 18582 8990
rect 18524 8922 18536 8956
rect 18570 8922 18582 8956
rect 18524 8888 18582 8922
rect 18524 8854 18536 8888
rect 18570 8854 18582 8888
rect 18524 8820 18582 8854
rect 18524 8786 18536 8820
rect 18570 8786 18582 8820
rect 18524 8752 18582 8786
rect 18524 8718 18536 8752
rect 18570 8718 18582 8752
rect 18524 8684 18582 8718
rect 18524 8650 18536 8684
rect 18570 8650 18582 8684
rect 18524 8616 18582 8650
rect 18524 8582 18536 8616
rect 18570 8582 18582 8616
rect 18524 8548 18582 8582
rect 18524 8514 18536 8548
rect 18570 8514 18582 8548
rect 18524 8480 18582 8514
rect 18524 8446 18536 8480
rect 18570 8446 18582 8480
rect 18524 8412 18582 8446
rect 18524 8378 18536 8412
rect 18570 8378 18582 8412
rect 18524 8344 18582 8378
rect 18524 8310 18536 8344
rect 18570 8310 18582 8344
rect 18524 8276 18582 8310
rect 18524 8242 18536 8276
rect 18570 8242 18582 8276
rect 18524 8221 18582 8242
rect 19582 11200 19640 11221
rect 19582 11166 19594 11200
rect 19628 11166 19640 11200
rect 19582 11132 19640 11166
rect 19582 11098 19594 11132
rect 19628 11098 19640 11132
rect 19582 11064 19640 11098
rect 19582 11030 19594 11064
rect 19628 11030 19640 11064
rect 19582 10996 19640 11030
rect 19582 10962 19594 10996
rect 19628 10962 19640 10996
rect 19582 10928 19640 10962
rect 19582 10894 19594 10928
rect 19628 10894 19640 10928
rect 19582 10860 19640 10894
rect 19582 10826 19594 10860
rect 19628 10826 19640 10860
rect 19582 10792 19640 10826
rect 19582 10758 19594 10792
rect 19628 10758 19640 10792
rect 19582 10724 19640 10758
rect 19582 10690 19594 10724
rect 19628 10690 19640 10724
rect 19582 10656 19640 10690
rect 19582 10622 19594 10656
rect 19628 10622 19640 10656
rect 19582 10588 19640 10622
rect 19582 10554 19594 10588
rect 19628 10554 19640 10588
rect 19582 10520 19640 10554
rect 19582 10486 19594 10520
rect 19628 10486 19640 10520
rect 19582 10452 19640 10486
rect 19582 10418 19594 10452
rect 19628 10418 19640 10452
rect 19582 10384 19640 10418
rect 19582 10350 19594 10384
rect 19628 10350 19640 10384
rect 19582 10316 19640 10350
rect 19582 10282 19594 10316
rect 19628 10282 19640 10316
rect 19582 10248 19640 10282
rect 19582 10214 19594 10248
rect 19628 10214 19640 10248
rect 19582 10180 19640 10214
rect 19582 10146 19594 10180
rect 19628 10146 19640 10180
rect 19582 10112 19640 10146
rect 19582 10078 19594 10112
rect 19628 10078 19640 10112
rect 19582 10044 19640 10078
rect 19582 10010 19594 10044
rect 19628 10010 19640 10044
rect 19582 9976 19640 10010
rect 19582 9942 19594 9976
rect 19628 9942 19640 9976
rect 19582 9908 19640 9942
rect 19582 9874 19594 9908
rect 19628 9874 19640 9908
rect 19582 9840 19640 9874
rect 19582 9806 19594 9840
rect 19628 9806 19640 9840
rect 19582 9772 19640 9806
rect 19582 9738 19594 9772
rect 19628 9738 19640 9772
rect 19582 9704 19640 9738
rect 19582 9670 19594 9704
rect 19628 9670 19640 9704
rect 19582 9636 19640 9670
rect 19582 9602 19594 9636
rect 19628 9602 19640 9636
rect 19582 9568 19640 9602
rect 19582 9534 19594 9568
rect 19628 9534 19640 9568
rect 19582 9500 19640 9534
rect 19582 9466 19594 9500
rect 19628 9466 19640 9500
rect 19582 9432 19640 9466
rect 19582 9398 19594 9432
rect 19628 9398 19640 9432
rect 19582 9364 19640 9398
rect 19582 9330 19594 9364
rect 19628 9330 19640 9364
rect 19582 9296 19640 9330
rect 19582 9262 19594 9296
rect 19628 9262 19640 9296
rect 19582 9228 19640 9262
rect 19582 9194 19594 9228
rect 19628 9194 19640 9228
rect 19582 9160 19640 9194
rect 19582 9126 19594 9160
rect 19628 9126 19640 9160
rect 19582 9092 19640 9126
rect 19582 9058 19594 9092
rect 19628 9058 19640 9092
rect 19582 9024 19640 9058
rect 19582 8990 19594 9024
rect 19628 8990 19640 9024
rect 19582 8956 19640 8990
rect 19582 8922 19594 8956
rect 19628 8922 19640 8956
rect 19582 8888 19640 8922
rect 19582 8854 19594 8888
rect 19628 8854 19640 8888
rect 19582 8820 19640 8854
rect 19582 8786 19594 8820
rect 19628 8786 19640 8820
rect 19582 8752 19640 8786
rect 19582 8718 19594 8752
rect 19628 8718 19640 8752
rect 19582 8684 19640 8718
rect 19582 8650 19594 8684
rect 19628 8650 19640 8684
rect 19582 8616 19640 8650
rect 19582 8582 19594 8616
rect 19628 8582 19640 8616
rect 19582 8548 19640 8582
rect 19582 8514 19594 8548
rect 19628 8514 19640 8548
rect 19582 8480 19640 8514
rect 19582 8446 19594 8480
rect 19628 8446 19640 8480
rect 19582 8412 19640 8446
rect 19582 8378 19594 8412
rect 19628 8378 19640 8412
rect 19582 8344 19640 8378
rect 19582 8310 19594 8344
rect 19628 8310 19640 8344
rect 19582 8276 19640 8310
rect 19582 8242 19594 8276
rect 19628 8242 19640 8276
rect 19582 8221 19640 8242
rect 23209 13356 24209 13368
rect 23209 13322 23250 13356
rect 23284 13322 23318 13356
rect 23352 13322 23386 13356
rect 23420 13322 23454 13356
rect 23488 13322 23522 13356
rect 23556 13322 23590 13356
rect 23624 13322 23658 13356
rect 23692 13322 23726 13356
rect 23760 13322 23794 13356
rect 23828 13322 23862 13356
rect 23896 13322 23930 13356
rect 23964 13322 23998 13356
rect 24032 13322 24066 13356
rect 24100 13322 24134 13356
rect 24168 13322 24209 13356
rect 23209 13310 24209 13322
rect 23209 12298 24209 12310
rect 23209 12264 23250 12298
rect 23284 12264 23318 12298
rect 23352 12264 23386 12298
rect 23420 12264 23454 12298
rect 23488 12264 23522 12298
rect 23556 12264 23590 12298
rect 23624 12264 23658 12298
rect 23692 12264 23726 12298
rect 23760 12264 23794 12298
rect 23828 12264 23862 12298
rect 23896 12264 23930 12298
rect 23964 12264 23998 12298
rect 24032 12264 24066 12298
rect 24100 12264 24134 12298
rect 24168 12264 24209 12298
rect 23209 12252 24209 12264
rect 24769 13350 25769 13362
rect 24769 13316 24810 13350
rect 24844 13316 24878 13350
rect 24912 13316 24946 13350
rect 24980 13316 25014 13350
rect 25048 13316 25082 13350
rect 25116 13316 25150 13350
rect 25184 13316 25218 13350
rect 25252 13316 25286 13350
rect 25320 13316 25354 13350
rect 25388 13316 25422 13350
rect 25456 13316 25490 13350
rect 25524 13316 25558 13350
rect 25592 13316 25626 13350
rect 25660 13316 25694 13350
rect 25728 13316 25769 13350
rect 24769 13304 25769 13316
rect 24769 12292 25769 12304
rect 24769 12258 24810 12292
rect 24844 12258 24878 12292
rect 24912 12258 24946 12292
rect 24980 12258 25014 12292
rect 25048 12258 25082 12292
rect 25116 12258 25150 12292
rect 25184 12258 25218 12292
rect 25252 12258 25286 12292
rect 25320 12258 25354 12292
rect 25388 12258 25422 12292
rect 25456 12258 25490 12292
rect 25524 12258 25558 12292
rect 25592 12258 25626 12292
rect 25660 12258 25694 12292
rect 25728 12258 25769 12292
rect 24769 12246 25769 12258
rect 24769 11234 25769 11246
rect 24769 11200 24810 11234
rect 24844 11200 24878 11234
rect 24912 11200 24946 11234
rect 24980 11200 25014 11234
rect 25048 11200 25082 11234
rect 25116 11200 25150 11234
rect 25184 11200 25218 11234
rect 25252 11200 25286 11234
rect 25320 11200 25354 11234
rect 25388 11200 25422 11234
rect 25456 11200 25490 11234
rect 25524 11200 25558 11234
rect 25592 11200 25626 11234
rect 25660 11200 25694 11234
rect 25728 11200 25769 11234
rect 24769 11188 25769 11200
rect 24769 10176 25769 10188
rect 24769 10142 24810 10176
rect 24844 10142 24878 10176
rect 24912 10142 24946 10176
rect 24980 10142 25014 10176
rect 25048 10142 25082 10176
rect 25116 10142 25150 10176
rect 25184 10142 25218 10176
rect 25252 10142 25286 10176
rect 25320 10142 25354 10176
rect 25388 10142 25422 10176
rect 25456 10142 25490 10176
rect 25524 10142 25558 10176
rect 25592 10142 25626 10176
rect 25660 10142 25694 10176
rect 25728 10142 25769 10176
rect 24769 10130 25769 10142
rect 24769 9118 25769 9130
rect 24769 9084 24810 9118
rect 24844 9084 24878 9118
rect 24912 9084 24946 9118
rect 24980 9084 25014 9118
rect 25048 9084 25082 9118
rect 25116 9084 25150 9118
rect 25184 9084 25218 9118
rect 25252 9084 25286 9118
rect 25320 9084 25354 9118
rect 25388 9084 25422 9118
rect 25456 9084 25490 9118
rect 25524 9084 25558 9118
rect 25592 9084 25626 9118
rect 25660 9084 25694 9118
rect 25728 9084 25769 9118
rect 24769 9072 25769 9084
<< pdiffc >>
rect 23468 15462 23502 15496
rect 23558 15462 23592 15496
rect 23648 15462 23682 15496
rect 23738 15462 23772 15496
rect 23828 15462 23862 15496
rect 23918 15462 23952 15496
rect 24008 15462 24042 15496
rect 23468 15372 23502 15406
rect 23558 15372 23592 15406
rect 23648 15372 23682 15406
rect 23738 15372 23772 15406
rect 23828 15372 23862 15406
rect 23918 15372 23952 15406
rect 24008 15372 24042 15406
rect 23468 15282 23502 15316
rect 23558 15282 23592 15316
rect 23648 15282 23682 15316
rect 23738 15282 23772 15316
rect 23828 15282 23862 15316
rect 23918 15282 23952 15316
rect 24008 15282 24042 15316
rect 23468 15192 23502 15226
rect 23558 15192 23592 15226
rect 23648 15192 23682 15226
rect 23738 15192 23772 15226
rect 23828 15192 23862 15226
rect 23918 15192 23952 15226
rect 24008 15192 24042 15226
rect 23468 15102 23502 15136
rect 23558 15102 23592 15136
rect 23648 15102 23682 15136
rect 23738 15102 23772 15136
rect 23828 15102 23862 15136
rect 23918 15102 23952 15136
rect 24008 15102 24042 15136
rect 23468 15012 23502 15046
rect 23558 15012 23592 15046
rect 23648 15012 23682 15046
rect 23738 15012 23772 15046
rect 23828 15012 23862 15046
rect 23918 15012 23952 15046
rect 24008 15012 24042 15046
rect 23468 14922 23502 14956
rect 23558 14922 23592 14956
rect 23648 14922 23682 14956
rect 23738 14922 23772 14956
rect 23828 14922 23862 14956
rect 23918 14922 23952 14956
rect 24008 14922 24042 14956
rect 13140 10944 13174 10978
rect 13230 10944 13264 10978
rect 13320 10944 13354 10978
rect 13410 10944 13444 10978
rect 13500 10944 13534 10978
rect 13590 10944 13624 10978
rect 13680 10944 13714 10978
rect 13140 10854 13174 10888
rect 13230 10854 13264 10888
rect 13320 10854 13354 10888
rect 13410 10854 13444 10888
rect 13500 10854 13534 10888
rect 13590 10854 13624 10888
rect 13680 10854 13714 10888
rect 13140 10764 13174 10798
rect 13230 10764 13264 10798
rect 13320 10764 13354 10798
rect 13410 10764 13444 10798
rect 13500 10764 13534 10798
rect 13590 10764 13624 10798
rect 13680 10764 13714 10798
rect 13140 10674 13174 10708
rect 13230 10674 13264 10708
rect 13320 10674 13354 10708
rect 13410 10674 13444 10708
rect 13500 10674 13534 10708
rect 13590 10674 13624 10708
rect 13680 10674 13714 10708
rect 13140 10584 13174 10618
rect 13230 10584 13264 10618
rect 13320 10584 13354 10618
rect 13410 10584 13444 10618
rect 13500 10584 13534 10618
rect 13590 10584 13624 10618
rect 13680 10584 13714 10618
rect 13140 10494 13174 10528
rect 13230 10494 13264 10528
rect 13320 10494 13354 10528
rect 13410 10494 13444 10528
rect 13500 10494 13534 10528
rect 13590 10494 13624 10528
rect 13680 10494 13714 10528
rect 13140 10404 13174 10438
rect 13230 10404 13264 10438
rect 13320 10404 13354 10438
rect 13410 10404 13444 10438
rect 13500 10404 13534 10438
rect 13590 10404 13624 10438
rect 13680 10404 13714 10438
rect 13140 9454 13174 9488
rect 13230 9454 13264 9488
rect 13320 9454 13354 9488
rect 13410 9454 13444 9488
rect 13500 9454 13534 9488
rect 13590 9454 13624 9488
rect 13680 9454 13714 9488
rect 13140 9364 13174 9398
rect 13230 9364 13264 9398
rect 13320 9364 13354 9398
rect 13410 9364 13444 9398
rect 13500 9364 13534 9398
rect 13590 9364 13624 9398
rect 13680 9364 13714 9398
rect 13140 9274 13174 9308
rect 13230 9274 13264 9308
rect 13320 9274 13354 9308
rect 13410 9274 13444 9308
rect 13500 9274 13534 9308
rect 13590 9274 13624 9308
rect 13680 9274 13714 9308
rect 13140 9184 13174 9218
rect 13230 9184 13264 9218
rect 13320 9184 13354 9218
rect 13410 9184 13444 9218
rect 13500 9184 13534 9218
rect 13590 9184 13624 9218
rect 13680 9184 13714 9218
rect 13140 9094 13174 9128
rect 13230 9094 13264 9128
rect 13320 9094 13354 9128
rect 13410 9094 13444 9128
rect 13500 9094 13534 9128
rect 13590 9094 13624 9128
rect 13680 9094 13714 9128
rect 13140 9004 13174 9038
rect 13230 9004 13264 9038
rect 13320 9004 13354 9038
rect 13410 9004 13444 9038
rect 13500 9004 13534 9038
rect 13590 9004 13624 9038
rect 13680 9004 13714 9038
rect 13140 8914 13174 8948
rect 13230 8914 13264 8948
rect 13320 8914 13354 8948
rect 13410 8914 13444 8948
rect 13500 8914 13534 8948
rect 13590 8914 13624 8948
rect 13680 8914 13714 8948
rect 13130 8044 13164 8078
rect 13220 8044 13254 8078
rect 13310 8044 13344 8078
rect 13400 8044 13434 8078
rect 13490 8044 13524 8078
rect 13580 8044 13614 8078
rect 13670 8044 13704 8078
rect 13130 7954 13164 7988
rect 13220 7954 13254 7988
rect 13310 7954 13344 7988
rect 13400 7954 13434 7988
rect 13490 7954 13524 7988
rect 13580 7954 13614 7988
rect 13670 7954 13704 7988
rect 13130 7864 13164 7898
rect 13220 7864 13254 7898
rect 13310 7864 13344 7898
rect 13400 7864 13434 7898
rect 13490 7864 13524 7898
rect 13580 7864 13614 7898
rect 13670 7864 13704 7898
rect 13130 7774 13164 7808
rect 13220 7774 13254 7808
rect 13310 7774 13344 7808
rect 13400 7774 13434 7808
rect 13490 7774 13524 7808
rect 13580 7774 13614 7808
rect 13670 7774 13704 7808
rect 13130 7684 13164 7718
rect 13220 7684 13254 7718
rect 13310 7684 13344 7718
rect 13400 7684 13434 7718
rect 13490 7684 13524 7718
rect 13580 7684 13614 7718
rect 13670 7684 13704 7718
rect 13130 7594 13164 7628
rect 13220 7594 13254 7628
rect 13310 7594 13344 7628
rect 13400 7594 13434 7628
rect 13490 7594 13524 7628
rect 13580 7594 13614 7628
rect 13670 7594 13704 7628
rect 13130 7504 13164 7538
rect 13220 7504 13254 7538
rect 13310 7504 13344 7538
rect 13400 7504 13434 7538
rect 13490 7504 13524 7538
rect 13580 7504 13614 7538
rect 13670 7504 13704 7538
rect 13130 6694 13164 6728
rect 13220 6694 13254 6728
rect 13310 6694 13344 6728
rect 13400 6694 13434 6728
rect 13490 6694 13524 6728
rect 13580 6694 13614 6728
rect 13670 6694 13704 6728
rect 13130 6604 13164 6638
rect 13220 6604 13254 6638
rect 13310 6604 13344 6638
rect 13400 6604 13434 6638
rect 13490 6604 13524 6638
rect 13580 6604 13614 6638
rect 13670 6604 13704 6638
rect 13130 6514 13164 6548
rect 13220 6514 13254 6548
rect 13310 6514 13344 6548
rect 13400 6514 13434 6548
rect 13490 6514 13524 6548
rect 13580 6514 13614 6548
rect 13670 6514 13704 6548
rect 13130 6424 13164 6458
rect 13220 6424 13254 6458
rect 13310 6424 13344 6458
rect 13400 6424 13434 6458
rect 13490 6424 13524 6458
rect 13580 6424 13614 6458
rect 13670 6424 13704 6458
rect 13130 6334 13164 6368
rect 13220 6334 13254 6368
rect 13310 6334 13344 6368
rect 13400 6334 13434 6368
rect 13490 6334 13524 6368
rect 13580 6334 13614 6368
rect 13670 6334 13704 6368
rect 13130 6244 13164 6278
rect 13220 6244 13254 6278
rect 13310 6244 13344 6278
rect 13400 6244 13434 6278
rect 13490 6244 13524 6278
rect 13580 6244 13614 6278
rect 13670 6244 13704 6278
rect 13130 6154 13164 6188
rect 13220 6154 13254 6188
rect 13310 6154 13344 6188
rect 13400 6154 13434 6188
rect 13490 6154 13524 6188
rect 13580 6154 13614 6188
rect 13670 6154 13704 6188
rect 14780 6724 14814 6758
rect 14870 6724 14904 6758
rect 14960 6724 14994 6758
rect 15050 6724 15084 6758
rect 15140 6724 15174 6758
rect 15230 6724 15264 6758
rect 15320 6724 15354 6758
rect 14780 6634 14814 6668
rect 14870 6634 14904 6668
rect 14960 6634 14994 6668
rect 15050 6634 15084 6668
rect 15140 6634 15174 6668
rect 15230 6634 15264 6668
rect 15320 6634 15354 6668
rect 14780 6544 14814 6578
rect 14870 6544 14904 6578
rect 14960 6544 14994 6578
rect 15050 6544 15084 6578
rect 15140 6544 15174 6578
rect 15230 6544 15264 6578
rect 15320 6544 15354 6578
rect 14780 6454 14814 6488
rect 14870 6454 14904 6488
rect 14960 6454 14994 6488
rect 15050 6454 15084 6488
rect 15140 6454 15174 6488
rect 15230 6454 15264 6488
rect 15320 6454 15354 6488
rect 14780 6364 14814 6398
rect 14870 6364 14904 6398
rect 14960 6364 14994 6398
rect 15050 6364 15084 6398
rect 15140 6364 15174 6398
rect 15230 6364 15264 6398
rect 15320 6364 15354 6398
rect 14780 6274 14814 6308
rect 14870 6274 14904 6308
rect 14960 6274 14994 6308
rect 15050 6274 15084 6308
rect 15140 6274 15174 6308
rect 15230 6274 15264 6308
rect 15320 6274 15354 6308
rect 14780 6184 14814 6218
rect 14870 6184 14904 6218
rect 14960 6184 14994 6218
rect 15050 6184 15084 6218
rect 15140 6184 15174 6218
rect 15230 6184 15264 6218
rect 15320 6184 15354 6218
rect 13130 5344 13164 5378
rect 13220 5344 13254 5378
rect 13310 5344 13344 5378
rect 13400 5344 13434 5378
rect 13490 5344 13524 5378
rect 13580 5344 13614 5378
rect 13670 5344 13704 5378
rect 13130 5254 13164 5288
rect 13220 5254 13254 5288
rect 13310 5254 13344 5288
rect 13400 5254 13434 5288
rect 13490 5254 13524 5288
rect 13580 5254 13614 5288
rect 13670 5254 13704 5288
rect 13130 5164 13164 5198
rect 13220 5164 13254 5198
rect 13310 5164 13344 5198
rect 13400 5164 13434 5198
rect 13490 5164 13524 5198
rect 13580 5164 13614 5198
rect 13670 5164 13704 5198
rect 13130 5074 13164 5108
rect 13220 5074 13254 5108
rect 13310 5074 13344 5108
rect 13400 5074 13434 5108
rect 13490 5074 13524 5108
rect 13580 5074 13614 5108
rect 13670 5074 13704 5108
rect 13130 4984 13164 5018
rect 13220 4984 13254 5018
rect 13310 4984 13344 5018
rect 13400 4984 13434 5018
rect 13490 4984 13524 5018
rect 13580 4984 13614 5018
rect 13670 4984 13704 5018
rect 13130 4894 13164 4928
rect 13220 4894 13254 4928
rect 13310 4894 13344 4928
rect 13400 4894 13434 4928
rect 13490 4894 13524 4928
rect 13580 4894 13614 4928
rect 13670 4894 13704 4928
rect 13130 4804 13164 4838
rect 13220 4804 13254 4838
rect 13310 4804 13344 4838
rect 13400 4804 13434 4838
rect 13490 4804 13524 4838
rect 13580 4804 13614 4838
rect 13670 4804 13704 4838
rect 14780 5364 14814 5398
rect 14870 5364 14904 5398
rect 14960 5364 14994 5398
rect 15050 5364 15084 5398
rect 15140 5364 15174 5398
rect 15230 5364 15264 5398
rect 15320 5364 15354 5398
rect 14780 5274 14814 5308
rect 14870 5274 14904 5308
rect 14960 5274 14994 5308
rect 15050 5274 15084 5308
rect 15140 5274 15174 5308
rect 15230 5274 15264 5308
rect 15320 5274 15354 5308
rect 14780 5184 14814 5218
rect 14870 5184 14904 5218
rect 14960 5184 14994 5218
rect 15050 5184 15084 5218
rect 15140 5184 15174 5218
rect 15230 5184 15264 5218
rect 15320 5184 15354 5218
rect 14780 5094 14814 5128
rect 14870 5094 14904 5128
rect 14960 5094 14994 5128
rect 15050 5094 15084 5128
rect 15140 5094 15174 5128
rect 15230 5094 15264 5128
rect 15320 5094 15354 5128
rect 14780 5004 14814 5038
rect 14870 5004 14904 5038
rect 14960 5004 14994 5038
rect 15050 5004 15084 5038
rect 15140 5004 15174 5038
rect 15230 5004 15264 5038
rect 15320 5004 15354 5038
rect 14780 4914 14814 4948
rect 14870 4914 14904 4948
rect 14960 4914 14994 4948
rect 15050 4914 15084 4948
rect 15140 4914 15174 4948
rect 15230 4914 15264 4948
rect 15320 4914 15354 4948
rect 14780 4824 14814 4858
rect 14870 4824 14904 4858
rect 14960 4824 14994 4858
rect 15050 4824 15084 4858
rect 15140 4824 15174 4858
rect 15230 4824 15264 4858
rect 15320 4824 15354 4858
<< mvndiffc >>
rect 23150 17061 23184 17095
rect 23150 16993 23184 17027
rect 23150 16925 23184 16959
rect 23150 16857 23184 16891
rect 23150 16789 23184 16823
rect 23150 16721 23184 16755
rect 23150 16653 23184 16687
rect 23150 16585 23184 16619
rect 23150 16517 23184 16551
rect 23150 16449 23184 16483
rect 23150 16381 23184 16415
rect 23150 16313 23184 16347
rect 23150 16245 23184 16279
rect 23150 16177 23184 16211
rect 24208 17061 24242 17095
rect 24208 16993 24242 17027
rect 24208 16925 24242 16959
rect 24208 16857 24242 16891
rect 24208 16789 24242 16823
rect 24208 16721 24242 16755
rect 24208 16653 24242 16687
rect 24208 16585 24242 16619
rect 24208 16517 24242 16551
rect 24208 16449 24242 16483
rect 24208 16381 24242 16415
rect 24208 16313 24242 16347
rect 24208 16245 24242 16279
rect 24208 16177 24242 16211
rect -7459 14770 -7425 14804
rect -7459 14702 -7425 14736
rect -7459 14634 -7425 14668
rect -7459 14566 -7425 14600
rect -7459 14498 -7425 14532
rect -7459 14430 -7425 14464
rect -7459 14362 -7425 14396
rect -7459 14294 -7425 14328
rect -7459 14226 -7425 14260
rect -7459 14158 -7425 14192
rect -7459 14090 -7425 14124
rect -7459 14022 -7425 14056
rect -7459 13954 -7425 13988
rect -7459 13886 -7425 13920
rect -7459 13818 -7425 13852
rect -7459 13750 -7425 13784
rect -7459 13682 -7425 13716
rect -7459 13614 -7425 13648
rect -7459 13546 -7425 13580
rect -7459 13478 -7425 13512
rect -7459 13410 -7425 13444
rect -7459 13342 -7425 13376
rect -7459 13274 -7425 13308
rect -7459 13206 -7425 13240
rect -7459 13138 -7425 13172
rect -7459 13070 -7425 13104
rect -7459 13002 -7425 13036
rect -7459 12934 -7425 12968
rect -7459 12866 -7425 12900
rect -7201 14770 -7167 14804
rect -7201 14702 -7167 14736
rect -7201 14634 -7167 14668
rect -7201 14566 -7167 14600
rect -7201 14498 -7167 14532
rect -7201 14430 -7167 14464
rect -7201 14362 -7167 14396
rect -7201 14294 -7167 14328
rect -7201 14226 -7167 14260
rect -7201 14158 -7167 14192
rect -7201 14090 -7167 14124
rect -7201 14022 -7167 14056
rect -7201 13954 -7167 13988
rect -7201 13886 -7167 13920
rect -7201 13818 -7167 13852
rect -7201 13750 -7167 13784
rect -7201 13682 -7167 13716
rect -7201 13614 -7167 13648
rect -7201 13546 -7167 13580
rect -7201 13478 -7167 13512
rect -7201 13410 -7167 13444
rect -7201 13342 -7167 13376
rect -7201 13274 -7167 13308
rect -7201 13206 -7167 13240
rect -7201 13138 -7167 13172
rect -7201 13070 -7167 13104
rect -7201 13002 -7167 13036
rect -7201 12934 -7167 12968
rect -7201 12866 -7167 12900
rect -6943 14770 -6909 14804
rect -6943 14702 -6909 14736
rect -6943 14634 -6909 14668
rect -6943 14566 -6909 14600
rect -6943 14498 -6909 14532
rect -6943 14430 -6909 14464
rect -6943 14362 -6909 14396
rect -6943 14294 -6909 14328
rect -6943 14226 -6909 14260
rect -6943 14158 -6909 14192
rect -6943 14090 -6909 14124
rect -6943 14022 -6909 14056
rect -6943 13954 -6909 13988
rect -6943 13886 -6909 13920
rect -6943 13818 -6909 13852
rect -6943 13750 -6909 13784
rect -6943 13682 -6909 13716
rect -6943 13614 -6909 13648
rect -6943 13546 -6909 13580
rect -6943 13478 -6909 13512
rect -6943 13410 -6909 13444
rect -6943 13342 -6909 13376
rect -6943 13274 -6909 13308
rect -6943 13206 -6909 13240
rect -6943 13138 -6909 13172
rect -6943 13070 -6909 13104
rect -6943 13002 -6909 13036
rect -6943 12934 -6909 12968
rect -6943 12866 -6909 12900
rect -6685 14770 -6651 14804
rect -6685 14702 -6651 14736
rect -6685 14634 -6651 14668
rect -6685 14566 -6651 14600
rect -6685 14498 -6651 14532
rect -6685 14430 -6651 14464
rect -6685 14362 -6651 14396
rect -6685 14294 -6651 14328
rect -6685 14226 -6651 14260
rect -6685 14158 -6651 14192
rect -6685 14090 -6651 14124
rect -6685 14022 -6651 14056
rect -6685 13954 -6651 13988
rect -6685 13886 -6651 13920
rect -6685 13818 -6651 13852
rect -6685 13750 -6651 13784
rect -6685 13682 -6651 13716
rect -6685 13614 -6651 13648
rect -6685 13546 -6651 13580
rect -6685 13478 -6651 13512
rect -6685 13410 -6651 13444
rect -6685 13342 -6651 13376
rect -6685 13274 -6651 13308
rect -6685 13206 -6651 13240
rect -6685 13138 -6651 13172
rect -6685 13070 -6651 13104
rect -6685 13002 -6651 13036
rect -6685 12934 -6651 12968
rect -6685 12866 -6651 12900
rect -6427 14770 -6393 14804
rect -6427 14702 -6393 14736
rect -6427 14634 -6393 14668
rect -6427 14566 -6393 14600
rect -6427 14498 -6393 14532
rect -6427 14430 -6393 14464
rect -6427 14362 -6393 14396
rect -6427 14294 -6393 14328
rect -6427 14226 -6393 14260
rect -6427 14158 -6393 14192
rect -6427 14090 -6393 14124
rect -6427 14022 -6393 14056
rect -6427 13954 -6393 13988
rect -6427 13886 -6393 13920
rect -6427 13818 -6393 13852
rect -6427 13750 -6393 13784
rect -6427 13682 -6393 13716
rect -6427 13614 -6393 13648
rect -6427 13546 -6393 13580
rect -6427 13478 -6393 13512
rect -6427 13410 -6393 13444
rect -6427 13342 -6393 13376
rect -6427 13274 -6393 13308
rect -6427 13206 -6393 13240
rect -6427 13138 -6393 13172
rect -6427 13070 -6393 13104
rect -6427 13002 -6393 13036
rect -6427 12934 -6393 12968
rect -6427 12866 -6393 12900
rect -6169 14770 -6135 14804
rect -6169 14702 -6135 14736
rect -6169 14634 -6135 14668
rect -6169 14566 -6135 14600
rect -6169 14498 -6135 14532
rect -6169 14430 -6135 14464
rect -6169 14362 -6135 14396
rect -6169 14294 -6135 14328
rect -6169 14226 -6135 14260
rect -6169 14158 -6135 14192
rect -6169 14090 -6135 14124
rect -6169 14022 -6135 14056
rect -6169 13954 -6135 13988
rect -6169 13886 -6135 13920
rect -6169 13818 -6135 13852
rect -6169 13750 -6135 13784
rect -6169 13682 -6135 13716
rect -6169 13614 -6135 13648
rect -6169 13546 -6135 13580
rect -6169 13478 -6135 13512
rect -6169 13410 -6135 13444
rect -6169 13342 -6135 13376
rect -6169 13274 -6135 13308
rect -6169 13206 -6135 13240
rect -6169 13138 -6135 13172
rect -6169 13070 -6135 13104
rect -6169 13002 -6135 13036
rect -6169 12934 -6135 12968
rect -6169 12866 -6135 12900
rect -5911 14770 -5877 14804
rect -5911 14702 -5877 14736
rect -5911 14634 -5877 14668
rect -5911 14566 -5877 14600
rect -5911 14498 -5877 14532
rect -5911 14430 -5877 14464
rect -5911 14362 -5877 14396
rect -5911 14294 -5877 14328
rect -5911 14226 -5877 14260
rect -5911 14158 -5877 14192
rect -5911 14090 -5877 14124
rect -5911 14022 -5877 14056
rect -5911 13954 -5877 13988
rect -5911 13886 -5877 13920
rect -5911 13818 -5877 13852
rect -5911 13750 -5877 13784
rect -5911 13682 -5877 13716
rect -5911 13614 -5877 13648
rect -5911 13546 -5877 13580
rect -5911 13478 -5877 13512
rect -5911 13410 -5877 13444
rect -5911 13342 -5877 13376
rect -5911 13274 -5877 13308
rect -5911 13206 -5877 13240
rect -5911 13138 -5877 13172
rect -5911 13070 -5877 13104
rect -5911 13002 -5877 13036
rect -5911 12934 -5877 12968
rect -5911 12866 -5877 12900
rect -5653 14770 -5619 14804
rect -5653 14702 -5619 14736
rect -5653 14634 -5619 14668
rect -5653 14566 -5619 14600
rect -5653 14498 -5619 14532
rect -5653 14430 -5619 14464
rect -5653 14362 -5619 14396
rect -5653 14294 -5619 14328
rect -5653 14226 -5619 14260
rect -5653 14158 -5619 14192
rect -5653 14090 -5619 14124
rect -5653 14022 -5619 14056
rect -5653 13954 -5619 13988
rect -5653 13886 -5619 13920
rect -5653 13818 -5619 13852
rect -5653 13750 -5619 13784
rect -5653 13682 -5619 13716
rect -5653 13614 -5619 13648
rect -5653 13546 -5619 13580
rect -5653 13478 -5619 13512
rect -5653 13410 -5619 13444
rect -5653 13342 -5619 13376
rect -5653 13274 -5619 13308
rect -5653 13206 -5619 13240
rect -5653 13138 -5619 13172
rect -5653 13070 -5619 13104
rect -5653 13002 -5619 13036
rect -5653 12934 -5619 12968
rect -5653 12866 -5619 12900
rect -5395 14770 -5361 14804
rect -5395 14702 -5361 14736
rect -5395 14634 -5361 14668
rect -5395 14566 -5361 14600
rect -5395 14498 -5361 14532
rect -5395 14430 -5361 14464
rect -5395 14362 -5361 14396
rect -5395 14294 -5361 14328
rect -5395 14226 -5361 14260
rect -5395 14158 -5361 14192
rect -5395 14090 -5361 14124
rect -5395 14022 -5361 14056
rect -5395 13954 -5361 13988
rect -5395 13886 -5361 13920
rect -5395 13818 -5361 13852
rect -5395 13750 -5361 13784
rect -5395 13682 -5361 13716
rect -5395 13614 -5361 13648
rect -5395 13546 -5361 13580
rect -5395 13478 -5361 13512
rect -5395 13410 -5361 13444
rect -5395 13342 -5361 13376
rect -5395 13274 -5361 13308
rect -5395 13206 -5361 13240
rect -5395 13138 -5361 13172
rect -5395 13070 -5361 13104
rect -5395 13002 -5361 13036
rect -5395 12934 -5361 12968
rect -5395 12866 -5361 12900
rect -5137 14770 -5103 14804
rect -5137 14702 -5103 14736
rect -5137 14634 -5103 14668
rect -5137 14566 -5103 14600
rect -5137 14498 -5103 14532
rect -5137 14430 -5103 14464
rect -5137 14362 -5103 14396
rect -5137 14294 -5103 14328
rect -5137 14226 -5103 14260
rect -5137 14158 -5103 14192
rect -5137 14090 -5103 14124
rect -5137 14022 -5103 14056
rect -5137 13954 -5103 13988
rect -5137 13886 -5103 13920
rect -5137 13818 -5103 13852
rect -5137 13750 -5103 13784
rect -5137 13682 -5103 13716
rect -5137 13614 -5103 13648
rect -5137 13546 -5103 13580
rect -5137 13478 -5103 13512
rect -5137 13410 -5103 13444
rect -5137 13342 -5103 13376
rect -5137 13274 -5103 13308
rect -5137 13206 -5103 13240
rect -5137 13138 -5103 13172
rect -5137 13070 -5103 13104
rect -5137 13002 -5103 13036
rect -5137 12934 -5103 12968
rect -5137 12866 -5103 12900
rect -4879 14770 -4845 14804
rect -4879 14702 -4845 14736
rect -4879 14634 -4845 14668
rect -4879 14566 -4845 14600
rect -4879 14498 -4845 14532
rect -4879 14430 -4845 14464
rect -4879 14362 -4845 14396
rect -4879 14294 -4845 14328
rect -4879 14226 -4845 14260
rect -4879 14158 -4845 14192
rect -4879 14090 -4845 14124
rect -4879 14022 -4845 14056
rect -4879 13954 -4845 13988
rect -4879 13886 -4845 13920
rect -4879 13818 -4845 13852
rect -4879 13750 -4845 13784
rect -4879 13682 -4845 13716
rect -4879 13614 -4845 13648
rect -4879 13546 -4845 13580
rect -4879 13478 -4845 13512
rect -4879 13410 -4845 13444
rect -4879 13342 -4845 13376
rect -4879 13274 -4845 13308
rect -4879 13206 -4845 13240
rect -4879 13138 -4845 13172
rect -4879 13070 -4845 13104
rect -4879 13002 -4845 13036
rect -4879 12934 -4845 12968
rect -4879 12866 -4845 12900
rect -8815 11089 -8781 11123
rect -8815 11021 -8781 11055
rect -8815 10953 -8781 10987
rect -8815 10885 -8781 10919
rect -8815 10817 -8781 10851
rect -8815 10749 -8781 10783
rect -8815 10681 -8781 10715
rect -8815 10613 -8781 10647
rect -8815 10545 -8781 10579
rect -8815 10477 -8781 10511
rect -8815 10409 -8781 10443
rect -8815 10341 -8781 10375
rect -8815 10273 -8781 10307
rect -8815 10205 -8781 10239
rect -8557 11089 -8523 11123
rect -8557 11021 -8523 11055
rect -8557 10953 -8523 10987
rect -8557 10885 -8523 10919
rect -8557 10817 -8523 10851
rect -8557 10749 -8523 10783
rect -8557 10681 -8523 10715
rect -8557 10613 -8523 10647
rect -8557 10545 -8523 10579
rect -8557 10477 -8523 10511
rect -8557 10409 -8523 10443
rect -8557 10341 -8523 10375
rect -8557 10273 -8523 10307
rect -8557 10205 -8523 10239
rect -8299 11089 -8265 11123
rect -8299 11021 -8265 11055
rect -8299 10953 -8265 10987
rect -8299 10885 -8265 10919
rect -8299 10817 -8265 10851
rect -8299 10749 -8265 10783
rect -8299 10681 -8265 10715
rect -8299 10613 -8265 10647
rect -8299 10545 -8265 10579
rect -8299 10477 -8265 10511
rect -8299 10409 -8265 10443
rect -8299 10341 -8265 10375
rect -8299 10273 -8265 10307
rect -8299 10205 -8265 10239
rect -8041 11089 -8007 11123
rect -8041 11021 -8007 11055
rect -8041 10953 -8007 10987
rect -8041 10885 -8007 10919
rect -8041 10817 -8007 10851
rect -8041 10749 -8007 10783
rect -8041 10681 -8007 10715
rect -8041 10613 -8007 10647
rect -8041 10545 -8007 10579
rect -8041 10477 -8007 10511
rect -8041 10409 -8007 10443
rect -8041 10341 -8007 10375
rect -8041 10273 -8007 10307
rect -8041 10205 -8007 10239
rect -7783 11089 -7749 11123
rect -7783 11021 -7749 11055
rect -7783 10953 -7749 10987
rect -7783 10885 -7749 10919
rect -7783 10817 -7749 10851
rect -7783 10749 -7749 10783
rect -7783 10681 -7749 10715
rect -7783 10613 -7749 10647
rect -7783 10545 -7749 10579
rect -7783 10477 -7749 10511
rect -7783 10409 -7749 10443
rect -7783 10341 -7749 10375
rect -7783 10273 -7749 10307
rect -7783 10205 -7749 10239
rect -7525 11089 -7491 11123
rect -7525 11021 -7491 11055
rect -7525 10953 -7491 10987
rect -7525 10885 -7491 10919
rect -7525 10817 -7491 10851
rect -7525 10749 -7491 10783
rect -7525 10681 -7491 10715
rect -7525 10613 -7491 10647
rect -7525 10545 -7491 10579
rect -7525 10477 -7491 10511
rect -7525 10409 -7491 10443
rect -7525 10341 -7491 10375
rect -7525 10273 -7491 10307
rect -7525 10205 -7491 10239
rect -7267 11089 -7233 11123
rect -7267 11021 -7233 11055
rect -7267 10953 -7233 10987
rect -7267 10885 -7233 10919
rect -7267 10817 -7233 10851
rect -7267 10749 -7233 10783
rect -7267 10681 -7233 10715
rect -7267 10613 -7233 10647
rect -7267 10545 -7233 10579
rect -7267 10477 -7233 10511
rect -7267 10409 -7233 10443
rect -7267 10341 -7233 10375
rect -7267 10273 -7233 10307
rect -7267 10205 -7233 10239
rect -7009 11089 -6975 11123
rect -7009 11021 -6975 11055
rect -7009 10953 -6975 10987
rect -7009 10885 -6975 10919
rect -7009 10817 -6975 10851
rect -7009 10749 -6975 10783
rect -7009 10681 -6975 10715
rect -7009 10613 -6975 10647
rect -7009 10545 -6975 10579
rect -7009 10477 -6975 10511
rect -7009 10409 -6975 10443
rect -7009 10341 -6975 10375
rect -7009 10273 -6975 10307
rect -7009 10205 -6975 10239
rect -6751 11089 -6717 11123
rect -6751 11021 -6717 11055
rect -6751 10953 -6717 10987
rect -6751 10885 -6717 10919
rect -6751 10817 -6717 10851
rect -6751 10749 -6717 10783
rect -6751 10681 -6717 10715
rect -6751 10613 -6717 10647
rect -6751 10545 -6717 10579
rect -6751 10477 -6717 10511
rect -6751 10409 -6717 10443
rect -6751 10341 -6717 10375
rect -6751 10273 -6717 10307
rect -6751 10205 -6717 10239
rect -6493 11089 -6459 11123
rect -6493 11021 -6459 11055
rect -6493 10953 -6459 10987
rect -6493 10885 -6459 10919
rect -6493 10817 -6459 10851
rect -6493 10749 -6459 10783
rect -6493 10681 -6459 10715
rect -6493 10613 -6459 10647
rect -6493 10545 -6459 10579
rect -6493 10477 -6459 10511
rect -6493 10409 -6459 10443
rect -6493 10341 -6459 10375
rect -6493 10273 -6459 10307
rect -6493 10205 -6459 10239
rect -6235 11089 -6201 11123
rect -6235 11021 -6201 11055
rect -6235 10953 -6201 10987
rect -6235 10885 -6201 10919
rect -6235 10817 -6201 10851
rect -6235 10749 -6201 10783
rect -6235 10681 -6201 10715
rect -6235 10613 -6201 10647
rect -6235 10545 -6201 10579
rect -6235 10477 -6201 10511
rect -6235 10409 -6201 10443
rect -6235 10341 -6201 10375
rect -6235 10273 -6201 10307
rect -6235 10205 -6201 10239
rect -5977 11089 -5943 11123
rect -5977 11021 -5943 11055
rect -5977 10953 -5943 10987
rect -5977 10885 -5943 10919
rect -5977 10817 -5943 10851
rect -5977 10749 -5943 10783
rect -5977 10681 -5943 10715
rect -5977 10613 -5943 10647
rect -5977 10545 -5943 10579
rect -5977 10477 -5943 10511
rect -5977 10409 -5943 10443
rect -5977 10341 -5943 10375
rect -5977 10273 -5943 10307
rect -5977 10205 -5943 10239
rect -5719 11089 -5685 11123
rect -5719 11021 -5685 11055
rect -5719 10953 -5685 10987
rect -5719 10885 -5685 10919
rect -5719 10817 -5685 10851
rect -5719 10749 -5685 10783
rect -5719 10681 -5685 10715
rect -5719 10613 -5685 10647
rect -5719 10545 -5685 10579
rect -5719 10477 -5685 10511
rect -5719 10409 -5685 10443
rect -5719 10341 -5685 10375
rect -5719 10273 -5685 10307
rect -5719 10205 -5685 10239
rect -5461 11089 -5427 11123
rect -5461 11021 -5427 11055
rect -5461 10953 -5427 10987
rect -5461 10885 -5427 10919
rect -5461 10817 -5427 10851
rect -5461 10749 -5427 10783
rect -5461 10681 -5427 10715
rect -5461 10613 -5427 10647
rect -5461 10545 -5427 10579
rect -5461 10477 -5427 10511
rect -5461 10409 -5427 10443
rect -5461 10341 -5427 10375
rect -5461 10273 -5427 10307
rect -5461 10205 -5427 10239
rect -5203 11089 -5169 11123
rect -5203 11021 -5169 11055
rect -5203 10953 -5169 10987
rect -5203 10885 -5169 10919
rect -5203 10817 -5169 10851
rect -5203 10749 -5169 10783
rect -5203 10681 -5169 10715
rect -5203 10613 -5169 10647
rect -5203 10545 -5169 10579
rect -5203 10477 -5169 10511
rect -5203 10409 -5169 10443
rect -5203 10341 -5169 10375
rect -5203 10273 -5169 10307
rect -5203 10205 -5169 10239
rect -4945 11089 -4911 11123
rect -4945 11021 -4911 11055
rect -4945 10953 -4911 10987
rect -4945 10885 -4911 10919
rect -4945 10817 -4911 10851
rect -4945 10749 -4911 10783
rect -4945 10681 -4911 10715
rect -4945 10613 -4911 10647
rect -4945 10545 -4911 10579
rect -4945 10477 -4911 10511
rect -4945 10409 -4911 10443
rect -4945 10341 -4911 10375
rect -4945 10273 -4911 10307
rect -4945 10205 -4911 10239
rect -4687 11089 -4653 11123
rect -4687 11021 -4653 11055
rect -4687 10953 -4653 10987
rect -4687 10885 -4653 10919
rect -4687 10817 -4653 10851
rect -4687 10749 -4653 10783
rect -4687 10681 -4653 10715
rect -4687 10613 -4653 10647
rect -4687 10545 -4653 10579
rect -4687 10477 -4653 10511
rect -4687 10409 -4653 10443
rect -4687 10341 -4653 10375
rect -4687 10273 -4653 10307
rect -4687 10205 -4653 10239
rect -4429 11089 -4395 11123
rect -4429 11021 -4395 11055
rect -4429 10953 -4395 10987
rect -4429 10885 -4395 10919
rect -4429 10817 -4395 10851
rect -4429 10749 -4395 10783
rect -4429 10681 -4395 10715
rect -4429 10613 -4395 10647
rect -4429 10545 -4395 10579
rect -4429 10477 -4395 10511
rect -4429 10409 -4395 10443
rect -4429 10341 -4395 10375
rect -4429 10273 -4395 10307
rect -4429 10205 -4395 10239
rect -4171 11089 -4137 11123
rect -4171 11021 -4137 11055
rect -4171 10953 -4137 10987
rect -4171 10885 -4137 10919
rect -4171 10817 -4137 10851
rect -4171 10749 -4137 10783
rect -4171 10681 -4137 10715
rect -4171 10613 -4137 10647
rect -4171 10545 -4137 10579
rect -4171 10477 -4137 10511
rect -4171 10409 -4137 10443
rect -4171 10341 -4137 10375
rect -4171 10273 -4137 10307
rect -4171 10205 -4137 10239
rect -3913 11089 -3879 11123
rect -3913 11021 -3879 11055
rect -3913 10953 -3879 10987
rect -3913 10885 -3879 10919
rect -3913 10817 -3879 10851
rect -3913 10749 -3879 10783
rect -3913 10681 -3879 10715
rect -3913 10613 -3879 10647
rect -3913 10545 -3879 10579
rect -3913 10477 -3879 10511
rect -3913 10409 -3879 10443
rect -3913 10341 -3879 10375
rect -3913 10273 -3879 10307
rect -3913 10205 -3879 10239
rect -3655 11089 -3621 11123
rect -3655 11021 -3621 11055
rect -3655 10953 -3621 10987
rect -3655 10885 -3621 10919
rect -3655 10817 -3621 10851
rect -3655 10749 -3621 10783
rect -3655 10681 -3621 10715
rect -3655 10613 -3621 10647
rect -3655 10545 -3621 10579
rect -3655 10477 -3621 10511
rect -3655 10409 -3621 10443
rect -3655 10341 -3621 10375
rect -3655 10273 -3621 10307
rect -3655 10205 -3621 10239
rect -7780 9724 -7746 9758
rect -7780 9656 -7746 9690
rect -7780 9588 -7746 9622
rect -7780 9520 -7746 9554
rect -7780 9452 -7746 9486
rect -7780 9384 -7746 9418
rect -7780 9316 -7746 9350
rect -7780 9248 -7746 9282
rect -7780 9180 -7746 9214
rect -7780 9112 -7746 9146
rect -7780 9044 -7746 9078
rect -7780 8976 -7746 9010
rect -7780 8908 -7746 8942
rect -7780 8840 -7746 8874
rect -7522 9724 -7488 9758
rect -7522 9656 -7488 9690
rect -7522 9588 -7488 9622
rect -7522 9520 -7488 9554
rect -7522 9452 -7488 9486
rect -7522 9384 -7488 9418
rect -7522 9316 -7488 9350
rect -7522 9248 -7488 9282
rect -7522 9180 -7488 9214
rect -7522 9112 -7488 9146
rect -7522 9044 -7488 9078
rect -7522 8976 -7488 9010
rect -7522 8908 -7488 8942
rect -7522 8840 -7488 8874
rect -7314 9724 -7280 9758
rect -7314 9656 -7280 9690
rect -7314 9588 -7280 9622
rect -7314 9520 -7280 9554
rect -7314 9452 -7280 9486
rect -7314 9384 -7280 9418
rect -7314 9316 -7280 9350
rect -7314 9248 -7280 9282
rect -7314 9180 -7280 9214
rect -7314 9112 -7280 9146
rect -7314 9044 -7280 9078
rect -7314 8976 -7280 9010
rect -7314 8908 -7280 8942
rect -7314 8840 -7280 8874
rect -7056 9724 -7022 9758
rect -7056 9656 -7022 9690
rect -7056 9588 -7022 9622
rect -7056 9520 -7022 9554
rect -7056 9452 -7022 9486
rect -7056 9384 -7022 9418
rect -7056 9316 -7022 9350
rect -7056 9248 -7022 9282
rect -7056 9180 -7022 9214
rect -7056 9112 -7022 9146
rect -7056 9044 -7022 9078
rect -7056 8976 -7022 9010
rect -7056 8908 -7022 8942
rect -7056 8840 -7022 8874
rect -6798 9724 -6764 9758
rect -6798 9656 -6764 9690
rect -6798 9588 -6764 9622
rect -6798 9520 -6764 9554
rect -6798 9452 -6764 9486
rect -6798 9384 -6764 9418
rect -6798 9316 -6764 9350
rect -6798 9248 -6764 9282
rect -6798 9180 -6764 9214
rect -6798 9112 -6764 9146
rect -6798 9044 -6764 9078
rect -6798 8976 -6764 9010
rect -6798 8908 -6764 8942
rect -6798 8840 -6764 8874
rect -6540 9724 -6506 9758
rect -6540 9656 -6506 9690
rect -6540 9588 -6506 9622
rect -6540 9520 -6506 9554
rect -6540 9452 -6506 9486
rect -6540 9384 -6506 9418
rect -6540 9316 -6506 9350
rect -6540 9248 -6506 9282
rect -6540 9180 -6506 9214
rect -6540 9112 -6506 9146
rect -6540 9044 -6506 9078
rect -6540 8976 -6506 9010
rect -6540 8908 -6506 8942
rect -6540 8840 -6506 8874
rect -6282 9724 -6248 9758
rect -6282 9656 -6248 9690
rect -6282 9588 -6248 9622
rect -6282 9520 -6248 9554
rect -6282 9452 -6248 9486
rect -6282 9384 -6248 9418
rect -6282 9316 -6248 9350
rect -6282 9248 -6248 9282
rect -6282 9180 -6248 9214
rect -6282 9112 -6248 9146
rect -6282 9044 -6248 9078
rect -6282 8976 -6248 9010
rect -6282 8908 -6248 8942
rect -6282 8840 -6248 8874
rect -6024 9724 -5990 9758
rect -6024 9656 -5990 9690
rect -6024 9588 -5990 9622
rect -6024 9520 -5990 9554
rect -6024 9452 -5990 9486
rect -6024 9384 -5990 9418
rect -6024 9316 -5990 9350
rect -6024 9248 -5990 9282
rect -6024 9180 -5990 9214
rect -6024 9112 -5990 9146
rect -6024 9044 -5990 9078
rect -6024 8976 -5990 9010
rect -6024 8908 -5990 8942
rect -6024 8840 -5990 8874
rect -5766 9724 -5732 9758
rect -5766 9656 -5732 9690
rect -5766 9588 -5732 9622
rect -5766 9520 -5732 9554
rect -5766 9452 -5732 9486
rect -5766 9384 -5732 9418
rect -5766 9316 -5732 9350
rect -5766 9248 -5732 9282
rect -5766 9180 -5732 9214
rect -5766 9112 -5732 9146
rect -5766 9044 -5732 9078
rect -5766 8976 -5732 9010
rect -5766 8908 -5732 8942
rect -5766 8840 -5732 8874
rect -5508 9724 -5474 9758
rect -5508 9656 -5474 9690
rect -5508 9588 -5474 9622
rect -5508 9520 -5474 9554
rect -5508 9452 -5474 9486
rect -5508 9384 -5474 9418
rect -5508 9316 -5474 9350
rect -5508 9248 -5474 9282
rect -5508 9180 -5474 9214
rect -5508 9112 -5474 9146
rect -5508 9044 -5474 9078
rect -5508 8976 -5474 9010
rect -5508 8908 -5474 8942
rect -5508 8840 -5474 8874
rect -5250 9724 -5216 9758
rect -5250 9656 -5216 9690
rect -5250 9588 -5216 9622
rect -5250 9520 -5216 9554
rect -5250 9452 -5216 9486
rect -5250 9384 -5216 9418
rect -5250 9316 -5216 9350
rect -5250 9248 -5216 9282
rect -5250 9180 -5216 9214
rect -5250 9112 -5216 9146
rect -5250 9044 -5216 9078
rect -5250 8976 -5216 9010
rect -5250 8908 -5216 8942
rect -5250 8840 -5216 8874
rect -4992 9724 -4958 9758
rect -4992 9656 -4958 9690
rect -4992 9588 -4958 9622
rect -4992 9520 -4958 9554
rect -4992 9452 -4958 9486
rect -4992 9384 -4958 9418
rect -4992 9316 -4958 9350
rect -4992 9248 -4958 9282
rect -4992 9180 -4958 9214
rect -4992 9112 -4958 9146
rect -4992 9044 -4958 9078
rect -4992 8976 -4958 9010
rect -4992 8908 -4958 8942
rect -4992 8840 -4958 8874
rect -4734 9724 -4700 9758
rect -4734 9656 -4700 9690
rect -4734 9588 -4700 9622
rect -4734 9520 -4700 9554
rect -4734 9452 -4700 9486
rect -4734 9384 -4700 9418
rect -4734 9316 -4700 9350
rect -4734 9248 -4700 9282
rect -4734 9180 -4700 9214
rect -4734 9112 -4700 9146
rect -4734 9044 -4700 9078
rect -4734 8976 -4700 9010
rect -4734 8908 -4700 8942
rect -4734 8840 -4700 8874
rect -7780 7473 -7746 7507
rect -7780 7405 -7746 7439
rect -7780 7337 -7746 7371
rect -7780 7269 -7746 7303
rect -7780 7201 -7746 7235
rect -7780 7133 -7746 7167
rect -7780 7065 -7746 7099
rect -7780 6997 -7746 7031
rect -7780 6929 -7746 6963
rect -7780 6861 -7746 6895
rect -7780 6793 -7746 6827
rect -7780 6725 -7746 6759
rect -7780 6657 -7746 6691
rect -7780 6589 -7746 6623
rect -7780 6521 -7746 6555
rect -7780 6453 -7746 6487
rect -7780 6385 -7746 6419
rect -7780 6317 -7746 6351
rect -7780 6249 -7746 6283
rect -7780 6181 -7746 6215
rect -7780 6113 -7746 6147
rect -7780 6045 -7746 6079
rect -7780 5977 -7746 6011
rect -7780 5909 -7746 5943
rect -7780 5841 -7746 5875
rect -7780 5773 -7746 5807
rect -7780 5705 -7746 5739
rect -7780 5637 -7746 5671
rect -7780 5569 -7746 5603
rect -7522 7473 -7488 7507
rect -7522 7405 -7488 7439
rect -7522 7337 -7488 7371
rect -7522 7269 -7488 7303
rect -7522 7201 -7488 7235
rect -7522 7133 -7488 7167
rect -7522 7065 -7488 7099
rect -7522 6997 -7488 7031
rect -7522 6929 -7488 6963
rect -7522 6861 -7488 6895
rect -7522 6793 -7488 6827
rect -7522 6725 -7488 6759
rect -7522 6657 -7488 6691
rect -7522 6589 -7488 6623
rect -7522 6521 -7488 6555
rect -7522 6453 -7488 6487
rect -7522 6385 -7488 6419
rect -7522 6317 -7488 6351
rect -7522 6249 -7488 6283
rect -7522 6181 -7488 6215
rect -7522 6113 -7488 6147
rect -7522 6045 -7488 6079
rect -7522 5977 -7488 6011
rect -7522 5909 -7488 5943
rect -7522 5841 -7488 5875
rect -7522 5773 -7488 5807
rect -7522 5705 -7488 5739
rect -7522 5637 -7488 5671
rect -7522 5569 -7488 5603
rect -7264 7473 -7230 7507
rect -7264 7405 -7230 7439
rect -7264 7337 -7230 7371
rect -7264 7269 -7230 7303
rect -7264 7201 -7230 7235
rect -7264 7133 -7230 7167
rect -7264 7065 -7230 7099
rect -7264 6997 -7230 7031
rect -7264 6929 -7230 6963
rect -7264 6861 -7230 6895
rect -7264 6793 -7230 6827
rect -7264 6725 -7230 6759
rect -7264 6657 -7230 6691
rect -7264 6589 -7230 6623
rect -7264 6521 -7230 6555
rect -7264 6453 -7230 6487
rect -7264 6385 -7230 6419
rect -7264 6317 -7230 6351
rect -7264 6249 -7230 6283
rect -7264 6181 -7230 6215
rect -7264 6113 -7230 6147
rect -7264 6045 -7230 6079
rect -7264 5977 -7230 6011
rect -7264 5909 -7230 5943
rect -7264 5841 -7230 5875
rect -7264 5773 -7230 5807
rect -7264 5705 -7230 5739
rect -7264 5637 -7230 5671
rect -7264 5569 -7230 5603
rect -7006 7473 -6972 7507
rect -7006 7405 -6972 7439
rect -7006 7337 -6972 7371
rect -7006 7269 -6972 7303
rect -7006 7201 -6972 7235
rect -7006 7133 -6972 7167
rect -7006 7065 -6972 7099
rect -7006 6997 -6972 7031
rect -7006 6929 -6972 6963
rect -7006 6861 -6972 6895
rect -7006 6793 -6972 6827
rect -7006 6725 -6972 6759
rect -7006 6657 -6972 6691
rect -7006 6589 -6972 6623
rect -7006 6521 -6972 6555
rect -7006 6453 -6972 6487
rect -7006 6385 -6972 6419
rect -7006 6317 -6972 6351
rect -7006 6249 -6972 6283
rect -7006 6181 -6972 6215
rect -7006 6113 -6972 6147
rect -7006 6045 -6972 6079
rect -7006 5977 -6972 6011
rect -7006 5909 -6972 5943
rect -7006 5841 -6972 5875
rect -7006 5773 -6972 5807
rect -7006 5705 -6972 5739
rect -7006 5637 -6972 5671
rect -7006 5569 -6972 5603
rect -6748 7473 -6714 7507
rect -6748 7405 -6714 7439
rect -6748 7337 -6714 7371
rect -6748 7269 -6714 7303
rect -6748 7201 -6714 7235
rect -6748 7133 -6714 7167
rect -6748 7065 -6714 7099
rect -6748 6997 -6714 7031
rect -6748 6929 -6714 6963
rect -6748 6861 -6714 6895
rect -6748 6793 -6714 6827
rect -6748 6725 -6714 6759
rect -6748 6657 -6714 6691
rect -6748 6589 -6714 6623
rect -6748 6521 -6714 6555
rect -6748 6453 -6714 6487
rect -6748 6385 -6714 6419
rect -6748 6317 -6714 6351
rect -6748 6249 -6714 6283
rect -6748 6181 -6714 6215
rect -6748 6113 -6714 6147
rect -6748 6045 -6714 6079
rect -6748 5977 -6714 6011
rect -6748 5909 -6714 5943
rect -6748 5841 -6714 5875
rect -6748 5773 -6714 5807
rect -6748 5705 -6714 5739
rect -6748 5637 -6714 5671
rect -6748 5569 -6714 5603
rect -6490 7473 -6456 7507
rect -6490 7405 -6456 7439
rect -6490 7337 -6456 7371
rect -6490 7269 -6456 7303
rect -6490 7201 -6456 7235
rect -6490 7133 -6456 7167
rect -6490 7065 -6456 7099
rect -6490 6997 -6456 7031
rect -6490 6929 -6456 6963
rect -6490 6861 -6456 6895
rect -6490 6793 -6456 6827
rect -6490 6725 -6456 6759
rect -6490 6657 -6456 6691
rect -6490 6589 -6456 6623
rect -6490 6521 -6456 6555
rect -6490 6453 -6456 6487
rect -6490 6385 -6456 6419
rect -6490 6317 -6456 6351
rect -6490 6249 -6456 6283
rect -6490 6181 -6456 6215
rect -6490 6113 -6456 6147
rect -6490 6045 -6456 6079
rect -6490 5977 -6456 6011
rect -6490 5909 -6456 5943
rect -6490 5841 -6456 5875
rect -6490 5773 -6456 5807
rect -6490 5705 -6456 5739
rect -6490 5637 -6456 5671
rect -6490 5569 -6456 5603
rect -6232 7473 -6198 7507
rect -6232 7405 -6198 7439
rect -6232 7337 -6198 7371
rect -6232 7269 -6198 7303
rect -6232 7201 -6198 7235
rect -6232 7133 -6198 7167
rect -6232 7065 -6198 7099
rect -6232 6997 -6198 7031
rect -6232 6929 -6198 6963
rect -6232 6861 -6198 6895
rect -6232 6793 -6198 6827
rect -6232 6725 -6198 6759
rect -6232 6657 -6198 6691
rect -6232 6589 -6198 6623
rect -6232 6521 -6198 6555
rect -6232 6453 -6198 6487
rect -6232 6385 -6198 6419
rect -6232 6317 -6198 6351
rect -6232 6249 -6198 6283
rect -6232 6181 -6198 6215
rect -6232 6113 -6198 6147
rect -6232 6045 -6198 6079
rect -6232 5977 -6198 6011
rect -6232 5909 -6198 5943
rect -6232 5841 -6198 5875
rect -6232 5773 -6198 5807
rect -6232 5705 -6198 5739
rect -6232 5637 -6198 5671
rect -6232 5569 -6198 5603
rect -5974 7473 -5940 7507
rect -5974 7405 -5940 7439
rect -5974 7337 -5940 7371
rect -5974 7269 -5940 7303
rect -5974 7201 -5940 7235
rect -5974 7133 -5940 7167
rect -5974 7065 -5940 7099
rect -5974 6997 -5940 7031
rect -5974 6929 -5940 6963
rect -5974 6861 -5940 6895
rect -5974 6793 -5940 6827
rect -5974 6725 -5940 6759
rect -5974 6657 -5940 6691
rect -5974 6589 -5940 6623
rect -5974 6521 -5940 6555
rect -5974 6453 -5940 6487
rect -5974 6385 -5940 6419
rect -5974 6317 -5940 6351
rect -5974 6249 -5940 6283
rect -5974 6181 -5940 6215
rect -5974 6113 -5940 6147
rect -5974 6045 -5940 6079
rect -5974 5977 -5940 6011
rect -5974 5909 -5940 5943
rect -5974 5841 -5940 5875
rect -5974 5773 -5940 5807
rect -5974 5705 -5940 5739
rect -5974 5637 -5940 5671
rect -5974 5569 -5940 5603
rect -5716 7473 -5682 7507
rect -5716 7405 -5682 7439
rect -5716 7337 -5682 7371
rect -5716 7269 -5682 7303
rect -5716 7201 -5682 7235
rect -5716 7133 -5682 7167
rect -5716 7065 -5682 7099
rect -5716 6997 -5682 7031
rect -5716 6929 -5682 6963
rect -5716 6861 -5682 6895
rect -5716 6793 -5682 6827
rect -5716 6725 -5682 6759
rect -5716 6657 -5682 6691
rect -5716 6589 -5682 6623
rect -5716 6521 -5682 6555
rect -5716 6453 -5682 6487
rect -5716 6385 -5682 6419
rect -5716 6317 -5682 6351
rect -5716 6249 -5682 6283
rect -5716 6181 -5682 6215
rect -5716 6113 -5682 6147
rect -5716 6045 -5682 6079
rect -5716 5977 -5682 6011
rect -5716 5909 -5682 5943
rect -5716 5841 -5682 5875
rect -5716 5773 -5682 5807
rect -5716 5705 -5682 5739
rect -5716 5637 -5682 5671
rect -5716 5569 -5682 5603
rect -5458 7473 -5424 7507
rect -5458 7405 -5424 7439
rect -5458 7337 -5424 7371
rect -5458 7269 -5424 7303
rect -5458 7201 -5424 7235
rect -5458 7133 -5424 7167
rect -5458 7065 -5424 7099
rect -5458 6997 -5424 7031
rect -5458 6929 -5424 6963
rect -5458 6861 -5424 6895
rect -5458 6793 -5424 6827
rect -5458 6725 -5424 6759
rect -5458 6657 -5424 6691
rect -5458 6589 -5424 6623
rect -5458 6521 -5424 6555
rect -5458 6453 -5424 6487
rect -5458 6385 -5424 6419
rect -5458 6317 -5424 6351
rect -5458 6249 -5424 6283
rect -5458 6181 -5424 6215
rect -5458 6113 -5424 6147
rect -5458 6045 -5424 6079
rect -5458 5977 -5424 6011
rect -5458 5909 -5424 5943
rect -5458 5841 -5424 5875
rect -5458 5773 -5424 5807
rect -5458 5705 -5424 5739
rect -5458 5637 -5424 5671
rect -5458 5569 -5424 5603
rect -5200 7473 -5166 7507
rect -5200 7405 -5166 7439
rect -5200 7337 -5166 7371
rect -5200 7269 -5166 7303
rect -5200 7201 -5166 7235
rect -5200 7133 -5166 7167
rect -5200 7065 -5166 7099
rect -5200 6997 -5166 7031
rect -5200 6929 -5166 6963
rect -5200 6861 -5166 6895
rect -5200 6793 -5166 6827
rect -5200 6725 -5166 6759
rect -5200 6657 -5166 6691
rect -5200 6589 -5166 6623
rect -5200 6521 -5166 6555
rect -5200 6453 -5166 6487
rect -5200 6385 -5166 6419
rect -5200 6317 -5166 6351
rect -5200 6249 -5166 6283
rect -5200 6181 -5166 6215
rect -5200 6113 -5166 6147
rect -5200 6045 -5166 6079
rect -5200 5977 -5166 6011
rect -5200 5909 -5166 5943
rect -5200 5841 -5166 5875
rect -5200 5773 -5166 5807
rect -5200 5705 -5166 5739
rect -5200 5637 -5166 5671
rect -5200 5569 -5166 5603
rect -4942 7473 -4908 7507
rect -4942 7405 -4908 7439
rect -4942 7337 -4908 7371
rect -4942 7269 -4908 7303
rect -4942 7201 -4908 7235
rect -4942 7133 -4908 7167
rect -4942 7065 -4908 7099
rect -4942 6997 -4908 7031
rect -4942 6929 -4908 6963
rect -4942 6861 -4908 6895
rect -4942 6793 -4908 6827
rect -4942 6725 -4908 6759
rect -4942 6657 -4908 6691
rect -4942 6589 -4908 6623
rect -4942 6521 -4908 6555
rect -4942 6453 -4908 6487
rect -4942 6385 -4908 6419
rect -4942 6317 -4908 6351
rect -4942 6249 -4908 6283
rect -4942 6181 -4908 6215
rect -4942 6113 -4908 6147
rect -4942 6045 -4908 6079
rect -4942 5977 -4908 6011
rect -4942 5909 -4908 5943
rect -4942 5841 -4908 5875
rect -4942 5773 -4908 5807
rect -4942 5705 -4908 5739
rect -4942 5637 -4908 5671
rect -4942 5569 -4908 5603
rect -4684 7473 -4650 7507
rect -4684 7405 -4650 7439
rect -4684 7337 -4650 7371
rect -4684 7269 -4650 7303
rect -4684 7201 -4650 7235
rect -4684 7133 -4650 7167
rect -4684 7065 -4650 7099
rect -4684 6997 -4650 7031
rect -4684 6929 -4650 6963
rect -4684 6861 -4650 6895
rect -4684 6793 -4650 6827
rect -4684 6725 -4650 6759
rect -4684 6657 -4650 6691
rect -4684 6589 -4650 6623
rect -4684 6521 -4650 6555
rect -4684 6453 -4650 6487
rect -4684 6385 -4650 6419
rect -4684 6317 -4650 6351
rect -4684 6249 -4650 6283
rect -4684 6181 -4650 6215
rect -4684 6113 -4650 6147
rect -4684 6045 -4650 6079
rect -4684 5977 -4650 6011
rect -4684 5909 -4650 5943
rect -4684 5841 -4650 5875
rect -4684 5773 -4650 5807
rect -4684 5705 -4650 5739
rect -4684 5637 -4650 5671
rect -4684 5569 -4650 5603
rect -4426 7473 -4392 7507
rect -4426 7405 -4392 7439
rect -4426 7337 -4392 7371
rect -4426 7269 -4392 7303
rect -4426 7201 -4392 7235
rect -4426 7133 -4392 7167
rect -4426 7065 -4392 7099
rect -4426 6997 -4392 7031
rect -4426 6929 -4392 6963
rect -4426 6861 -4392 6895
rect -4426 6793 -4392 6827
rect -4426 6725 -4392 6759
rect -4426 6657 -4392 6691
rect -4426 6589 -4392 6623
rect -4426 6521 -4392 6555
rect -4426 6453 -4392 6487
rect -4426 6385 -4392 6419
rect -4426 6317 -4392 6351
rect -4426 6249 -4392 6283
rect -4426 6181 -4392 6215
rect -4426 6113 -4392 6147
rect -4426 6045 -4392 6079
rect -4426 5977 -4392 6011
rect -4426 5909 -4392 5943
rect -4426 5841 -4392 5875
rect -4426 5773 -4392 5807
rect -4426 5705 -4392 5739
rect -4426 5637 -4392 5671
rect -4426 5569 -4392 5603
rect -4168 7473 -4134 7507
rect -4168 7405 -4134 7439
rect -4168 7337 -4134 7371
rect -4168 7269 -4134 7303
rect -4168 7201 -4134 7235
rect -4168 7133 -4134 7167
rect -4168 7065 -4134 7099
rect -4168 6997 -4134 7031
rect -4168 6929 -4134 6963
rect -4168 6861 -4134 6895
rect -4168 6793 -4134 6827
rect -4168 6725 -4134 6759
rect -4168 6657 -4134 6691
rect -4168 6589 -4134 6623
rect -4168 6521 -4134 6555
rect -4168 6453 -4134 6487
rect -4168 6385 -4134 6419
rect -4168 6317 -4134 6351
rect -4168 6249 -4134 6283
rect -4168 6181 -4134 6215
rect -4168 6113 -4134 6147
rect -4168 6045 -4134 6079
rect -4168 5977 -4134 6011
rect -4168 5909 -4134 5943
rect -4168 5841 -4134 5875
rect -4168 5773 -4134 5807
rect -4168 5705 -4134 5739
rect -4168 5637 -4134 5671
rect -4168 5569 -4134 5603
rect -3910 7473 -3876 7507
rect -3910 7405 -3876 7439
rect -3910 7337 -3876 7371
rect -3910 7269 -3876 7303
rect -3910 7201 -3876 7235
rect -3910 7133 -3876 7167
rect -3910 7065 -3876 7099
rect -3910 6997 -3876 7031
rect -3910 6929 -3876 6963
rect -3910 6861 -3876 6895
rect -3910 6793 -3876 6827
rect -3910 6725 -3876 6759
rect -3910 6657 -3876 6691
rect -3910 6589 -3876 6623
rect -3910 6521 -3876 6555
rect -3910 6453 -3876 6487
rect -3910 6385 -3876 6419
rect -3910 6317 -3876 6351
rect -3910 6249 -3876 6283
rect -3910 6181 -3876 6215
rect -3910 6113 -3876 6147
rect -3910 6045 -3876 6079
rect -3910 5977 -3876 6011
rect -3910 5909 -3876 5943
rect -3910 5841 -3876 5875
rect -3910 5773 -3876 5807
rect -3910 5705 -3876 5739
rect -3910 5637 -3876 5671
rect -3910 5569 -3876 5603
rect -3652 7473 -3618 7507
rect -3652 7405 -3618 7439
rect -3652 7337 -3618 7371
rect -3652 7269 -3618 7303
rect -3652 7201 -3618 7235
rect -3652 7133 -3618 7167
rect -3652 7065 -3618 7099
rect -3652 6997 -3618 7031
rect -3652 6929 -3618 6963
rect -3652 6861 -3618 6895
rect -3652 6793 -3618 6827
rect -3652 6725 -3618 6759
rect -3652 6657 -3618 6691
rect -3652 6589 -3618 6623
rect -3652 6521 -3618 6555
rect -3652 6453 -3618 6487
rect -3652 6385 -3618 6419
rect -3652 6317 -3618 6351
rect -3652 6249 -3618 6283
rect -3652 6181 -3618 6215
rect -3652 6113 -3618 6147
rect -3652 6045 -3618 6079
rect -3652 5977 -3618 6011
rect -3652 5909 -3618 5943
rect -3652 5841 -3618 5875
rect -3652 5773 -3618 5807
rect -3652 5705 -3618 5739
rect -3652 5637 -3618 5671
rect -3652 5569 -3618 5603
rect 17434 7493 17468 7527
rect 17434 7425 17468 7459
rect 17434 7357 17468 7391
rect 17434 7289 17468 7323
rect 17434 7221 17468 7255
rect 17434 7153 17468 7187
rect 17434 7085 17468 7119
rect 17434 7017 17468 7051
rect 17434 6949 17468 6983
rect 17434 6881 17468 6915
rect 17434 6813 17468 6847
rect 17434 6745 17468 6779
rect 17434 6677 17468 6711
rect 17434 6609 17468 6643
rect 17434 6541 17468 6575
rect 17434 6473 17468 6507
rect 17434 6405 17468 6439
rect 17434 6337 17468 6371
rect 17434 6269 17468 6303
rect 17434 6201 17468 6235
rect 17434 6133 17468 6167
rect 17434 6065 17468 6099
rect 17434 5997 17468 6031
rect 17434 5929 17468 5963
rect 17434 5861 17468 5895
rect 17434 5793 17468 5827
rect 17434 5725 17468 5759
rect 17434 5657 17468 5691
rect 17434 5589 17468 5623
rect 17434 5521 17468 5555
rect 17434 5453 17468 5487
rect 17434 5385 17468 5419
rect 17434 5317 17468 5351
rect 17434 5249 17468 5283
rect 17434 5181 17468 5215
rect 17434 5113 17468 5147
rect 17434 5045 17468 5079
rect 17434 4977 17468 5011
rect 17434 4909 17468 4943
rect 17434 4841 17468 4875
rect 17434 4773 17468 4807
rect 17434 4705 17468 4739
rect 17434 4637 17468 4671
rect 17434 4569 17468 4603
rect 18492 7493 18526 7527
rect 18492 7425 18526 7459
rect 18492 7357 18526 7391
rect 18492 7289 18526 7323
rect 18492 7221 18526 7255
rect 18492 7153 18526 7187
rect 18492 7085 18526 7119
rect 18492 7017 18526 7051
rect 18492 6949 18526 6983
rect 18492 6881 18526 6915
rect 18492 6813 18526 6847
rect 18492 6745 18526 6779
rect 18492 6677 18526 6711
rect 18492 6609 18526 6643
rect 18492 6541 18526 6575
rect 18492 6473 18526 6507
rect 18492 6405 18526 6439
rect 18492 6337 18526 6371
rect 18492 6269 18526 6303
rect 18492 6201 18526 6235
rect 18492 6133 18526 6167
rect 18492 6065 18526 6099
rect 18492 5997 18526 6031
rect 18492 5929 18526 5963
rect 18492 5861 18526 5895
rect 18492 5793 18526 5827
rect 18492 5725 18526 5759
rect 18492 5657 18526 5691
rect 18492 5589 18526 5623
rect 18492 5521 18526 5555
rect 18492 5453 18526 5487
rect 18492 5385 18526 5419
rect 18492 5317 18526 5351
rect 18492 5249 18526 5283
rect 18492 5181 18526 5215
rect 18492 5113 18526 5147
rect 18492 5045 18526 5079
rect 18492 4977 18526 5011
rect 18492 4909 18526 4943
rect 18492 4841 18526 4875
rect 18492 4773 18526 4807
rect 18492 4705 18526 4739
rect 18492 4637 18526 4671
rect 18492 4569 18526 4603
rect 18884 7493 18918 7527
rect 18884 7425 18918 7459
rect 18884 7357 18918 7391
rect 18884 7289 18918 7323
rect 18884 7221 18918 7255
rect 18884 7153 18918 7187
rect 18884 7085 18918 7119
rect 18884 7017 18918 7051
rect 18884 6949 18918 6983
rect 18884 6881 18918 6915
rect 18884 6813 18918 6847
rect 18884 6745 18918 6779
rect 18884 6677 18918 6711
rect 18884 6609 18918 6643
rect 18884 6541 18918 6575
rect 18884 6473 18918 6507
rect 18884 6405 18918 6439
rect 18884 6337 18918 6371
rect 18884 6269 18918 6303
rect 18884 6201 18918 6235
rect 18884 6133 18918 6167
rect 18884 6065 18918 6099
rect 18884 5997 18918 6031
rect 18884 5929 18918 5963
rect 18884 5861 18918 5895
rect 18884 5793 18918 5827
rect 18884 5725 18918 5759
rect 18884 5657 18918 5691
rect 18884 5589 18918 5623
rect 18884 5521 18918 5555
rect 18884 5453 18918 5487
rect 18884 5385 18918 5419
rect 18884 5317 18918 5351
rect 18884 5249 18918 5283
rect 18884 5181 18918 5215
rect 18884 5113 18918 5147
rect 18884 5045 18918 5079
rect 18884 4977 18918 5011
rect 18884 4909 18918 4943
rect 18884 4841 18918 4875
rect 18884 4773 18918 4807
rect 18884 4705 18918 4739
rect 18884 4637 18918 4671
rect 18884 4569 18918 4603
rect 19942 7493 19976 7527
rect 19942 7425 19976 7459
rect 19942 7357 19976 7391
rect 19942 7289 19976 7323
rect 19942 7221 19976 7255
rect 19942 7153 19976 7187
rect 19942 7085 19976 7119
rect 19942 7017 19976 7051
rect 19942 6949 19976 6983
rect 19942 6881 19976 6915
rect 19942 6813 19976 6847
rect 19942 6745 19976 6779
rect 19942 6677 19976 6711
rect 19942 6609 19976 6643
rect 19942 6541 19976 6575
rect 19942 6473 19976 6507
rect 19942 6405 19976 6439
rect 19942 6337 19976 6371
rect 19942 6269 19976 6303
rect 19942 6201 19976 6235
rect 19942 6133 19976 6167
rect 19942 6065 19976 6099
rect 19942 5997 19976 6031
rect 19942 5929 19976 5963
rect 19942 5861 19976 5895
rect 19942 5793 19976 5827
rect 19942 5725 19976 5759
rect 19942 5657 19976 5691
rect 19942 5589 19976 5623
rect 19942 5521 19976 5555
rect 19942 5453 19976 5487
rect 19942 5385 19976 5419
rect 19942 5317 19976 5351
rect 19942 5249 19976 5283
rect 19942 5181 19976 5215
rect 19942 5113 19976 5147
rect 19942 5045 19976 5079
rect 19942 4977 19976 5011
rect 19942 4909 19976 4943
rect 19942 4841 19976 4875
rect 19942 4773 19976 4807
rect 19942 4705 19976 4739
rect 19942 4637 19976 4671
rect 19942 4569 19976 4603
rect 38133 15520 38167 15554
rect 38133 15452 38167 15486
rect 38133 15384 38167 15418
rect 38133 15316 38167 15350
rect 38133 15248 38167 15282
rect 38133 15180 38167 15214
rect 38133 15112 38167 15146
rect 38133 15044 38167 15078
rect 38133 14976 38167 15010
rect 38133 14908 38167 14942
rect 38133 14840 38167 14874
rect 38133 14772 38167 14806
rect 38133 14704 38167 14738
rect 38133 14636 38167 14670
rect 38133 14568 38167 14602
rect 38133 14500 38167 14534
rect 38133 14432 38167 14466
rect 38133 14364 38167 14398
rect 38133 14296 38167 14330
rect 38133 14228 38167 14262
rect 38133 14160 38167 14194
rect 38133 14092 38167 14126
rect 38133 14024 38167 14058
rect 38133 13956 38167 13990
rect 38133 13888 38167 13922
rect 38133 13820 38167 13854
rect 38133 13752 38167 13786
rect 38133 13684 38167 13718
rect 38133 13616 38167 13650
rect 38391 15520 38425 15554
rect 38391 15452 38425 15486
rect 38391 15384 38425 15418
rect 38391 15316 38425 15350
rect 38391 15248 38425 15282
rect 38391 15180 38425 15214
rect 38391 15112 38425 15146
rect 38391 15044 38425 15078
rect 38391 14976 38425 15010
rect 38391 14908 38425 14942
rect 38391 14840 38425 14874
rect 38391 14772 38425 14806
rect 38391 14704 38425 14738
rect 38391 14636 38425 14670
rect 38391 14568 38425 14602
rect 38391 14500 38425 14534
rect 38391 14432 38425 14466
rect 38391 14364 38425 14398
rect 38391 14296 38425 14330
rect 38391 14228 38425 14262
rect 38391 14160 38425 14194
rect 38391 14092 38425 14126
rect 38391 14024 38425 14058
rect 38391 13956 38425 13990
rect 38391 13888 38425 13922
rect 38391 13820 38425 13854
rect 38391 13752 38425 13786
rect 38391 13684 38425 13718
rect 38391 13616 38425 13650
rect 38649 15520 38683 15554
rect 38649 15452 38683 15486
rect 38649 15384 38683 15418
rect 38649 15316 38683 15350
rect 38649 15248 38683 15282
rect 38649 15180 38683 15214
rect 38649 15112 38683 15146
rect 38649 15044 38683 15078
rect 38649 14976 38683 15010
rect 38649 14908 38683 14942
rect 38649 14840 38683 14874
rect 38649 14772 38683 14806
rect 38649 14704 38683 14738
rect 38649 14636 38683 14670
rect 38649 14568 38683 14602
rect 38649 14500 38683 14534
rect 38649 14432 38683 14466
rect 38649 14364 38683 14398
rect 38649 14296 38683 14330
rect 38649 14228 38683 14262
rect 38649 14160 38683 14194
rect 38649 14092 38683 14126
rect 38649 14024 38683 14058
rect 38649 13956 38683 13990
rect 38649 13888 38683 13922
rect 38649 13820 38683 13854
rect 38649 13752 38683 13786
rect 38649 13684 38683 13718
rect 38649 13616 38683 13650
rect 38907 15520 38941 15554
rect 38907 15452 38941 15486
rect 38907 15384 38941 15418
rect 38907 15316 38941 15350
rect 38907 15248 38941 15282
rect 38907 15180 38941 15214
rect 38907 15112 38941 15146
rect 38907 15044 38941 15078
rect 38907 14976 38941 15010
rect 38907 14908 38941 14942
rect 38907 14840 38941 14874
rect 38907 14772 38941 14806
rect 38907 14704 38941 14738
rect 38907 14636 38941 14670
rect 38907 14568 38941 14602
rect 38907 14500 38941 14534
rect 38907 14432 38941 14466
rect 38907 14364 38941 14398
rect 38907 14296 38941 14330
rect 38907 14228 38941 14262
rect 38907 14160 38941 14194
rect 38907 14092 38941 14126
rect 38907 14024 38941 14058
rect 38907 13956 38941 13990
rect 38907 13888 38941 13922
rect 38907 13820 38941 13854
rect 38907 13752 38941 13786
rect 38907 13684 38941 13718
rect 38907 13616 38941 13650
rect 39165 15520 39199 15554
rect 39165 15452 39199 15486
rect 39165 15384 39199 15418
rect 39165 15316 39199 15350
rect 39165 15248 39199 15282
rect 39165 15180 39199 15214
rect 39165 15112 39199 15146
rect 39165 15044 39199 15078
rect 39165 14976 39199 15010
rect 39165 14908 39199 14942
rect 39165 14840 39199 14874
rect 39165 14772 39199 14806
rect 39165 14704 39199 14738
rect 39165 14636 39199 14670
rect 39165 14568 39199 14602
rect 39165 14500 39199 14534
rect 39165 14432 39199 14466
rect 39165 14364 39199 14398
rect 39165 14296 39199 14330
rect 39165 14228 39199 14262
rect 39165 14160 39199 14194
rect 39165 14092 39199 14126
rect 39165 14024 39199 14058
rect 39165 13956 39199 13990
rect 39165 13888 39199 13922
rect 39165 13820 39199 13854
rect 39165 13752 39199 13786
rect 39165 13684 39199 13718
rect 39165 13616 39199 13650
rect 39423 15520 39457 15554
rect 39423 15452 39457 15486
rect 39423 15384 39457 15418
rect 39423 15316 39457 15350
rect 39423 15248 39457 15282
rect 39423 15180 39457 15214
rect 39423 15112 39457 15146
rect 39423 15044 39457 15078
rect 39423 14976 39457 15010
rect 39423 14908 39457 14942
rect 39423 14840 39457 14874
rect 39423 14772 39457 14806
rect 39423 14704 39457 14738
rect 39423 14636 39457 14670
rect 39423 14568 39457 14602
rect 39423 14500 39457 14534
rect 39423 14432 39457 14466
rect 39423 14364 39457 14398
rect 39423 14296 39457 14330
rect 39423 14228 39457 14262
rect 39423 14160 39457 14194
rect 39423 14092 39457 14126
rect 39423 14024 39457 14058
rect 39423 13956 39457 13990
rect 39423 13888 39457 13922
rect 39423 13820 39457 13854
rect 39423 13752 39457 13786
rect 39423 13684 39457 13718
rect 39423 13616 39457 13650
rect 39681 15520 39715 15554
rect 39681 15452 39715 15486
rect 39681 15384 39715 15418
rect 39681 15316 39715 15350
rect 39681 15248 39715 15282
rect 39681 15180 39715 15214
rect 39681 15112 39715 15146
rect 39681 15044 39715 15078
rect 39681 14976 39715 15010
rect 39681 14908 39715 14942
rect 39681 14840 39715 14874
rect 39681 14772 39715 14806
rect 39681 14704 39715 14738
rect 39681 14636 39715 14670
rect 39681 14568 39715 14602
rect 39681 14500 39715 14534
rect 39681 14432 39715 14466
rect 39681 14364 39715 14398
rect 39681 14296 39715 14330
rect 39681 14228 39715 14262
rect 39681 14160 39715 14194
rect 39681 14092 39715 14126
rect 39681 14024 39715 14058
rect 39681 13956 39715 13990
rect 39681 13888 39715 13922
rect 39681 13820 39715 13854
rect 39681 13752 39715 13786
rect 39681 13684 39715 13718
rect 39681 13616 39715 13650
rect 39939 15520 39973 15554
rect 39939 15452 39973 15486
rect 39939 15384 39973 15418
rect 39939 15316 39973 15350
rect 39939 15248 39973 15282
rect 39939 15180 39973 15214
rect 39939 15112 39973 15146
rect 39939 15044 39973 15078
rect 39939 14976 39973 15010
rect 39939 14908 39973 14942
rect 39939 14840 39973 14874
rect 39939 14772 39973 14806
rect 39939 14704 39973 14738
rect 39939 14636 39973 14670
rect 39939 14568 39973 14602
rect 39939 14500 39973 14534
rect 39939 14432 39973 14466
rect 39939 14364 39973 14398
rect 39939 14296 39973 14330
rect 39939 14228 39973 14262
rect 39939 14160 39973 14194
rect 39939 14092 39973 14126
rect 39939 14024 39973 14058
rect 39939 13956 39973 13990
rect 39939 13888 39973 13922
rect 39939 13820 39973 13854
rect 39939 13752 39973 13786
rect 39939 13684 39973 13718
rect 39939 13616 39973 13650
rect 40197 15520 40231 15554
rect 40197 15452 40231 15486
rect 40197 15384 40231 15418
rect 40197 15316 40231 15350
rect 40197 15248 40231 15282
rect 40197 15180 40231 15214
rect 40197 15112 40231 15146
rect 40197 15044 40231 15078
rect 40197 14976 40231 15010
rect 40197 14908 40231 14942
rect 40197 14840 40231 14874
rect 40197 14772 40231 14806
rect 40197 14704 40231 14738
rect 40197 14636 40231 14670
rect 40197 14568 40231 14602
rect 40197 14500 40231 14534
rect 40197 14432 40231 14466
rect 40197 14364 40231 14398
rect 40197 14296 40231 14330
rect 40197 14228 40231 14262
rect 40197 14160 40231 14194
rect 40197 14092 40231 14126
rect 40197 14024 40231 14058
rect 40197 13956 40231 13990
rect 40197 13888 40231 13922
rect 40197 13820 40231 13854
rect 40197 13752 40231 13786
rect 40197 13684 40231 13718
rect 40197 13616 40231 13650
rect 40455 15520 40489 15554
rect 40455 15452 40489 15486
rect 40455 15384 40489 15418
rect 40455 15316 40489 15350
rect 40455 15248 40489 15282
rect 40455 15180 40489 15214
rect 40455 15112 40489 15146
rect 40455 15044 40489 15078
rect 40455 14976 40489 15010
rect 40455 14908 40489 14942
rect 40455 14840 40489 14874
rect 40455 14772 40489 14806
rect 40455 14704 40489 14738
rect 40455 14636 40489 14670
rect 40455 14568 40489 14602
rect 40455 14500 40489 14534
rect 40455 14432 40489 14466
rect 40455 14364 40489 14398
rect 40455 14296 40489 14330
rect 40455 14228 40489 14262
rect 40455 14160 40489 14194
rect 40455 14092 40489 14126
rect 40455 14024 40489 14058
rect 40455 13956 40489 13990
rect 40455 13888 40489 13922
rect 40455 13820 40489 13854
rect 40455 13752 40489 13786
rect 40455 13684 40489 13718
rect 40455 13616 40489 13650
rect 40713 15520 40747 15554
rect 40713 15452 40747 15486
rect 40713 15384 40747 15418
rect 40713 15316 40747 15350
rect 40713 15248 40747 15282
rect 40713 15180 40747 15214
rect 40713 15112 40747 15146
rect 40713 15044 40747 15078
rect 40713 14976 40747 15010
rect 40713 14908 40747 14942
rect 40713 14840 40747 14874
rect 40713 14772 40747 14806
rect 40713 14704 40747 14738
rect 40713 14636 40747 14670
rect 40713 14568 40747 14602
rect 40713 14500 40747 14534
rect 40713 14432 40747 14466
rect 40713 14364 40747 14398
rect 40713 14296 40747 14330
rect 40713 14228 40747 14262
rect 40713 14160 40747 14194
rect 40713 14092 40747 14126
rect 40713 14024 40747 14058
rect 40713 13956 40747 13990
rect 40713 13888 40747 13922
rect 40713 13820 40747 13854
rect 40713 13752 40747 13786
rect 40713 13684 40747 13718
rect 40713 13616 40747 13650
rect 23171 11782 23205 11816
rect 23239 11782 23273 11816
rect 23307 11782 23341 11816
rect 23375 11782 23409 11816
rect 23443 11782 23477 11816
rect 23511 11782 23545 11816
rect 23579 11782 23613 11816
rect 23647 11782 23681 11816
rect 23715 11782 23749 11816
rect 23783 11782 23817 11816
rect 23851 11782 23885 11816
rect 23919 11782 23953 11816
rect 23987 11782 24021 11816
rect 24055 11782 24089 11816
rect 23171 10724 23205 10758
rect 23239 10724 23273 10758
rect 23307 10724 23341 10758
rect 23375 10724 23409 10758
rect 23443 10724 23477 10758
rect 23511 10724 23545 10758
rect 23579 10724 23613 10758
rect 23647 10724 23681 10758
rect 23715 10724 23749 10758
rect 23783 10724 23817 10758
rect 23851 10724 23885 10758
rect 23919 10724 23953 10758
rect 23987 10724 24021 10758
rect 24055 10724 24089 10758
rect 23651 7846 23685 7880
rect 23719 7846 23753 7880
rect 23787 7846 23821 7880
rect 23855 7846 23889 7880
rect 23923 7846 23957 7880
rect 23991 7846 24025 7880
rect 24059 7846 24093 7880
rect 24127 7846 24161 7880
rect 24195 7846 24229 7880
rect 24263 7846 24297 7880
rect 24331 7846 24365 7880
rect 24399 7846 24433 7880
rect 24467 7846 24501 7880
rect 24535 7846 24569 7880
rect 23651 6788 23685 6822
rect 23719 6788 23753 6822
rect 23787 6788 23821 6822
rect 23855 6788 23889 6822
rect 23923 6788 23957 6822
rect 23991 6788 24025 6822
rect 24059 6788 24093 6822
rect 24127 6788 24161 6822
rect 24195 6788 24229 6822
rect 24263 6788 24297 6822
rect 24331 6788 24365 6822
rect 24399 6788 24433 6822
rect 24467 6788 24501 6822
rect 24535 6788 24569 6822
rect 23651 5730 23685 5764
rect 23719 5730 23753 5764
rect 23787 5730 23821 5764
rect 23855 5730 23889 5764
rect 23923 5730 23957 5764
rect 23991 5730 24025 5764
rect 24059 5730 24093 5764
rect 24127 5730 24161 5764
rect 24195 5730 24229 5764
rect 24263 5730 24297 5764
rect 24331 5730 24365 5764
rect 24399 5730 24433 5764
rect 24467 5730 24501 5764
rect 24535 5730 24569 5764
rect 23651 4672 23685 4706
rect 23719 4672 23753 4706
rect 23787 4672 23821 4706
rect 23855 4672 23889 4706
rect 23923 4672 23957 4706
rect 23991 4672 24025 4706
rect 24059 4672 24093 4706
rect 24127 4672 24161 4706
rect 24195 4672 24229 4706
rect 24263 4672 24297 4706
rect 24331 4672 24365 4706
rect 24399 4672 24433 4706
rect 24467 4672 24501 4706
rect 24535 4672 24569 4706
rect 23651 3614 23685 3648
rect 23719 3614 23753 3648
rect 23787 3614 23821 3648
rect 23855 3614 23889 3648
rect 23923 3614 23957 3648
rect 23991 3614 24025 3648
rect 24059 3614 24093 3648
rect 24127 3614 24161 3648
rect 24195 3614 24229 3648
rect 24263 3614 24297 3648
rect 24331 3614 24365 3648
rect 24399 3614 24433 3648
rect 24467 3614 24501 3648
rect 24535 3614 24569 3648
rect 25151 7846 25185 7880
rect 25219 7846 25253 7880
rect 25287 7846 25321 7880
rect 25355 7846 25389 7880
rect 25423 7846 25457 7880
rect 25491 7846 25525 7880
rect 25559 7846 25593 7880
rect 25627 7846 25661 7880
rect 25695 7846 25729 7880
rect 25763 7846 25797 7880
rect 25831 7846 25865 7880
rect 25899 7846 25933 7880
rect 25967 7846 26001 7880
rect 26035 7846 26069 7880
rect 25151 6788 25185 6822
rect 25219 6788 25253 6822
rect 25287 6788 25321 6822
rect 25355 6788 25389 6822
rect 25423 6788 25457 6822
rect 25491 6788 25525 6822
rect 25559 6788 25593 6822
rect 25627 6788 25661 6822
rect 25695 6788 25729 6822
rect 25763 6788 25797 6822
rect 25831 6788 25865 6822
rect 25899 6788 25933 6822
rect 25967 6788 26001 6822
rect 26035 6788 26069 6822
rect 25151 5730 25185 5764
rect 25219 5730 25253 5764
rect 25287 5730 25321 5764
rect 25355 5730 25389 5764
rect 25423 5730 25457 5764
rect 25491 5730 25525 5764
rect 25559 5730 25593 5764
rect 25627 5730 25661 5764
rect 25695 5730 25729 5764
rect 25763 5730 25797 5764
rect 25831 5730 25865 5764
rect 25899 5730 25933 5764
rect 25967 5730 26001 5764
rect 26035 5730 26069 5764
rect 25151 4672 25185 4706
rect 25219 4672 25253 4706
rect 25287 4672 25321 4706
rect 25355 4672 25389 4706
rect 25423 4672 25457 4706
rect 25491 4672 25525 4706
rect 25559 4672 25593 4706
rect 25627 4672 25661 4706
rect 25695 4672 25729 4706
rect 25763 4672 25797 4706
rect 25831 4672 25865 4706
rect 25899 4672 25933 4706
rect 25967 4672 26001 4706
rect 26035 4672 26069 4706
rect 25151 3614 25185 3648
rect 25219 3614 25253 3648
rect 25287 3614 25321 3648
rect 25355 3614 25389 3648
rect 25423 3614 25457 3648
rect 25491 3614 25525 3648
rect 25559 3614 25593 3648
rect 25627 3614 25661 3648
rect 25695 3614 25729 3648
rect 25763 3614 25797 3648
rect 25831 3614 25865 3648
rect 25899 3614 25933 3648
rect 25967 3614 26001 3648
rect 26035 3614 26069 3648
rect 36777 11839 36811 11873
rect 36777 11771 36811 11805
rect 36777 11703 36811 11737
rect 36777 11635 36811 11669
rect 36777 11567 36811 11601
rect 36777 11499 36811 11533
rect 36777 11431 36811 11465
rect 36777 11363 36811 11397
rect 36777 11295 36811 11329
rect 36777 11227 36811 11261
rect 36777 11159 36811 11193
rect 36777 11091 36811 11125
rect 36777 11023 36811 11057
rect 36777 10955 36811 10989
rect 37035 11839 37069 11873
rect 37035 11771 37069 11805
rect 37035 11703 37069 11737
rect 37035 11635 37069 11669
rect 37035 11567 37069 11601
rect 37035 11499 37069 11533
rect 37035 11431 37069 11465
rect 37035 11363 37069 11397
rect 37035 11295 37069 11329
rect 37035 11227 37069 11261
rect 37035 11159 37069 11193
rect 37035 11091 37069 11125
rect 37035 11023 37069 11057
rect 37035 10955 37069 10989
rect 37293 11839 37327 11873
rect 37293 11771 37327 11805
rect 37293 11703 37327 11737
rect 37293 11635 37327 11669
rect 37293 11567 37327 11601
rect 37293 11499 37327 11533
rect 37293 11431 37327 11465
rect 37293 11363 37327 11397
rect 37293 11295 37327 11329
rect 37293 11227 37327 11261
rect 37293 11159 37327 11193
rect 37293 11091 37327 11125
rect 37293 11023 37327 11057
rect 37293 10955 37327 10989
rect 37551 11839 37585 11873
rect 37551 11771 37585 11805
rect 37551 11703 37585 11737
rect 37551 11635 37585 11669
rect 37551 11567 37585 11601
rect 37551 11499 37585 11533
rect 37551 11431 37585 11465
rect 37551 11363 37585 11397
rect 37551 11295 37585 11329
rect 37551 11227 37585 11261
rect 37551 11159 37585 11193
rect 37551 11091 37585 11125
rect 37551 11023 37585 11057
rect 37551 10955 37585 10989
rect 37809 11839 37843 11873
rect 37809 11771 37843 11805
rect 37809 11703 37843 11737
rect 37809 11635 37843 11669
rect 37809 11567 37843 11601
rect 37809 11499 37843 11533
rect 37809 11431 37843 11465
rect 37809 11363 37843 11397
rect 37809 11295 37843 11329
rect 37809 11227 37843 11261
rect 37809 11159 37843 11193
rect 37809 11091 37843 11125
rect 37809 11023 37843 11057
rect 37809 10955 37843 10989
rect 38067 11839 38101 11873
rect 38067 11771 38101 11805
rect 38067 11703 38101 11737
rect 38067 11635 38101 11669
rect 38067 11567 38101 11601
rect 38067 11499 38101 11533
rect 38067 11431 38101 11465
rect 38067 11363 38101 11397
rect 38067 11295 38101 11329
rect 38067 11227 38101 11261
rect 38067 11159 38101 11193
rect 38067 11091 38101 11125
rect 38067 11023 38101 11057
rect 38067 10955 38101 10989
rect 38325 11839 38359 11873
rect 38325 11771 38359 11805
rect 38325 11703 38359 11737
rect 38325 11635 38359 11669
rect 38325 11567 38359 11601
rect 38325 11499 38359 11533
rect 38325 11431 38359 11465
rect 38325 11363 38359 11397
rect 38325 11295 38359 11329
rect 38325 11227 38359 11261
rect 38325 11159 38359 11193
rect 38325 11091 38359 11125
rect 38325 11023 38359 11057
rect 38325 10955 38359 10989
rect 38583 11839 38617 11873
rect 38583 11771 38617 11805
rect 38583 11703 38617 11737
rect 38583 11635 38617 11669
rect 38583 11567 38617 11601
rect 38583 11499 38617 11533
rect 38583 11431 38617 11465
rect 38583 11363 38617 11397
rect 38583 11295 38617 11329
rect 38583 11227 38617 11261
rect 38583 11159 38617 11193
rect 38583 11091 38617 11125
rect 38583 11023 38617 11057
rect 38583 10955 38617 10989
rect 38841 11839 38875 11873
rect 38841 11771 38875 11805
rect 38841 11703 38875 11737
rect 38841 11635 38875 11669
rect 38841 11567 38875 11601
rect 38841 11499 38875 11533
rect 38841 11431 38875 11465
rect 38841 11363 38875 11397
rect 38841 11295 38875 11329
rect 38841 11227 38875 11261
rect 38841 11159 38875 11193
rect 38841 11091 38875 11125
rect 38841 11023 38875 11057
rect 38841 10955 38875 10989
rect 39099 11839 39133 11873
rect 39099 11771 39133 11805
rect 39099 11703 39133 11737
rect 39099 11635 39133 11669
rect 39099 11567 39133 11601
rect 39099 11499 39133 11533
rect 39099 11431 39133 11465
rect 39099 11363 39133 11397
rect 39099 11295 39133 11329
rect 39099 11227 39133 11261
rect 39099 11159 39133 11193
rect 39099 11091 39133 11125
rect 39099 11023 39133 11057
rect 39099 10955 39133 10989
rect 39357 11839 39391 11873
rect 39357 11771 39391 11805
rect 39357 11703 39391 11737
rect 39357 11635 39391 11669
rect 39357 11567 39391 11601
rect 39357 11499 39391 11533
rect 39357 11431 39391 11465
rect 39357 11363 39391 11397
rect 39357 11295 39391 11329
rect 39357 11227 39391 11261
rect 39357 11159 39391 11193
rect 39357 11091 39391 11125
rect 39357 11023 39391 11057
rect 39357 10955 39391 10989
rect 39615 11839 39649 11873
rect 39615 11771 39649 11805
rect 39615 11703 39649 11737
rect 39615 11635 39649 11669
rect 39615 11567 39649 11601
rect 39615 11499 39649 11533
rect 39615 11431 39649 11465
rect 39615 11363 39649 11397
rect 39615 11295 39649 11329
rect 39615 11227 39649 11261
rect 39615 11159 39649 11193
rect 39615 11091 39649 11125
rect 39615 11023 39649 11057
rect 39615 10955 39649 10989
rect 39873 11839 39907 11873
rect 39873 11771 39907 11805
rect 39873 11703 39907 11737
rect 39873 11635 39907 11669
rect 39873 11567 39907 11601
rect 39873 11499 39907 11533
rect 39873 11431 39907 11465
rect 39873 11363 39907 11397
rect 39873 11295 39907 11329
rect 39873 11227 39907 11261
rect 39873 11159 39907 11193
rect 39873 11091 39907 11125
rect 39873 11023 39907 11057
rect 39873 10955 39907 10989
rect 40131 11839 40165 11873
rect 40131 11771 40165 11805
rect 40131 11703 40165 11737
rect 40131 11635 40165 11669
rect 40131 11567 40165 11601
rect 40131 11499 40165 11533
rect 40131 11431 40165 11465
rect 40131 11363 40165 11397
rect 40131 11295 40165 11329
rect 40131 11227 40165 11261
rect 40131 11159 40165 11193
rect 40131 11091 40165 11125
rect 40131 11023 40165 11057
rect 40131 10955 40165 10989
rect 40389 11839 40423 11873
rect 40389 11771 40423 11805
rect 40389 11703 40423 11737
rect 40389 11635 40423 11669
rect 40389 11567 40423 11601
rect 40389 11499 40423 11533
rect 40389 11431 40423 11465
rect 40389 11363 40423 11397
rect 40389 11295 40423 11329
rect 40389 11227 40423 11261
rect 40389 11159 40423 11193
rect 40389 11091 40423 11125
rect 40389 11023 40423 11057
rect 40389 10955 40423 10989
rect 40647 11839 40681 11873
rect 40647 11771 40681 11805
rect 40647 11703 40681 11737
rect 40647 11635 40681 11669
rect 40647 11567 40681 11601
rect 40647 11499 40681 11533
rect 40647 11431 40681 11465
rect 40647 11363 40681 11397
rect 40647 11295 40681 11329
rect 40647 11227 40681 11261
rect 40647 11159 40681 11193
rect 40647 11091 40681 11125
rect 40647 11023 40681 11057
rect 40647 10955 40681 10989
rect 40905 11839 40939 11873
rect 40905 11771 40939 11805
rect 40905 11703 40939 11737
rect 40905 11635 40939 11669
rect 40905 11567 40939 11601
rect 40905 11499 40939 11533
rect 40905 11431 40939 11465
rect 40905 11363 40939 11397
rect 40905 11295 40939 11329
rect 40905 11227 40939 11261
rect 40905 11159 40939 11193
rect 40905 11091 40939 11125
rect 40905 11023 40939 11057
rect 40905 10955 40939 10989
rect 41163 11839 41197 11873
rect 41163 11771 41197 11805
rect 41163 11703 41197 11737
rect 41163 11635 41197 11669
rect 41163 11567 41197 11601
rect 41163 11499 41197 11533
rect 41163 11431 41197 11465
rect 41163 11363 41197 11397
rect 41163 11295 41197 11329
rect 41163 11227 41197 11261
rect 41163 11159 41197 11193
rect 41163 11091 41197 11125
rect 41163 11023 41197 11057
rect 41163 10955 41197 10989
rect 41421 11839 41455 11873
rect 41421 11771 41455 11805
rect 41421 11703 41455 11737
rect 41421 11635 41455 11669
rect 41421 11567 41455 11601
rect 41421 11499 41455 11533
rect 41421 11431 41455 11465
rect 41421 11363 41455 11397
rect 41421 11295 41455 11329
rect 41421 11227 41455 11261
rect 41421 11159 41455 11193
rect 41421 11091 41455 11125
rect 41421 11023 41455 11057
rect 41421 10955 41455 10989
rect 41679 11839 41713 11873
rect 41679 11771 41713 11805
rect 41679 11703 41713 11737
rect 41679 11635 41713 11669
rect 41679 11567 41713 11601
rect 41679 11499 41713 11533
rect 41679 11431 41713 11465
rect 41679 11363 41713 11397
rect 41679 11295 41713 11329
rect 41679 11227 41713 11261
rect 41679 11159 41713 11193
rect 41679 11091 41713 11125
rect 41679 11023 41713 11057
rect 41679 10955 41713 10989
rect 41937 11839 41971 11873
rect 41937 11771 41971 11805
rect 41937 11703 41971 11737
rect 41937 11635 41971 11669
rect 41937 11567 41971 11601
rect 41937 11499 41971 11533
rect 41937 11431 41971 11465
rect 41937 11363 41971 11397
rect 41937 11295 41971 11329
rect 41937 11227 41971 11261
rect 41937 11159 41971 11193
rect 41937 11091 41971 11125
rect 41937 11023 41971 11057
rect 41937 10955 41971 10989
rect 37812 10474 37846 10508
rect 37812 10406 37846 10440
rect 37812 10338 37846 10372
rect 37812 10270 37846 10304
rect 37812 10202 37846 10236
rect 37812 10134 37846 10168
rect 37812 10066 37846 10100
rect 37812 9998 37846 10032
rect 37812 9930 37846 9964
rect 37812 9862 37846 9896
rect 37812 9794 37846 9828
rect 37812 9726 37846 9760
rect 37812 9658 37846 9692
rect 37812 9590 37846 9624
rect 38070 10474 38104 10508
rect 38070 10406 38104 10440
rect 38070 10338 38104 10372
rect 38070 10270 38104 10304
rect 38070 10202 38104 10236
rect 38070 10134 38104 10168
rect 38070 10066 38104 10100
rect 38070 9998 38104 10032
rect 38070 9930 38104 9964
rect 38070 9862 38104 9896
rect 38070 9794 38104 9828
rect 38070 9726 38104 9760
rect 38070 9658 38104 9692
rect 38070 9590 38104 9624
rect 38278 10474 38312 10508
rect 38278 10406 38312 10440
rect 38278 10338 38312 10372
rect 38278 10270 38312 10304
rect 38278 10202 38312 10236
rect 38278 10134 38312 10168
rect 38278 10066 38312 10100
rect 38278 9998 38312 10032
rect 38278 9930 38312 9964
rect 38278 9862 38312 9896
rect 38278 9794 38312 9828
rect 38278 9726 38312 9760
rect 38278 9658 38312 9692
rect 38278 9590 38312 9624
rect 38536 10474 38570 10508
rect 38536 10406 38570 10440
rect 38536 10338 38570 10372
rect 38536 10270 38570 10304
rect 38536 10202 38570 10236
rect 38536 10134 38570 10168
rect 38536 10066 38570 10100
rect 38536 9998 38570 10032
rect 38536 9930 38570 9964
rect 38536 9862 38570 9896
rect 38536 9794 38570 9828
rect 38536 9726 38570 9760
rect 38536 9658 38570 9692
rect 38536 9590 38570 9624
rect 38794 10474 38828 10508
rect 38794 10406 38828 10440
rect 38794 10338 38828 10372
rect 38794 10270 38828 10304
rect 38794 10202 38828 10236
rect 38794 10134 38828 10168
rect 38794 10066 38828 10100
rect 38794 9998 38828 10032
rect 38794 9930 38828 9964
rect 38794 9862 38828 9896
rect 38794 9794 38828 9828
rect 38794 9726 38828 9760
rect 38794 9658 38828 9692
rect 38794 9590 38828 9624
rect 39052 10474 39086 10508
rect 39052 10406 39086 10440
rect 39052 10338 39086 10372
rect 39052 10270 39086 10304
rect 39052 10202 39086 10236
rect 39052 10134 39086 10168
rect 39052 10066 39086 10100
rect 39052 9998 39086 10032
rect 39052 9930 39086 9964
rect 39052 9862 39086 9896
rect 39052 9794 39086 9828
rect 39052 9726 39086 9760
rect 39052 9658 39086 9692
rect 39052 9590 39086 9624
rect 39310 10474 39344 10508
rect 39310 10406 39344 10440
rect 39310 10338 39344 10372
rect 39310 10270 39344 10304
rect 39310 10202 39344 10236
rect 39310 10134 39344 10168
rect 39310 10066 39344 10100
rect 39310 9998 39344 10032
rect 39310 9930 39344 9964
rect 39310 9862 39344 9896
rect 39310 9794 39344 9828
rect 39310 9726 39344 9760
rect 39310 9658 39344 9692
rect 39310 9590 39344 9624
rect 39568 10474 39602 10508
rect 39568 10406 39602 10440
rect 39568 10338 39602 10372
rect 39568 10270 39602 10304
rect 39568 10202 39602 10236
rect 39568 10134 39602 10168
rect 39568 10066 39602 10100
rect 39568 9998 39602 10032
rect 39568 9930 39602 9964
rect 39568 9862 39602 9896
rect 39568 9794 39602 9828
rect 39568 9726 39602 9760
rect 39568 9658 39602 9692
rect 39568 9590 39602 9624
rect 39826 10474 39860 10508
rect 39826 10406 39860 10440
rect 39826 10338 39860 10372
rect 39826 10270 39860 10304
rect 39826 10202 39860 10236
rect 39826 10134 39860 10168
rect 39826 10066 39860 10100
rect 39826 9998 39860 10032
rect 39826 9930 39860 9964
rect 39826 9862 39860 9896
rect 39826 9794 39860 9828
rect 39826 9726 39860 9760
rect 39826 9658 39860 9692
rect 39826 9590 39860 9624
rect 40084 10474 40118 10508
rect 40084 10406 40118 10440
rect 40084 10338 40118 10372
rect 40084 10270 40118 10304
rect 40084 10202 40118 10236
rect 40084 10134 40118 10168
rect 40084 10066 40118 10100
rect 40084 9998 40118 10032
rect 40084 9930 40118 9964
rect 40084 9862 40118 9896
rect 40084 9794 40118 9828
rect 40084 9726 40118 9760
rect 40084 9658 40118 9692
rect 40084 9590 40118 9624
rect 40342 10474 40376 10508
rect 40342 10406 40376 10440
rect 40342 10338 40376 10372
rect 40342 10270 40376 10304
rect 40342 10202 40376 10236
rect 40342 10134 40376 10168
rect 40342 10066 40376 10100
rect 40342 9998 40376 10032
rect 40342 9930 40376 9964
rect 40342 9862 40376 9896
rect 40342 9794 40376 9828
rect 40342 9726 40376 9760
rect 40342 9658 40376 9692
rect 40342 9590 40376 9624
rect 40600 10474 40634 10508
rect 40600 10406 40634 10440
rect 40600 10338 40634 10372
rect 40600 10270 40634 10304
rect 40600 10202 40634 10236
rect 40600 10134 40634 10168
rect 40600 10066 40634 10100
rect 40600 9998 40634 10032
rect 40600 9930 40634 9964
rect 40600 9862 40634 9896
rect 40600 9794 40634 9828
rect 40600 9726 40634 9760
rect 40600 9658 40634 9692
rect 40600 9590 40634 9624
rect 40858 10474 40892 10508
rect 40858 10406 40892 10440
rect 40858 10338 40892 10372
rect 40858 10270 40892 10304
rect 40858 10202 40892 10236
rect 40858 10134 40892 10168
rect 40858 10066 40892 10100
rect 40858 9998 40892 10032
rect 40858 9930 40892 9964
rect 40858 9862 40892 9896
rect 40858 9794 40892 9828
rect 40858 9726 40892 9760
rect 40858 9658 40892 9692
rect 40858 9590 40892 9624
rect 37812 8223 37846 8257
rect 37812 8155 37846 8189
rect 37812 8087 37846 8121
rect 37812 8019 37846 8053
rect 37812 7951 37846 7985
rect 37812 7883 37846 7917
rect 37812 7815 37846 7849
rect 37812 7747 37846 7781
rect 37812 7679 37846 7713
rect 37812 7611 37846 7645
rect 37812 7543 37846 7577
rect 37812 7475 37846 7509
rect 37812 7407 37846 7441
rect 37812 7339 37846 7373
rect 37812 7271 37846 7305
rect 37812 7203 37846 7237
rect 37812 7135 37846 7169
rect 37812 7067 37846 7101
rect 37812 6999 37846 7033
rect 37812 6931 37846 6965
rect 37812 6863 37846 6897
rect 37812 6795 37846 6829
rect 37812 6727 37846 6761
rect 37812 6659 37846 6693
rect 37812 6591 37846 6625
rect 37812 6523 37846 6557
rect 37812 6455 37846 6489
rect 37812 6387 37846 6421
rect 37812 6319 37846 6353
rect 38070 8223 38104 8257
rect 38070 8155 38104 8189
rect 38070 8087 38104 8121
rect 38070 8019 38104 8053
rect 38070 7951 38104 7985
rect 38070 7883 38104 7917
rect 38070 7815 38104 7849
rect 38070 7747 38104 7781
rect 38070 7679 38104 7713
rect 38070 7611 38104 7645
rect 38070 7543 38104 7577
rect 38070 7475 38104 7509
rect 38070 7407 38104 7441
rect 38070 7339 38104 7373
rect 38070 7271 38104 7305
rect 38070 7203 38104 7237
rect 38070 7135 38104 7169
rect 38070 7067 38104 7101
rect 38070 6999 38104 7033
rect 38070 6931 38104 6965
rect 38070 6863 38104 6897
rect 38070 6795 38104 6829
rect 38070 6727 38104 6761
rect 38070 6659 38104 6693
rect 38070 6591 38104 6625
rect 38070 6523 38104 6557
rect 38070 6455 38104 6489
rect 38070 6387 38104 6421
rect 38070 6319 38104 6353
rect 38328 8223 38362 8257
rect 38328 8155 38362 8189
rect 38328 8087 38362 8121
rect 38328 8019 38362 8053
rect 38328 7951 38362 7985
rect 38328 7883 38362 7917
rect 38328 7815 38362 7849
rect 38328 7747 38362 7781
rect 38328 7679 38362 7713
rect 38328 7611 38362 7645
rect 38328 7543 38362 7577
rect 38328 7475 38362 7509
rect 38328 7407 38362 7441
rect 38328 7339 38362 7373
rect 38328 7271 38362 7305
rect 38328 7203 38362 7237
rect 38328 7135 38362 7169
rect 38328 7067 38362 7101
rect 38328 6999 38362 7033
rect 38328 6931 38362 6965
rect 38328 6863 38362 6897
rect 38328 6795 38362 6829
rect 38328 6727 38362 6761
rect 38328 6659 38362 6693
rect 38328 6591 38362 6625
rect 38328 6523 38362 6557
rect 38328 6455 38362 6489
rect 38328 6387 38362 6421
rect 38328 6319 38362 6353
rect 38586 8223 38620 8257
rect 38586 8155 38620 8189
rect 38586 8087 38620 8121
rect 38586 8019 38620 8053
rect 38586 7951 38620 7985
rect 38586 7883 38620 7917
rect 38586 7815 38620 7849
rect 38586 7747 38620 7781
rect 38586 7679 38620 7713
rect 38586 7611 38620 7645
rect 38586 7543 38620 7577
rect 38586 7475 38620 7509
rect 38586 7407 38620 7441
rect 38586 7339 38620 7373
rect 38586 7271 38620 7305
rect 38586 7203 38620 7237
rect 38586 7135 38620 7169
rect 38586 7067 38620 7101
rect 38586 6999 38620 7033
rect 38586 6931 38620 6965
rect 38586 6863 38620 6897
rect 38586 6795 38620 6829
rect 38586 6727 38620 6761
rect 38586 6659 38620 6693
rect 38586 6591 38620 6625
rect 38586 6523 38620 6557
rect 38586 6455 38620 6489
rect 38586 6387 38620 6421
rect 38586 6319 38620 6353
rect 38844 8223 38878 8257
rect 38844 8155 38878 8189
rect 38844 8087 38878 8121
rect 38844 8019 38878 8053
rect 38844 7951 38878 7985
rect 38844 7883 38878 7917
rect 38844 7815 38878 7849
rect 38844 7747 38878 7781
rect 38844 7679 38878 7713
rect 38844 7611 38878 7645
rect 38844 7543 38878 7577
rect 38844 7475 38878 7509
rect 38844 7407 38878 7441
rect 38844 7339 38878 7373
rect 38844 7271 38878 7305
rect 38844 7203 38878 7237
rect 38844 7135 38878 7169
rect 38844 7067 38878 7101
rect 38844 6999 38878 7033
rect 38844 6931 38878 6965
rect 38844 6863 38878 6897
rect 38844 6795 38878 6829
rect 38844 6727 38878 6761
rect 38844 6659 38878 6693
rect 38844 6591 38878 6625
rect 38844 6523 38878 6557
rect 38844 6455 38878 6489
rect 38844 6387 38878 6421
rect 38844 6319 38878 6353
rect 39102 8223 39136 8257
rect 39102 8155 39136 8189
rect 39102 8087 39136 8121
rect 39102 8019 39136 8053
rect 39102 7951 39136 7985
rect 39102 7883 39136 7917
rect 39102 7815 39136 7849
rect 39102 7747 39136 7781
rect 39102 7679 39136 7713
rect 39102 7611 39136 7645
rect 39102 7543 39136 7577
rect 39102 7475 39136 7509
rect 39102 7407 39136 7441
rect 39102 7339 39136 7373
rect 39102 7271 39136 7305
rect 39102 7203 39136 7237
rect 39102 7135 39136 7169
rect 39102 7067 39136 7101
rect 39102 6999 39136 7033
rect 39102 6931 39136 6965
rect 39102 6863 39136 6897
rect 39102 6795 39136 6829
rect 39102 6727 39136 6761
rect 39102 6659 39136 6693
rect 39102 6591 39136 6625
rect 39102 6523 39136 6557
rect 39102 6455 39136 6489
rect 39102 6387 39136 6421
rect 39102 6319 39136 6353
rect 39360 8223 39394 8257
rect 39360 8155 39394 8189
rect 39360 8087 39394 8121
rect 39360 8019 39394 8053
rect 39360 7951 39394 7985
rect 39360 7883 39394 7917
rect 39360 7815 39394 7849
rect 39360 7747 39394 7781
rect 39360 7679 39394 7713
rect 39360 7611 39394 7645
rect 39360 7543 39394 7577
rect 39360 7475 39394 7509
rect 39360 7407 39394 7441
rect 39360 7339 39394 7373
rect 39360 7271 39394 7305
rect 39360 7203 39394 7237
rect 39360 7135 39394 7169
rect 39360 7067 39394 7101
rect 39360 6999 39394 7033
rect 39360 6931 39394 6965
rect 39360 6863 39394 6897
rect 39360 6795 39394 6829
rect 39360 6727 39394 6761
rect 39360 6659 39394 6693
rect 39360 6591 39394 6625
rect 39360 6523 39394 6557
rect 39360 6455 39394 6489
rect 39360 6387 39394 6421
rect 39360 6319 39394 6353
rect 39618 8223 39652 8257
rect 39618 8155 39652 8189
rect 39618 8087 39652 8121
rect 39618 8019 39652 8053
rect 39618 7951 39652 7985
rect 39618 7883 39652 7917
rect 39618 7815 39652 7849
rect 39618 7747 39652 7781
rect 39618 7679 39652 7713
rect 39618 7611 39652 7645
rect 39618 7543 39652 7577
rect 39618 7475 39652 7509
rect 39618 7407 39652 7441
rect 39618 7339 39652 7373
rect 39618 7271 39652 7305
rect 39618 7203 39652 7237
rect 39618 7135 39652 7169
rect 39618 7067 39652 7101
rect 39618 6999 39652 7033
rect 39618 6931 39652 6965
rect 39618 6863 39652 6897
rect 39618 6795 39652 6829
rect 39618 6727 39652 6761
rect 39618 6659 39652 6693
rect 39618 6591 39652 6625
rect 39618 6523 39652 6557
rect 39618 6455 39652 6489
rect 39618 6387 39652 6421
rect 39618 6319 39652 6353
rect 39876 8223 39910 8257
rect 39876 8155 39910 8189
rect 39876 8087 39910 8121
rect 39876 8019 39910 8053
rect 39876 7951 39910 7985
rect 39876 7883 39910 7917
rect 39876 7815 39910 7849
rect 39876 7747 39910 7781
rect 39876 7679 39910 7713
rect 39876 7611 39910 7645
rect 39876 7543 39910 7577
rect 39876 7475 39910 7509
rect 39876 7407 39910 7441
rect 39876 7339 39910 7373
rect 39876 7271 39910 7305
rect 39876 7203 39910 7237
rect 39876 7135 39910 7169
rect 39876 7067 39910 7101
rect 39876 6999 39910 7033
rect 39876 6931 39910 6965
rect 39876 6863 39910 6897
rect 39876 6795 39910 6829
rect 39876 6727 39910 6761
rect 39876 6659 39910 6693
rect 39876 6591 39910 6625
rect 39876 6523 39910 6557
rect 39876 6455 39910 6489
rect 39876 6387 39910 6421
rect 39876 6319 39910 6353
rect 40134 8223 40168 8257
rect 40134 8155 40168 8189
rect 40134 8087 40168 8121
rect 40134 8019 40168 8053
rect 40134 7951 40168 7985
rect 40134 7883 40168 7917
rect 40134 7815 40168 7849
rect 40134 7747 40168 7781
rect 40134 7679 40168 7713
rect 40134 7611 40168 7645
rect 40134 7543 40168 7577
rect 40134 7475 40168 7509
rect 40134 7407 40168 7441
rect 40134 7339 40168 7373
rect 40134 7271 40168 7305
rect 40134 7203 40168 7237
rect 40134 7135 40168 7169
rect 40134 7067 40168 7101
rect 40134 6999 40168 7033
rect 40134 6931 40168 6965
rect 40134 6863 40168 6897
rect 40134 6795 40168 6829
rect 40134 6727 40168 6761
rect 40134 6659 40168 6693
rect 40134 6591 40168 6625
rect 40134 6523 40168 6557
rect 40134 6455 40168 6489
rect 40134 6387 40168 6421
rect 40134 6319 40168 6353
rect 40392 8223 40426 8257
rect 40392 8155 40426 8189
rect 40392 8087 40426 8121
rect 40392 8019 40426 8053
rect 40392 7951 40426 7985
rect 40392 7883 40426 7917
rect 40392 7815 40426 7849
rect 40392 7747 40426 7781
rect 40392 7679 40426 7713
rect 40392 7611 40426 7645
rect 40392 7543 40426 7577
rect 40392 7475 40426 7509
rect 40392 7407 40426 7441
rect 40392 7339 40426 7373
rect 40392 7271 40426 7305
rect 40392 7203 40426 7237
rect 40392 7135 40426 7169
rect 40392 7067 40426 7101
rect 40392 6999 40426 7033
rect 40392 6931 40426 6965
rect 40392 6863 40426 6897
rect 40392 6795 40426 6829
rect 40392 6727 40426 6761
rect 40392 6659 40426 6693
rect 40392 6591 40426 6625
rect 40392 6523 40426 6557
rect 40392 6455 40426 6489
rect 40392 6387 40426 6421
rect 40392 6319 40426 6353
rect 40650 8223 40684 8257
rect 40650 8155 40684 8189
rect 40650 8087 40684 8121
rect 40650 8019 40684 8053
rect 40650 7951 40684 7985
rect 40650 7883 40684 7917
rect 40650 7815 40684 7849
rect 40650 7747 40684 7781
rect 40650 7679 40684 7713
rect 40650 7611 40684 7645
rect 40650 7543 40684 7577
rect 40650 7475 40684 7509
rect 40650 7407 40684 7441
rect 40650 7339 40684 7373
rect 40650 7271 40684 7305
rect 40650 7203 40684 7237
rect 40650 7135 40684 7169
rect 40650 7067 40684 7101
rect 40650 6999 40684 7033
rect 40650 6931 40684 6965
rect 40650 6863 40684 6897
rect 40650 6795 40684 6829
rect 40650 6727 40684 6761
rect 40650 6659 40684 6693
rect 40650 6591 40684 6625
rect 40650 6523 40684 6557
rect 40650 6455 40684 6489
rect 40650 6387 40684 6421
rect 40650 6319 40684 6353
rect 40908 8223 40942 8257
rect 40908 8155 40942 8189
rect 40908 8087 40942 8121
rect 40908 8019 40942 8053
rect 40908 7951 40942 7985
rect 40908 7883 40942 7917
rect 40908 7815 40942 7849
rect 40908 7747 40942 7781
rect 40908 7679 40942 7713
rect 40908 7611 40942 7645
rect 40908 7543 40942 7577
rect 40908 7475 40942 7509
rect 40908 7407 40942 7441
rect 40908 7339 40942 7373
rect 40908 7271 40942 7305
rect 40908 7203 40942 7237
rect 40908 7135 40942 7169
rect 40908 7067 40942 7101
rect 40908 6999 40942 7033
rect 40908 6931 40942 6965
rect 40908 6863 40942 6897
rect 40908 6795 40942 6829
rect 40908 6727 40942 6761
rect 40908 6659 40942 6693
rect 40908 6591 40942 6625
rect 40908 6523 40942 6557
rect 40908 6455 40942 6489
rect 40908 6387 40942 6421
rect 40908 6319 40942 6353
rect 41166 8223 41200 8257
rect 41166 8155 41200 8189
rect 41166 8087 41200 8121
rect 41166 8019 41200 8053
rect 41166 7951 41200 7985
rect 41166 7883 41200 7917
rect 41166 7815 41200 7849
rect 41166 7747 41200 7781
rect 41166 7679 41200 7713
rect 41166 7611 41200 7645
rect 41166 7543 41200 7577
rect 41166 7475 41200 7509
rect 41166 7407 41200 7441
rect 41166 7339 41200 7373
rect 41166 7271 41200 7305
rect 41166 7203 41200 7237
rect 41166 7135 41200 7169
rect 41166 7067 41200 7101
rect 41166 6999 41200 7033
rect 41166 6931 41200 6965
rect 41166 6863 41200 6897
rect 41166 6795 41200 6829
rect 41166 6727 41200 6761
rect 41166 6659 41200 6693
rect 41166 6591 41200 6625
rect 41166 6523 41200 6557
rect 41166 6455 41200 6489
rect 41166 6387 41200 6421
rect 41166 6319 41200 6353
rect 41424 8223 41458 8257
rect 41424 8155 41458 8189
rect 41424 8087 41458 8121
rect 41424 8019 41458 8053
rect 41424 7951 41458 7985
rect 41424 7883 41458 7917
rect 41424 7815 41458 7849
rect 41424 7747 41458 7781
rect 41424 7679 41458 7713
rect 41424 7611 41458 7645
rect 41424 7543 41458 7577
rect 41424 7475 41458 7509
rect 41424 7407 41458 7441
rect 41424 7339 41458 7373
rect 41424 7271 41458 7305
rect 41424 7203 41458 7237
rect 41424 7135 41458 7169
rect 41424 7067 41458 7101
rect 41424 6999 41458 7033
rect 41424 6931 41458 6965
rect 41424 6863 41458 6897
rect 41424 6795 41458 6829
rect 41424 6727 41458 6761
rect 41424 6659 41458 6693
rect 41424 6591 41458 6625
rect 41424 6523 41458 6557
rect 41424 6455 41458 6489
rect 41424 6387 41458 6421
rect 41424 6319 41458 6353
rect 41682 8223 41716 8257
rect 41682 8155 41716 8189
rect 41682 8087 41716 8121
rect 41682 8019 41716 8053
rect 41682 7951 41716 7985
rect 41682 7883 41716 7917
rect 41682 7815 41716 7849
rect 41682 7747 41716 7781
rect 41682 7679 41716 7713
rect 41682 7611 41716 7645
rect 41682 7543 41716 7577
rect 41682 7475 41716 7509
rect 41682 7407 41716 7441
rect 41682 7339 41716 7373
rect 41682 7271 41716 7305
rect 41682 7203 41716 7237
rect 41682 7135 41716 7169
rect 41682 7067 41716 7101
rect 41682 6999 41716 7033
rect 41682 6931 41716 6965
rect 41682 6863 41716 6897
rect 41682 6795 41716 6829
rect 41682 6727 41716 6761
rect 41682 6659 41716 6693
rect 41682 6591 41716 6625
rect 41682 6523 41716 6557
rect 41682 6455 41716 6489
rect 41682 6387 41716 6421
rect 41682 6319 41716 6353
rect 41940 8223 41974 8257
rect 41940 8155 41974 8189
rect 41940 8087 41974 8121
rect 41940 8019 41974 8053
rect 41940 7951 41974 7985
rect 41940 7883 41974 7917
rect 41940 7815 41974 7849
rect 41940 7747 41974 7781
rect 41940 7679 41974 7713
rect 41940 7611 41974 7645
rect 41940 7543 41974 7577
rect 41940 7475 41974 7509
rect 41940 7407 41974 7441
rect 41940 7339 41974 7373
rect 41940 7271 41974 7305
rect 41940 7203 41974 7237
rect 41940 7135 41974 7169
rect 41940 7067 41974 7101
rect 41940 6999 41974 7033
rect 41940 6931 41974 6965
rect 41940 6863 41974 6897
rect 41940 6795 41974 6829
rect 41940 6727 41974 6761
rect 41940 6659 41974 6693
rect 41940 6591 41974 6625
rect 41940 6523 41974 6557
rect 41940 6455 41974 6489
rect 41940 6387 41974 6421
rect 41940 6319 41974 6353
<< mvpdiffc >>
rect -6448 17149 -6414 17183
rect -6448 17081 -6414 17115
rect -6448 17013 -6414 17047
rect -6448 16945 -6414 16979
rect -6448 16877 -6414 16911
rect -6448 16809 -6414 16843
rect -6448 16741 -6414 16775
rect -6448 16673 -6414 16707
rect -6448 16605 -6414 16639
rect -6448 16537 -6414 16571
rect -6448 16469 -6414 16503
rect -6448 16401 -6414 16435
rect -6448 16333 -6414 16367
rect -6448 16265 -6414 16299
rect -6190 17149 -6156 17183
rect -6190 17081 -6156 17115
rect -6190 17013 -6156 17047
rect -6190 16945 -6156 16979
rect -6190 16877 -6156 16911
rect -6190 16809 -6156 16843
rect -6190 16741 -6156 16775
rect -6190 16673 -6156 16707
rect -6190 16605 -6156 16639
rect -6190 16537 -6156 16571
rect -6190 16469 -6156 16503
rect -6190 16401 -6156 16435
rect -6190 16333 -6156 16367
rect -6190 16265 -6156 16299
rect -5932 17149 -5898 17183
rect -5932 17081 -5898 17115
rect -5932 17013 -5898 17047
rect -5932 16945 -5898 16979
rect -5932 16877 -5898 16911
rect -5932 16809 -5898 16843
rect -5932 16741 -5898 16775
rect -5932 16673 -5898 16707
rect -5932 16605 -5898 16639
rect -5932 16537 -5898 16571
rect -5932 16469 -5898 16503
rect -5932 16401 -5898 16435
rect -5932 16333 -5898 16367
rect -5932 16265 -5898 16299
rect -2980 18028 -2946 18062
rect -2980 17960 -2946 17994
rect -2980 17892 -2946 17926
rect -2980 17824 -2946 17858
rect -2980 17756 -2946 17790
rect -2980 17688 -2946 17722
rect -2980 17620 -2946 17654
rect -2980 17552 -2946 17586
rect -2980 17484 -2946 17518
rect -2980 17416 -2946 17450
rect -2980 17348 -2946 17382
rect -2980 17280 -2946 17314
rect -2980 17212 -2946 17246
rect -2980 17144 -2946 17178
rect -2980 17076 -2946 17110
rect -2980 17008 -2946 17042
rect -2980 16940 -2946 16974
rect -2980 16872 -2946 16906
rect -2980 16804 -2946 16838
rect -2980 16736 -2946 16770
rect -2980 16668 -2946 16702
rect -2980 16600 -2946 16634
rect -2980 16532 -2946 16566
rect -2980 16464 -2946 16498
rect -2980 16396 -2946 16430
rect -2980 16328 -2946 16362
rect -2980 16260 -2946 16294
rect -2980 16192 -2946 16226
rect -2980 16124 -2946 16158
rect -2722 18028 -2688 18062
rect -2722 17960 -2688 17994
rect -2722 17892 -2688 17926
rect -2722 17824 -2688 17858
rect -2722 17756 -2688 17790
rect -2722 17688 -2688 17722
rect -2722 17620 -2688 17654
rect -2722 17552 -2688 17586
rect -2722 17484 -2688 17518
rect -2722 17416 -2688 17450
rect -2722 17348 -2688 17382
rect -2722 17280 -2688 17314
rect -2722 17212 -2688 17246
rect -2722 17144 -2688 17178
rect -2722 17076 -2688 17110
rect -2722 17008 -2688 17042
rect -2722 16940 -2688 16974
rect -2722 16872 -2688 16906
rect -2722 16804 -2688 16838
rect -2722 16736 -2688 16770
rect -2722 16668 -2688 16702
rect -2722 16600 -2688 16634
rect -2722 16532 -2688 16566
rect -2722 16464 -2688 16498
rect -2722 16396 -2688 16430
rect -2722 16328 -2688 16362
rect -2722 16260 -2688 16294
rect -2722 16192 -2688 16226
rect -2722 16124 -2688 16158
rect -2464 18028 -2430 18062
rect -2464 17960 -2430 17994
rect -2464 17892 -2430 17926
rect -2464 17824 -2430 17858
rect -2464 17756 -2430 17790
rect -2464 17688 -2430 17722
rect -2464 17620 -2430 17654
rect -2464 17552 -2430 17586
rect -2464 17484 -2430 17518
rect -2464 17416 -2430 17450
rect -2464 17348 -2430 17382
rect -2464 17280 -2430 17314
rect -2464 17212 -2430 17246
rect -2464 17144 -2430 17178
rect -2464 17076 -2430 17110
rect -2464 17008 -2430 17042
rect -2464 16940 -2430 16974
rect -2464 16872 -2430 16906
rect -2464 16804 -2430 16838
rect -2464 16736 -2430 16770
rect -2464 16668 -2430 16702
rect -2464 16600 -2430 16634
rect -2464 16532 -2430 16566
rect -2464 16464 -2430 16498
rect -2464 16396 -2430 16430
rect -2464 16328 -2430 16362
rect -2464 16260 -2430 16294
rect -2464 16192 -2430 16226
rect -2464 16124 -2430 16158
rect -2206 18028 -2172 18062
rect -2206 17960 -2172 17994
rect -2206 17892 -2172 17926
rect -2206 17824 -2172 17858
rect -2206 17756 -2172 17790
rect -2206 17688 -2172 17722
rect -2206 17620 -2172 17654
rect -2206 17552 -2172 17586
rect -2206 17484 -2172 17518
rect -2206 17416 -2172 17450
rect -2206 17348 -2172 17382
rect -2206 17280 -2172 17314
rect -2206 17212 -2172 17246
rect -2206 17144 -2172 17178
rect -2206 17076 -2172 17110
rect -2206 17008 -2172 17042
rect -2206 16940 -2172 16974
rect -2206 16872 -2172 16906
rect -2206 16804 -2172 16838
rect -2206 16736 -2172 16770
rect -2206 16668 -2172 16702
rect -2206 16600 -2172 16634
rect -2206 16532 -2172 16566
rect -2206 16464 -2172 16498
rect -2206 16396 -2172 16430
rect -2206 16328 -2172 16362
rect -2206 16260 -2172 16294
rect -2206 16192 -2172 16226
rect -2206 16124 -2172 16158
rect -1948 18028 -1914 18062
rect -1948 17960 -1914 17994
rect -1948 17892 -1914 17926
rect -1948 17824 -1914 17858
rect -1948 17756 -1914 17790
rect -1948 17688 -1914 17722
rect -1948 17620 -1914 17654
rect -1948 17552 -1914 17586
rect -1948 17484 -1914 17518
rect -1948 17416 -1914 17450
rect -1948 17348 -1914 17382
rect -1948 17280 -1914 17314
rect -1948 17212 -1914 17246
rect -1948 17144 -1914 17178
rect -1948 17076 -1914 17110
rect -1948 17008 -1914 17042
rect -1948 16940 -1914 16974
rect -1948 16872 -1914 16906
rect -1948 16804 -1914 16838
rect -1948 16736 -1914 16770
rect -1948 16668 -1914 16702
rect -1948 16600 -1914 16634
rect -1948 16532 -1914 16566
rect -1948 16464 -1914 16498
rect -1948 16396 -1914 16430
rect -1948 16328 -1914 16362
rect -1948 16260 -1914 16294
rect -1948 16192 -1914 16226
rect -1948 16124 -1914 16158
rect -1690 18028 -1656 18062
rect -1690 17960 -1656 17994
rect -1690 17892 -1656 17926
rect -1690 17824 -1656 17858
rect -1690 17756 -1656 17790
rect -1690 17688 -1656 17722
rect -1690 17620 -1656 17654
rect -1690 17552 -1656 17586
rect -1690 17484 -1656 17518
rect -1690 17416 -1656 17450
rect -1690 17348 -1656 17382
rect -1690 17280 -1656 17314
rect -1690 17212 -1656 17246
rect -1690 17144 -1656 17178
rect -1690 17076 -1656 17110
rect -1690 17008 -1656 17042
rect -1690 16940 -1656 16974
rect -1690 16872 -1656 16906
rect -1690 16804 -1656 16838
rect -1690 16736 -1656 16770
rect -1690 16668 -1656 16702
rect -1690 16600 -1656 16634
rect -1690 16532 -1656 16566
rect -1690 16464 -1656 16498
rect -1690 16396 -1656 16430
rect -1690 16328 -1656 16362
rect -1690 16260 -1656 16294
rect -1690 16192 -1656 16226
rect -1690 16124 -1656 16158
rect -1432 18028 -1398 18062
rect -1432 17960 -1398 17994
rect -1432 17892 -1398 17926
rect -1432 17824 -1398 17858
rect -1432 17756 -1398 17790
rect -1432 17688 -1398 17722
rect -1432 17620 -1398 17654
rect -1432 17552 -1398 17586
rect -1432 17484 -1398 17518
rect -1432 17416 -1398 17450
rect -1432 17348 -1398 17382
rect -1432 17280 -1398 17314
rect -1432 17212 -1398 17246
rect -1432 17144 -1398 17178
rect -1432 17076 -1398 17110
rect -1432 17008 -1398 17042
rect -1432 16940 -1398 16974
rect -1432 16872 -1398 16906
rect -1432 16804 -1398 16838
rect -1432 16736 -1398 16770
rect -1432 16668 -1398 16702
rect -1432 16600 -1398 16634
rect -1432 16532 -1398 16566
rect -1432 16464 -1398 16498
rect -1432 16396 -1398 16430
rect -1432 16328 -1398 16362
rect -1432 16260 -1398 16294
rect -1432 16192 -1398 16226
rect -1432 16124 -1398 16158
rect -1174 18028 -1140 18062
rect -1174 17960 -1140 17994
rect -1174 17892 -1140 17926
rect -1174 17824 -1140 17858
rect -1174 17756 -1140 17790
rect -1174 17688 -1140 17722
rect -1174 17620 -1140 17654
rect -1174 17552 -1140 17586
rect -1174 17484 -1140 17518
rect -1174 17416 -1140 17450
rect -1174 17348 -1140 17382
rect -1174 17280 -1140 17314
rect -1174 17212 -1140 17246
rect -1174 17144 -1140 17178
rect -1174 17076 -1140 17110
rect -1174 17008 -1140 17042
rect -1174 16940 -1140 16974
rect -1174 16872 -1140 16906
rect -1174 16804 -1140 16838
rect -1174 16736 -1140 16770
rect -1174 16668 -1140 16702
rect -1174 16600 -1140 16634
rect -1174 16532 -1140 16566
rect -1174 16464 -1140 16498
rect -1174 16396 -1140 16430
rect -1174 16328 -1140 16362
rect -1174 16260 -1140 16294
rect -1174 16192 -1140 16226
rect -1174 16124 -1140 16158
rect -916 18028 -882 18062
rect -916 17960 -882 17994
rect -916 17892 -882 17926
rect -916 17824 -882 17858
rect -916 17756 -882 17790
rect -916 17688 -882 17722
rect -916 17620 -882 17654
rect -916 17552 -882 17586
rect -916 17484 -882 17518
rect -916 17416 -882 17450
rect -916 17348 -882 17382
rect -916 17280 -882 17314
rect -916 17212 -882 17246
rect -916 17144 -882 17178
rect -916 17076 -882 17110
rect -916 17008 -882 17042
rect -916 16940 -882 16974
rect -916 16872 -882 16906
rect -916 16804 -882 16838
rect -916 16736 -882 16770
rect -916 16668 -882 16702
rect -916 16600 -882 16634
rect -916 16532 -882 16566
rect -916 16464 -882 16498
rect -916 16396 -882 16430
rect -916 16328 -882 16362
rect -916 16260 -882 16294
rect -916 16192 -882 16226
rect -916 16124 -882 16158
rect -658 18028 -624 18062
rect -658 17960 -624 17994
rect -658 17892 -624 17926
rect -658 17824 -624 17858
rect -658 17756 -624 17790
rect -658 17688 -624 17722
rect -658 17620 -624 17654
rect -658 17552 -624 17586
rect -658 17484 -624 17518
rect -658 17416 -624 17450
rect -658 17348 -624 17382
rect -658 17280 -624 17314
rect -658 17212 -624 17246
rect -658 17144 -624 17178
rect -658 17076 -624 17110
rect -658 17008 -624 17042
rect -658 16940 -624 16974
rect -658 16872 -624 16906
rect -658 16804 -624 16838
rect -658 16736 -624 16770
rect -658 16668 -624 16702
rect -658 16600 -624 16634
rect -658 16532 -624 16566
rect -658 16464 -624 16498
rect -658 16396 -624 16430
rect -658 16328 -624 16362
rect -658 16260 -624 16294
rect -658 16192 -624 16226
rect -658 16124 -624 16158
rect -400 18028 -366 18062
rect -400 17960 -366 17994
rect -400 17892 -366 17926
rect -400 17824 -366 17858
rect -400 17756 -366 17790
rect -400 17688 -366 17722
rect -400 17620 -366 17654
rect -400 17552 -366 17586
rect -400 17484 -366 17518
rect -400 17416 -366 17450
rect -400 17348 -366 17382
rect -400 17280 -366 17314
rect -400 17212 -366 17246
rect -400 17144 -366 17178
rect -400 17076 -366 17110
rect -400 17008 -366 17042
rect -400 16940 -366 16974
rect -400 16872 -366 16906
rect -400 16804 -366 16838
rect -400 16736 -366 16770
rect -400 16668 -366 16702
rect -400 16600 -366 16634
rect -400 16532 -366 16566
rect -400 16464 -366 16498
rect -400 16396 -366 16430
rect -400 16328 -366 16362
rect -400 16260 -366 16294
rect -400 16192 -366 16226
rect -400 16124 -366 16158
rect 23176 18672 23210 18706
rect 23176 18604 23210 18638
rect 23176 18536 23210 18570
rect 23176 18468 23210 18502
rect 23176 18400 23210 18434
rect 23176 18332 23210 18366
rect 23176 18264 23210 18298
rect 23176 18196 23210 18230
rect 23176 18128 23210 18162
rect 23176 18060 23210 18094
rect 23176 17992 23210 18026
rect 23176 17924 23210 17958
rect 23176 17856 23210 17890
rect 23176 17788 23210 17822
rect 24234 18672 24268 18706
rect 24234 18604 24268 18638
rect 24234 18536 24268 18570
rect 24234 18468 24268 18502
rect 24234 18400 24268 18434
rect 24234 18332 24268 18366
rect 24234 18264 24268 18298
rect 24234 18196 24268 18230
rect 24234 18128 24268 18162
rect 24234 18060 24268 18094
rect 24234 17992 24268 18026
rect 24234 17924 24268 17958
rect 24234 17856 24268 17890
rect 24234 17788 24268 17822
rect 24692 18678 24726 18712
rect 24692 18610 24726 18644
rect 24692 18542 24726 18576
rect 24692 18474 24726 18508
rect 24692 18406 24726 18440
rect 24692 18338 24726 18372
rect 24692 18270 24726 18304
rect 24692 18202 24726 18236
rect 24692 18134 24726 18168
rect 24692 18066 24726 18100
rect 24692 17998 24726 18032
rect 24692 17930 24726 17964
rect 24692 17862 24726 17896
rect 24692 17794 24726 17828
rect 24692 17726 24726 17760
rect 24692 17658 24726 17692
rect 24692 17590 24726 17624
rect 24692 17522 24726 17556
rect 24692 17454 24726 17488
rect 24692 17386 24726 17420
rect 24692 17318 24726 17352
rect 24692 17250 24726 17284
rect 24692 17182 24726 17216
rect 25750 18678 25784 18712
rect 25750 18610 25784 18644
rect 25750 18542 25784 18576
rect 25750 18474 25784 18508
rect 25750 18406 25784 18440
rect 25750 18338 25784 18372
rect 25750 18270 25784 18304
rect 25750 18202 25784 18236
rect 25750 18134 25784 18168
rect 25750 18066 25784 18100
rect 25750 17998 25784 18032
rect 25750 17930 25784 17964
rect 25750 17862 25784 17896
rect 25750 17794 25784 17828
rect 25750 17726 25784 17760
rect 25750 17658 25784 17692
rect 25750 17590 25784 17624
rect 25750 17522 25784 17556
rect 25750 17454 25784 17488
rect 25750 17386 25784 17420
rect 25750 17318 25784 17352
rect 25750 17250 25784 17284
rect 25750 17182 25784 17216
rect 26808 18678 26842 18712
rect 26808 18610 26842 18644
rect 26808 18542 26842 18576
rect 26808 18474 26842 18508
rect 26808 18406 26842 18440
rect 26808 18338 26842 18372
rect 26808 18270 26842 18304
rect 26808 18202 26842 18236
rect 26808 18134 26842 18168
rect 26808 18066 26842 18100
rect 26808 17998 26842 18032
rect 26808 17930 26842 17964
rect 26808 17862 26842 17896
rect 26808 17794 26842 17828
rect 26808 17726 26842 17760
rect 26808 17658 26842 17692
rect 26808 17590 26842 17624
rect 26808 17522 26842 17556
rect 26808 17454 26842 17488
rect 26808 17386 26842 17420
rect 26808 17318 26842 17352
rect 26808 17250 26842 17284
rect 26808 17182 26842 17216
rect 27866 18678 27900 18712
rect 27866 18610 27900 18644
rect 27866 18542 27900 18576
rect 27866 18474 27900 18508
rect 27866 18406 27900 18440
rect 27866 18338 27900 18372
rect 27866 18270 27900 18304
rect 27866 18202 27900 18236
rect 27866 18134 27900 18168
rect 27866 18066 27900 18100
rect 27866 17998 27900 18032
rect 27866 17930 27900 17964
rect 27866 17862 27900 17896
rect 27866 17794 27900 17828
rect 27866 17726 27900 17760
rect 27866 17658 27900 17692
rect 27866 17590 27900 17624
rect 27866 17522 27900 17556
rect 27866 17454 27900 17488
rect 27866 17386 27900 17420
rect 27866 17318 27900 17352
rect 27866 17250 27900 17284
rect 27866 17182 27900 17216
rect 39144 17899 39178 17933
rect 39144 17831 39178 17865
rect 39144 17763 39178 17797
rect 39144 17695 39178 17729
rect 39144 17627 39178 17661
rect 39144 17559 39178 17593
rect 39144 17491 39178 17525
rect 39144 17423 39178 17457
rect 39144 17355 39178 17389
rect 39144 17287 39178 17321
rect 39144 17219 39178 17253
rect 39144 17151 39178 17185
rect 39144 17083 39178 17117
rect 39144 17015 39178 17049
rect 39402 17899 39436 17933
rect 39402 17831 39436 17865
rect 39402 17763 39436 17797
rect 39402 17695 39436 17729
rect 39402 17627 39436 17661
rect 39402 17559 39436 17593
rect 39402 17491 39436 17525
rect 39402 17423 39436 17457
rect 39402 17355 39436 17389
rect 39402 17287 39436 17321
rect 39402 17219 39436 17253
rect 39402 17151 39436 17185
rect 39402 17083 39436 17117
rect 39402 17015 39436 17049
rect 39660 17899 39694 17933
rect 39660 17831 39694 17865
rect 39660 17763 39694 17797
rect 39660 17695 39694 17729
rect 39660 17627 39694 17661
rect 39660 17559 39694 17593
rect 39660 17491 39694 17525
rect 39660 17423 39694 17457
rect 39660 17355 39694 17389
rect 39660 17287 39694 17321
rect 39660 17219 39694 17253
rect 39660 17151 39694 17185
rect 39660 17083 39694 17117
rect 39660 17015 39694 17049
rect 42612 18778 42646 18812
rect 42612 18710 42646 18744
rect 42612 18642 42646 18676
rect 42612 18574 42646 18608
rect 42612 18506 42646 18540
rect 42612 18438 42646 18472
rect 42612 18370 42646 18404
rect 42612 18302 42646 18336
rect 42612 18234 42646 18268
rect 42612 18166 42646 18200
rect 42612 18098 42646 18132
rect 42612 18030 42646 18064
rect 42612 17962 42646 17996
rect 42612 17894 42646 17928
rect 42612 17826 42646 17860
rect 42612 17758 42646 17792
rect 42612 17690 42646 17724
rect 42612 17622 42646 17656
rect 42612 17554 42646 17588
rect 42612 17486 42646 17520
rect 42612 17418 42646 17452
rect 42612 17350 42646 17384
rect 42612 17282 42646 17316
rect 42612 17214 42646 17248
rect 42612 17146 42646 17180
rect 42612 17078 42646 17112
rect 42612 17010 42646 17044
rect 42612 16942 42646 16976
rect 42612 16874 42646 16908
rect 42870 18778 42904 18812
rect 42870 18710 42904 18744
rect 42870 18642 42904 18676
rect 42870 18574 42904 18608
rect 42870 18506 42904 18540
rect 42870 18438 42904 18472
rect 42870 18370 42904 18404
rect 42870 18302 42904 18336
rect 42870 18234 42904 18268
rect 42870 18166 42904 18200
rect 42870 18098 42904 18132
rect 42870 18030 42904 18064
rect 42870 17962 42904 17996
rect 42870 17894 42904 17928
rect 42870 17826 42904 17860
rect 42870 17758 42904 17792
rect 42870 17690 42904 17724
rect 42870 17622 42904 17656
rect 42870 17554 42904 17588
rect 42870 17486 42904 17520
rect 42870 17418 42904 17452
rect 42870 17350 42904 17384
rect 42870 17282 42904 17316
rect 42870 17214 42904 17248
rect 42870 17146 42904 17180
rect 42870 17078 42904 17112
rect 42870 17010 42904 17044
rect 42870 16942 42904 16976
rect 42870 16874 42904 16908
rect 43128 18778 43162 18812
rect 43128 18710 43162 18744
rect 43128 18642 43162 18676
rect 43128 18574 43162 18608
rect 43128 18506 43162 18540
rect 43128 18438 43162 18472
rect 43128 18370 43162 18404
rect 43128 18302 43162 18336
rect 43128 18234 43162 18268
rect 43128 18166 43162 18200
rect 43128 18098 43162 18132
rect 43128 18030 43162 18064
rect 43128 17962 43162 17996
rect 43128 17894 43162 17928
rect 43128 17826 43162 17860
rect 43128 17758 43162 17792
rect 43128 17690 43162 17724
rect 43128 17622 43162 17656
rect 43128 17554 43162 17588
rect 43128 17486 43162 17520
rect 43128 17418 43162 17452
rect 43128 17350 43162 17384
rect 43128 17282 43162 17316
rect 43128 17214 43162 17248
rect 43128 17146 43162 17180
rect 43128 17078 43162 17112
rect 43128 17010 43162 17044
rect 43128 16942 43162 16976
rect 43128 16874 43162 16908
rect 43386 18778 43420 18812
rect 43386 18710 43420 18744
rect 43386 18642 43420 18676
rect 43386 18574 43420 18608
rect 43386 18506 43420 18540
rect 43386 18438 43420 18472
rect 43386 18370 43420 18404
rect 43386 18302 43420 18336
rect 43386 18234 43420 18268
rect 43386 18166 43420 18200
rect 43386 18098 43420 18132
rect 43386 18030 43420 18064
rect 43386 17962 43420 17996
rect 43386 17894 43420 17928
rect 43386 17826 43420 17860
rect 43386 17758 43420 17792
rect 43386 17690 43420 17724
rect 43386 17622 43420 17656
rect 43386 17554 43420 17588
rect 43386 17486 43420 17520
rect 43386 17418 43420 17452
rect 43386 17350 43420 17384
rect 43386 17282 43420 17316
rect 43386 17214 43420 17248
rect 43386 17146 43420 17180
rect 43386 17078 43420 17112
rect 43386 17010 43420 17044
rect 43386 16942 43420 16976
rect 43386 16874 43420 16908
rect 43644 18778 43678 18812
rect 43644 18710 43678 18744
rect 43644 18642 43678 18676
rect 43644 18574 43678 18608
rect 43644 18506 43678 18540
rect 43644 18438 43678 18472
rect 43644 18370 43678 18404
rect 43644 18302 43678 18336
rect 43644 18234 43678 18268
rect 43644 18166 43678 18200
rect 43644 18098 43678 18132
rect 43644 18030 43678 18064
rect 43644 17962 43678 17996
rect 43644 17894 43678 17928
rect 43644 17826 43678 17860
rect 43644 17758 43678 17792
rect 43644 17690 43678 17724
rect 43644 17622 43678 17656
rect 43644 17554 43678 17588
rect 43644 17486 43678 17520
rect 43644 17418 43678 17452
rect 43644 17350 43678 17384
rect 43644 17282 43678 17316
rect 43644 17214 43678 17248
rect 43644 17146 43678 17180
rect 43644 17078 43678 17112
rect 43644 17010 43678 17044
rect 43644 16942 43678 16976
rect 43644 16874 43678 16908
rect 43902 18778 43936 18812
rect 43902 18710 43936 18744
rect 43902 18642 43936 18676
rect 43902 18574 43936 18608
rect 43902 18506 43936 18540
rect 43902 18438 43936 18472
rect 43902 18370 43936 18404
rect 43902 18302 43936 18336
rect 43902 18234 43936 18268
rect 43902 18166 43936 18200
rect 43902 18098 43936 18132
rect 43902 18030 43936 18064
rect 43902 17962 43936 17996
rect 43902 17894 43936 17928
rect 43902 17826 43936 17860
rect 43902 17758 43936 17792
rect 43902 17690 43936 17724
rect 43902 17622 43936 17656
rect 43902 17554 43936 17588
rect 43902 17486 43936 17520
rect 43902 17418 43936 17452
rect 43902 17350 43936 17384
rect 43902 17282 43936 17316
rect 43902 17214 43936 17248
rect 43902 17146 43936 17180
rect 43902 17078 43936 17112
rect 43902 17010 43936 17044
rect 43902 16942 43936 16976
rect 43902 16874 43936 16908
rect 44160 18778 44194 18812
rect 44160 18710 44194 18744
rect 44160 18642 44194 18676
rect 44160 18574 44194 18608
rect 44160 18506 44194 18540
rect 44160 18438 44194 18472
rect 44160 18370 44194 18404
rect 44160 18302 44194 18336
rect 44160 18234 44194 18268
rect 44160 18166 44194 18200
rect 44160 18098 44194 18132
rect 44160 18030 44194 18064
rect 44160 17962 44194 17996
rect 44160 17894 44194 17928
rect 44160 17826 44194 17860
rect 44160 17758 44194 17792
rect 44160 17690 44194 17724
rect 44160 17622 44194 17656
rect 44160 17554 44194 17588
rect 44160 17486 44194 17520
rect 44160 17418 44194 17452
rect 44160 17350 44194 17384
rect 44160 17282 44194 17316
rect 44160 17214 44194 17248
rect 44160 17146 44194 17180
rect 44160 17078 44194 17112
rect 44160 17010 44194 17044
rect 44160 16942 44194 16976
rect 44160 16874 44194 16908
rect 44418 18778 44452 18812
rect 44418 18710 44452 18744
rect 44418 18642 44452 18676
rect 44418 18574 44452 18608
rect 44418 18506 44452 18540
rect 44418 18438 44452 18472
rect 44418 18370 44452 18404
rect 44418 18302 44452 18336
rect 44418 18234 44452 18268
rect 44418 18166 44452 18200
rect 44418 18098 44452 18132
rect 44418 18030 44452 18064
rect 44418 17962 44452 17996
rect 44418 17894 44452 17928
rect 44418 17826 44452 17860
rect 44418 17758 44452 17792
rect 44418 17690 44452 17724
rect 44418 17622 44452 17656
rect 44418 17554 44452 17588
rect 44418 17486 44452 17520
rect 44418 17418 44452 17452
rect 44418 17350 44452 17384
rect 44418 17282 44452 17316
rect 44418 17214 44452 17248
rect 44418 17146 44452 17180
rect 44418 17078 44452 17112
rect 44418 17010 44452 17044
rect 44418 16942 44452 16976
rect 44418 16874 44452 16908
rect 44676 18778 44710 18812
rect 44676 18710 44710 18744
rect 44676 18642 44710 18676
rect 44676 18574 44710 18608
rect 44676 18506 44710 18540
rect 44676 18438 44710 18472
rect 44676 18370 44710 18404
rect 44676 18302 44710 18336
rect 44676 18234 44710 18268
rect 44676 18166 44710 18200
rect 44676 18098 44710 18132
rect 44676 18030 44710 18064
rect 44676 17962 44710 17996
rect 44676 17894 44710 17928
rect 44676 17826 44710 17860
rect 44676 17758 44710 17792
rect 44676 17690 44710 17724
rect 44676 17622 44710 17656
rect 44676 17554 44710 17588
rect 44676 17486 44710 17520
rect 44676 17418 44710 17452
rect 44676 17350 44710 17384
rect 44676 17282 44710 17316
rect 44676 17214 44710 17248
rect 44676 17146 44710 17180
rect 44676 17078 44710 17112
rect 44676 17010 44710 17044
rect 44676 16942 44710 16976
rect 44676 16874 44710 16908
rect 44934 18778 44968 18812
rect 44934 18710 44968 18744
rect 44934 18642 44968 18676
rect 44934 18574 44968 18608
rect 44934 18506 44968 18540
rect 44934 18438 44968 18472
rect 44934 18370 44968 18404
rect 44934 18302 44968 18336
rect 44934 18234 44968 18268
rect 44934 18166 44968 18200
rect 44934 18098 44968 18132
rect 44934 18030 44968 18064
rect 44934 17962 44968 17996
rect 44934 17894 44968 17928
rect 44934 17826 44968 17860
rect 44934 17758 44968 17792
rect 44934 17690 44968 17724
rect 44934 17622 44968 17656
rect 44934 17554 44968 17588
rect 44934 17486 44968 17520
rect 44934 17418 44968 17452
rect 44934 17350 44968 17384
rect 44934 17282 44968 17316
rect 44934 17214 44968 17248
rect 44934 17146 44968 17180
rect 44934 17078 44968 17112
rect 44934 17010 44968 17044
rect 44934 16942 44968 16976
rect 44934 16874 44968 16908
rect 45192 18778 45226 18812
rect 45192 18710 45226 18744
rect 45192 18642 45226 18676
rect 45192 18574 45226 18608
rect 45192 18506 45226 18540
rect 45192 18438 45226 18472
rect 45192 18370 45226 18404
rect 45192 18302 45226 18336
rect 45192 18234 45226 18268
rect 45192 18166 45226 18200
rect 45192 18098 45226 18132
rect 45192 18030 45226 18064
rect 45192 17962 45226 17996
rect 45192 17894 45226 17928
rect 45192 17826 45226 17860
rect 45192 17758 45226 17792
rect 45192 17690 45226 17724
rect 45192 17622 45226 17656
rect 45192 17554 45226 17588
rect 45192 17486 45226 17520
rect 45192 17418 45226 17452
rect 45192 17350 45226 17384
rect 45192 17282 45226 17316
rect 45192 17214 45226 17248
rect 45192 17146 45226 17180
rect 45192 17078 45226 17112
rect 45192 17010 45226 17044
rect 45192 16942 45226 16976
rect 45192 16874 45226 16908
rect 12994 14712 13028 14746
rect 12994 14644 13028 14678
rect 12994 14576 13028 14610
rect 12994 14508 13028 14542
rect 12994 14440 13028 14474
rect 12994 14372 13028 14406
rect 12994 14304 13028 14338
rect 12994 14236 13028 14270
rect 12994 14168 13028 14202
rect 12994 14100 13028 14134
rect 12994 14032 13028 14066
rect 12994 13964 13028 13998
rect 12994 13896 13028 13930
rect 12994 13828 13028 13862
rect 12994 13760 13028 13794
rect 12994 13692 13028 13726
rect 12994 13624 13028 13658
rect 12994 13556 13028 13590
rect 12994 13488 13028 13522
rect 12994 13420 13028 13454
rect 12994 13352 13028 13386
rect 12994 13284 13028 13318
rect 12994 13216 13028 13250
rect 12994 13148 13028 13182
rect 12994 13080 13028 13114
rect 12994 13012 13028 13046
rect 12994 12944 13028 12978
rect 12994 12876 13028 12910
rect 12994 12808 13028 12842
rect 12994 12740 13028 12774
rect 12994 12672 13028 12706
rect 12994 12604 13028 12638
rect 12994 12536 13028 12570
rect 12994 12468 13028 12502
rect 12994 12400 13028 12434
rect 12994 12332 13028 12366
rect 12994 12264 13028 12298
rect 12994 12196 13028 12230
rect 12994 12128 13028 12162
rect 12994 12060 13028 12094
rect 12994 11992 13028 12026
rect 12994 11924 13028 11958
rect 12994 11856 13028 11890
rect 12994 11788 13028 11822
rect 14052 14712 14086 14746
rect 14052 14644 14086 14678
rect 14052 14576 14086 14610
rect 14052 14508 14086 14542
rect 14052 14440 14086 14474
rect 14052 14372 14086 14406
rect 14052 14304 14086 14338
rect 14052 14236 14086 14270
rect 14052 14168 14086 14202
rect 14052 14100 14086 14134
rect 14052 14032 14086 14066
rect 14052 13964 14086 13998
rect 14052 13896 14086 13930
rect 14052 13828 14086 13862
rect 14052 13760 14086 13794
rect 14052 13692 14086 13726
rect 14052 13624 14086 13658
rect 14052 13556 14086 13590
rect 14052 13488 14086 13522
rect 14052 13420 14086 13454
rect 14052 13352 14086 13386
rect 14052 13284 14086 13318
rect 14052 13216 14086 13250
rect 14052 13148 14086 13182
rect 14052 13080 14086 13114
rect 14052 13012 14086 13046
rect 14052 12944 14086 12978
rect 14052 12876 14086 12910
rect 14052 12808 14086 12842
rect 14052 12740 14086 12774
rect 14052 12672 14086 12706
rect 14052 12604 14086 12638
rect 14052 12536 14086 12570
rect 14052 12468 14086 12502
rect 14052 12400 14086 12434
rect 14052 12332 14086 12366
rect 14052 12264 14086 12298
rect 14052 12196 14086 12230
rect 14052 12128 14086 12162
rect 14052 12060 14086 12094
rect 14052 11992 14086 12026
rect 14052 11924 14086 11958
rect 14052 11856 14086 11890
rect 14052 11788 14086 11822
rect 15110 14712 15144 14746
rect 15110 14644 15144 14678
rect 15110 14576 15144 14610
rect 15110 14508 15144 14542
rect 15110 14440 15144 14474
rect 15110 14372 15144 14406
rect 15110 14304 15144 14338
rect 15110 14236 15144 14270
rect 15110 14168 15144 14202
rect 15110 14100 15144 14134
rect 15110 14032 15144 14066
rect 15110 13964 15144 13998
rect 15110 13896 15144 13930
rect 15110 13828 15144 13862
rect 15110 13760 15144 13794
rect 15110 13692 15144 13726
rect 15110 13624 15144 13658
rect 15110 13556 15144 13590
rect 15110 13488 15144 13522
rect 15110 13420 15144 13454
rect 15110 13352 15144 13386
rect 15110 13284 15144 13318
rect 15110 13216 15144 13250
rect 15110 13148 15144 13182
rect 15110 13080 15144 13114
rect 15110 13012 15144 13046
rect 15110 12944 15144 12978
rect 15110 12876 15144 12910
rect 15110 12808 15144 12842
rect 15110 12740 15144 12774
rect 15110 12672 15144 12706
rect 15110 12604 15144 12638
rect 15110 12536 15144 12570
rect 15110 12468 15144 12502
rect 15110 12400 15144 12434
rect 15110 12332 15144 12366
rect 15110 12264 15144 12298
rect 15110 12196 15144 12230
rect 15110 12128 15144 12162
rect 15110 12060 15144 12094
rect 15110 11992 15144 12026
rect 15110 11924 15144 11958
rect 15110 11856 15144 11890
rect 15110 11788 15144 11822
rect 15564 14712 15598 14746
rect 15564 14644 15598 14678
rect 15564 14576 15598 14610
rect 15564 14508 15598 14542
rect 15564 14440 15598 14474
rect 15564 14372 15598 14406
rect 15564 14304 15598 14338
rect 15564 14236 15598 14270
rect 15564 14168 15598 14202
rect 15564 14100 15598 14134
rect 15564 14032 15598 14066
rect 15564 13964 15598 13998
rect 15564 13896 15598 13930
rect 15564 13828 15598 13862
rect 15564 13760 15598 13794
rect 15564 13692 15598 13726
rect 15564 13624 15598 13658
rect 15564 13556 15598 13590
rect 15564 13488 15598 13522
rect 15564 13420 15598 13454
rect 15564 13352 15598 13386
rect 15564 13284 15598 13318
rect 15564 13216 15598 13250
rect 15564 13148 15598 13182
rect 15564 13080 15598 13114
rect 15564 13012 15598 13046
rect 15564 12944 15598 12978
rect 15564 12876 15598 12910
rect 15564 12808 15598 12842
rect 15564 12740 15598 12774
rect 15564 12672 15598 12706
rect 15564 12604 15598 12638
rect 15564 12536 15598 12570
rect 15564 12468 15598 12502
rect 15564 12400 15598 12434
rect 15564 12332 15598 12366
rect 15564 12264 15598 12298
rect 15564 12196 15598 12230
rect 15564 12128 15598 12162
rect 15564 12060 15598 12094
rect 15564 11992 15598 12026
rect 15564 11924 15598 11958
rect 15564 11856 15598 11890
rect 15564 11788 15598 11822
rect 16622 14712 16656 14746
rect 16622 14644 16656 14678
rect 16622 14576 16656 14610
rect 16622 14508 16656 14542
rect 16622 14440 16656 14474
rect 16622 14372 16656 14406
rect 16622 14304 16656 14338
rect 16622 14236 16656 14270
rect 16622 14168 16656 14202
rect 16622 14100 16656 14134
rect 16622 14032 16656 14066
rect 16622 13964 16656 13998
rect 16622 13896 16656 13930
rect 16622 13828 16656 13862
rect 16622 13760 16656 13794
rect 16622 13692 16656 13726
rect 16622 13624 16656 13658
rect 16622 13556 16656 13590
rect 16622 13488 16656 13522
rect 16622 13420 16656 13454
rect 16622 13352 16656 13386
rect 16622 13284 16656 13318
rect 16622 13216 16656 13250
rect 16622 13148 16656 13182
rect 16622 13080 16656 13114
rect 16622 13012 16656 13046
rect 16622 12944 16656 12978
rect 16622 12876 16656 12910
rect 16622 12808 16656 12842
rect 16622 12740 16656 12774
rect 16622 12672 16656 12706
rect 16622 12604 16656 12638
rect 16622 12536 16656 12570
rect 16622 12468 16656 12502
rect 16622 12400 16656 12434
rect 16622 12332 16656 12366
rect 16622 12264 16656 12298
rect 16622 12196 16656 12230
rect 16622 12128 16656 12162
rect 16622 12060 16656 12094
rect 16622 11992 16656 12026
rect 16622 11924 16656 11958
rect 16622 11856 16656 11890
rect 16622 11788 16656 11822
rect 17074 14722 17108 14756
rect 17074 14654 17108 14688
rect 17074 14586 17108 14620
rect 17074 14518 17108 14552
rect 17074 14450 17108 14484
rect 17074 14382 17108 14416
rect 17074 14314 17108 14348
rect 17074 14246 17108 14280
rect 17074 14178 17108 14212
rect 17074 14110 17108 14144
rect 17074 14042 17108 14076
rect 17074 13974 17108 14008
rect 17074 13906 17108 13940
rect 17074 13838 17108 13872
rect 17074 13770 17108 13804
rect 17074 13702 17108 13736
rect 17074 13634 17108 13668
rect 17074 13566 17108 13600
rect 17074 13498 17108 13532
rect 17074 13430 17108 13464
rect 17074 13362 17108 13396
rect 17074 13294 17108 13328
rect 17074 13226 17108 13260
rect 17074 13158 17108 13192
rect 17074 13090 17108 13124
rect 17074 13022 17108 13056
rect 17074 12954 17108 12988
rect 17074 12886 17108 12920
rect 17074 12818 17108 12852
rect 17074 12750 17108 12784
rect 17074 12682 17108 12716
rect 17074 12614 17108 12648
rect 17074 12546 17108 12580
rect 17074 12478 17108 12512
rect 17074 12410 17108 12444
rect 17074 12342 17108 12376
rect 17074 12274 17108 12308
rect 17074 12206 17108 12240
rect 17074 12138 17108 12172
rect 17074 12070 17108 12104
rect 17074 12002 17108 12036
rect 17074 11934 17108 11968
rect 17074 11866 17108 11900
rect 17074 11798 17108 11832
rect 18132 14722 18166 14756
rect 18132 14654 18166 14688
rect 18132 14586 18166 14620
rect 18132 14518 18166 14552
rect 18132 14450 18166 14484
rect 18132 14382 18166 14416
rect 18132 14314 18166 14348
rect 18132 14246 18166 14280
rect 18132 14178 18166 14212
rect 18132 14110 18166 14144
rect 18132 14042 18166 14076
rect 18132 13974 18166 14008
rect 18132 13906 18166 13940
rect 18132 13838 18166 13872
rect 18132 13770 18166 13804
rect 18132 13702 18166 13736
rect 18132 13634 18166 13668
rect 18132 13566 18166 13600
rect 18132 13498 18166 13532
rect 18132 13430 18166 13464
rect 18132 13362 18166 13396
rect 18132 13294 18166 13328
rect 18132 13226 18166 13260
rect 18132 13158 18166 13192
rect 18132 13090 18166 13124
rect 18132 13022 18166 13056
rect 18132 12954 18166 12988
rect 18132 12886 18166 12920
rect 18132 12818 18166 12852
rect 18132 12750 18166 12784
rect 18132 12682 18166 12716
rect 18132 12614 18166 12648
rect 18132 12546 18166 12580
rect 18132 12478 18166 12512
rect 18132 12410 18166 12444
rect 18132 12342 18166 12376
rect 18132 12274 18166 12308
rect 18132 12206 18166 12240
rect 18132 12138 18166 12172
rect 18132 12070 18166 12104
rect 18132 12002 18166 12036
rect 18132 11934 18166 11968
rect 18132 11866 18166 11900
rect 18132 11798 18166 11832
rect 18538 14706 18572 14740
rect 18538 14638 18572 14672
rect 18538 14570 18572 14604
rect 18538 14502 18572 14536
rect 18538 14434 18572 14468
rect 18538 14366 18572 14400
rect 18538 14298 18572 14332
rect 18538 14230 18572 14264
rect 18538 14162 18572 14196
rect 18538 14094 18572 14128
rect 18538 14026 18572 14060
rect 18538 13958 18572 13992
rect 18538 13890 18572 13924
rect 18538 13822 18572 13856
rect 18538 13754 18572 13788
rect 18538 13686 18572 13720
rect 18538 13618 18572 13652
rect 18538 13550 18572 13584
rect 18538 13482 18572 13516
rect 18538 13414 18572 13448
rect 18538 13346 18572 13380
rect 18538 13278 18572 13312
rect 18538 13210 18572 13244
rect 18538 13142 18572 13176
rect 18538 13074 18572 13108
rect 18538 13006 18572 13040
rect 18538 12938 18572 12972
rect 18538 12870 18572 12904
rect 18538 12802 18572 12836
rect 18538 12734 18572 12768
rect 18538 12666 18572 12700
rect 18538 12598 18572 12632
rect 18538 12530 18572 12564
rect 18538 12462 18572 12496
rect 18538 12394 18572 12428
rect 18538 12326 18572 12360
rect 18538 12258 18572 12292
rect 18538 12190 18572 12224
rect 18538 12122 18572 12156
rect 18538 12054 18572 12088
rect 18538 11986 18572 12020
rect 18538 11918 18572 11952
rect 18538 11850 18572 11884
rect 18538 11782 18572 11816
rect 19596 14706 19630 14740
rect 19596 14638 19630 14672
rect 19596 14570 19630 14604
rect 19596 14502 19630 14536
rect 19596 14434 19630 14468
rect 19596 14366 19630 14400
rect 19596 14298 19630 14332
rect 19596 14230 19630 14264
rect 19596 14162 19630 14196
rect 19596 14094 19630 14128
rect 19596 14026 19630 14060
rect 19596 13958 19630 13992
rect 19596 13890 19630 13924
rect 19596 13822 19630 13856
rect 19596 13754 19630 13788
rect 19596 13686 19630 13720
rect 19596 13618 19630 13652
rect 19596 13550 19630 13584
rect 19596 13482 19630 13516
rect 19596 13414 19630 13448
rect 19596 13346 19630 13380
rect 19596 13278 19630 13312
rect 19596 13210 19630 13244
rect 19596 13142 19630 13176
rect 19596 13074 19630 13108
rect 19596 13006 19630 13040
rect 19596 12938 19630 12972
rect 19596 12870 19630 12904
rect 19596 12802 19630 12836
rect 19596 12734 19630 12768
rect 19596 12666 19630 12700
rect 19596 12598 19630 12632
rect 19596 12530 19630 12564
rect 19596 12462 19630 12496
rect 19596 12394 19630 12428
rect 19596 12326 19630 12360
rect 19596 12258 19630 12292
rect 19596 12190 19630 12224
rect 19596 12122 19630 12156
rect 19596 12054 19630 12088
rect 19596 11986 19630 12020
rect 19596 11918 19630 11952
rect 19596 11850 19630 11884
rect 19596 11782 19630 11816
rect 14954 11192 14988 11226
rect 14954 11124 14988 11158
rect 14954 11056 14988 11090
rect 14954 10988 14988 11022
rect 14954 10920 14988 10954
rect 14954 10852 14988 10886
rect 14954 10784 14988 10818
rect 14954 10716 14988 10750
rect 14954 10648 14988 10682
rect 14954 10580 14988 10614
rect 14954 10512 14988 10546
rect 14954 10444 14988 10478
rect 14954 10376 14988 10410
rect 14954 10308 14988 10342
rect 14954 10240 14988 10274
rect 14954 10172 14988 10206
rect 14954 10104 14988 10138
rect 14954 10036 14988 10070
rect 14954 9968 14988 10002
rect 14954 9900 14988 9934
rect 14954 9832 14988 9866
rect 14954 9764 14988 9798
rect 14954 9696 14988 9730
rect 14954 9628 14988 9662
rect 14954 9560 14988 9594
rect 14954 9492 14988 9526
rect 14954 9424 14988 9458
rect 14954 9356 14988 9390
rect 14954 9288 14988 9322
rect 14954 9220 14988 9254
rect 14954 9152 14988 9186
rect 14954 9084 14988 9118
rect 14954 9016 14988 9050
rect 14954 8948 14988 8982
rect 14954 8880 14988 8914
rect 14954 8812 14988 8846
rect 14954 8744 14988 8778
rect 14954 8676 14988 8710
rect 14954 8608 14988 8642
rect 14954 8540 14988 8574
rect 14954 8472 14988 8506
rect 14954 8404 14988 8438
rect 14954 8336 14988 8370
rect 14954 8268 14988 8302
rect 16012 11192 16046 11226
rect 16012 11124 16046 11158
rect 16012 11056 16046 11090
rect 16012 10988 16046 11022
rect 16012 10920 16046 10954
rect 16012 10852 16046 10886
rect 16012 10784 16046 10818
rect 16012 10716 16046 10750
rect 16012 10648 16046 10682
rect 16012 10580 16046 10614
rect 16012 10512 16046 10546
rect 16012 10444 16046 10478
rect 16012 10376 16046 10410
rect 16012 10308 16046 10342
rect 16012 10240 16046 10274
rect 16012 10172 16046 10206
rect 16012 10104 16046 10138
rect 16012 10036 16046 10070
rect 16012 9968 16046 10002
rect 16012 9900 16046 9934
rect 16012 9832 16046 9866
rect 16012 9764 16046 9798
rect 16012 9696 16046 9730
rect 16012 9628 16046 9662
rect 16012 9560 16046 9594
rect 16012 9492 16046 9526
rect 16012 9424 16046 9458
rect 16012 9356 16046 9390
rect 16012 9288 16046 9322
rect 16012 9220 16046 9254
rect 16012 9152 16046 9186
rect 16012 9084 16046 9118
rect 16012 9016 16046 9050
rect 16012 8948 16046 8982
rect 16012 8880 16046 8914
rect 16012 8812 16046 8846
rect 16012 8744 16046 8778
rect 16012 8676 16046 8710
rect 16012 8608 16046 8642
rect 16012 8540 16046 8574
rect 16012 8472 16046 8506
rect 16012 8404 16046 8438
rect 16012 8336 16046 8370
rect 16012 8268 16046 8302
rect 17070 11192 17104 11226
rect 17070 11124 17104 11158
rect 17070 11056 17104 11090
rect 17070 10988 17104 11022
rect 17070 10920 17104 10954
rect 17070 10852 17104 10886
rect 17070 10784 17104 10818
rect 17070 10716 17104 10750
rect 17070 10648 17104 10682
rect 17070 10580 17104 10614
rect 17070 10512 17104 10546
rect 17070 10444 17104 10478
rect 17070 10376 17104 10410
rect 17070 10308 17104 10342
rect 17070 10240 17104 10274
rect 17070 10172 17104 10206
rect 17070 10104 17104 10138
rect 17070 10036 17104 10070
rect 17070 9968 17104 10002
rect 17070 9900 17104 9934
rect 17070 9832 17104 9866
rect 17070 9764 17104 9798
rect 17070 9696 17104 9730
rect 17070 9628 17104 9662
rect 17070 9560 17104 9594
rect 17070 9492 17104 9526
rect 17070 9424 17104 9458
rect 17070 9356 17104 9390
rect 17070 9288 17104 9322
rect 17070 9220 17104 9254
rect 17070 9152 17104 9186
rect 17070 9084 17104 9118
rect 17070 9016 17104 9050
rect 17070 8948 17104 8982
rect 17070 8880 17104 8914
rect 17070 8812 17104 8846
rect 17070 8744 17104 8778
rect 17070 8676 17104 8710
rect 17070 8608 17104 8642
rect 17070 8540 17104 8574
rect 17070 8472 17104 8506
rect 17070 8404 17104 8438
rect 17070 8336 17104 8370
rect 17070 8268 17104 8302
rect 17478 11166 17512 11200
rect 17478 11098 17512 11132
rect 17478 11030 17512 11064
rect 17478 10962 17512 10996
rect 17478 10894 17512 10928
rect 17478 10826 17512 10860
rect 17478 10758 17512 10792
rect 17478 10690 17512 10724
rect 17478 10622 17512 10656
rect 17478 10554 17512 10588
rect 17478 10486 17512 10520
rect 17478 10418 17512 10452
rect 17478 10350 17512 10384
rect 17478 10282 17512 10316
rect 17478 10214 17512 10248
rect 17478 10146 17512 10180
rect 17478 10078 17512 10112
rect 17478 10010 17512 10044
rect 17478 9942 17512 9976
rect 17478 9874 17512 9908
rect 17478 9806 17512 9840
rect 17478 9738 17512 9772
rect 17478 9670 17512 9704
rect 17478 9602 17512 9636
rect 17478 9534 17512 9568
rect 17478 9466 17512 9500
rect 17478 9398 17512 9432
rect 17478 9330 17512 9364
rect 17478 9262 17512 9296
rect 17478 9194 17512 9228
rect 17478 9126 17512 9160
rect 17478 9058 17512 9092
rect 17478 8990 17512 9024
rect 17478 8922 17512 8956
rect 17478 8854 17512 8888
rect 17478 8786 17512 8820
rect 17478 8718 17512 8752
rect 17478 8650 17512 8684
rect 17478 8582 17512 8616
rect 17478 8514 17512 8548
rect 17478 8446 17512 8480
rect 17478 8378 17512 8412
rect 17478 8310 17512 8344
rect 17478 8242 17512 8276
rect 18536 11166 18570 11200
rect 18536 11098 18570 11132
rect 18536 11030 18570 11064
rect 18536 10962 18570 10996
rect 18536 10894 18570 10928
rect 18536 10826 18570 10860
rect 18536 10758 18570 10792
rect 18536 10690 18570 10724
rect 18536 10622 18570 10656
rect 18536 10554 18570 10588
rect 18536 10486 18570 10520
rect 18536 10418 18570 10452
rect 18536 10350 18570 10384
rect 18536 10282 18570 10316
rect 18536 10214 18570 10248
rect 18536 10146 18570 10180
rect 18536 10078 18570 10112
rect 18536 10010 18570 10044
rect 18536 9942 18570 9976
rect 18536 9874 18570 9908
rect 18536 9806 18570 9840
rect 18536 9738 18570 9772
rect 18536 9670 18570 9704
rect 18536 9602 18570 9636
rect 18536 9534 18570 9568
rect 18536 9466 18570 9500
rect 18536 9398 18570 9432
rect 18536 9330 18570 9364
rect 18536 9262 18570 9296
rect 18536 9194 18570 9228
rect 18536 9126 18570 9160
rect 18536 9058 18570 9092
rect 18536 8990 18570 9024
rect 18536 8922 18570 8956
rect 18536 8854 18570 8888
rect 18536 8786 18570 8820
rect 18536 8718 18570 8752
rect 18536 8650 18570 8684
rect 18536 8582 18570 8616
rect 18536 8514 18570 8548
rect 18536 8446 18570 8480
rect 18536 8378 18570 8412
rect 18536 8310 18570 8344
rect 18536 8242 18570 8276
rect 19594 11166 19628 11200
rect 19594 11098 19628 11132
rect 19594 11030 19628 11064
rect 19594 10962 19628 10996
rect 19594 10894 19628 10928
rect 19594 10826 19628 10860
rect 19594 10758 19628 10792
rect 19594 10690 19628 10724
rect 19594 10622 19628 10656
rect 19594 10554 19628 10588
rect 19594 10486 19628 10520
rect 19594 10418 19628 10452
rect 19594 10350 19628 10384
rect 19594 10282 19628 10316
rect 19594 10214 19628 10248
rect 19594 10146 19628 10180
rect 19594 10078 19628 10112
rect 19594 10010 19628 10044
rect 19594 9942 19628 9976
rect 19594 9874 19628 9908
rect 19594 9806 19628 9840
rect 19594 9738 19628 9772
rect 19594 9670 19628 9704
rect 19594 9602 19628 9636
rect 19594 9534 19628 9568
rect 19594 9466 19628 9500
rect 19594 9398 19628 9432
rect 19594 9330 19628 9364
rect 19594 9262 19628 9296
rect 19594 9194 19628 9228
rect 19594 9126 19628 9160
rect 19594 9058 19628 9092
rect 19594 8990 19628 9024
rect 19594 8922 19628 8956
rect 19594 8854 19628 8888
rect 19594 8786 19628 8820
rect 19594 8718 19628 8752
rect 19594 8650 19628 8684
rect 19594 8582 19628 8616
rect 19594 8514 19628 8548
rect 19594 8446 19628 8480
rect 19594 8378 19628 8412
rect 19594 8310 19628 8344
rect 19594 8242 19628 8276
rect 23250 13322 23284 13356
rect 23318 13322 23352 13356
rect 23386 13322 23420 13356
rect 23454 13322 23488 13356
rect 23522 13322 23556 13356
rect 23590 13322 23624 13356
rect 23658 13322 23692 13356
rect 23726 13322 23760 13356
rect 23794 13322 23828 13356
rect 23862 13322 23896 13356
rect 23930 13322 23964 13356
rect 23998 13322 24032 13356
rect 24066 13322 24100 13356
rect 24134 13322 24168 13356
rect 23250 12264 23284 12298
rect 23318 12264 23352 12298
rect 23386 12264 23420 12298
rect 23454 12264 23488 12298
rect 23522 12264 23556 12298
rect 23590 12264 23624 12298
rect 23658 12264 23692 12298
rect 23726 12264 23760 12298
rect 23794 12264 23828 12298
rect 23862 12264 23896 12298
rect 23930 12264 23964 12298
rect 23998 12264 24032 12298
rect 24066 12264 24100 12298
rect 24134 12264 24168 12298
rect 24810 13316 24844 13350
rect 24878 13316 24912 13350
rect 24946 13316 24980 13350
rect 25014 13316 25048 13350
rect 25082 13316 25116 13350
rect 25150 13316 25184 13350
rect 25218 13316 25252 13350
rect 25286 13316 25320 13350
rect 25354 13316 25388 13350
rect 25422 13316 25456 13350
rect 25490 13316 25524 13350
rect 25558 13316 25592 13350
rect 25626 13316 25660 13350
rect 25694 13316 25728 13350
rect 24810 12258 24844 12292
rect 24878 12258 24912 12292
rect 24946 12258 24980 12292
rect 25014 12258 25048 12292
rect 25082 12258 25116 12292
rect 25150 12258 25184 12292
rect 25218 12258 25252 12292
rect 25286 12258 25320 12292
rect 25354 12258 25388 12292
rect 25422 12258 25456 12292
rect 25490 12258 25524 12292
rect 25558 12258 25592 12292
rect 25626 12258 25660 12292
rect 25694 12258 25728 12292
rect 24810 11200 24844 11234
rect 24878 11200 24912 11234
rect 24946 11200 24980 11234
rect 25014 11200 25048 11234
rect 25082 11200 25116 11234
rect 25150 11200 25184 11234
rect 25218 11200 25252 11234
rect 25286 11200 25320 11234
rect 25354 11200 25388 11234
rect 25422 11200 25456 11234
rect 25490 11200 25524 11234
rect 25558 11200 25592 11234
rect 25626 11200 25660 11234
rect 25694 11200 25728 11234
rect 24810 10142 24844 10176
rect 24878 10142 24912 10176
rect 24946 10142 24980 10176
rect 25014 10142 25048 10176
rect 25082 10142 25116 10176
rect 25150 10142 25184 10176
rect 25218 10142 25252 10176
rect 25286 10142 25320 10176
rect 25354 10142 25388 10176
rect 25422 10142 25456 10176
rect 25490 10142 25524 10176
rect 25558 10142 25592 10176
rect 25626 10142 25660 10176
rect 25694 10142 25728 10176
rect 24810 9084 24844 9118
rect 24878 9084 24912 9118
rect 24946 9084 24980 9118
rect 25014 9084 25048 9118
rect 25082 9084 25116 9118
rect 25150 9084 25184 9118
rect 25218 9084 25252 9118
rect 25286 9084 25320 9118
rect 25354 9084 25388 9118
rect 25422 9084 25456 9118
rect 25490 9084 25524 9118
rect 25558 9084 25592 9118
rect 25626 9084 25660 9118
rect 25694 9084 25728 9118
<< psubdiff >>
rect 24460 16716 24559 16750
rect 24593 16716 24627 16750
rect 24661 16716 24695 16750
rect 24729 16716 24763 16750
rect 24797 16716 24831 16750
rect 24865 16716 24899 16750
rect 24933 16716 24967 16750
rect 25001 16716 25035 16750
rect 25069 16716 25103 16750
rect 25137 16716 25171 16750
rect 25205 16716 25239 16750
rect 25273 16716 25307 16750
rect 25341 16716 25375 16750
rect 25409 16716 25443 16750
rect 25477 16716 25511 16750
rect 25545 16716 25579 16750
rect 25613 16716 25647 16750
rect 25681 16716 25715 16750
rect 25749 16716 25783 16750
rect 25817 16716 25851 16750
rect 25885 16716 25919 16750
rect 25953 16716 25987 16750
rect 26021 16716 26055 16750
rect 26089 16716 26123 16750
rect 26157 16716 26191 16750
rect 26225 16716 26259 16750
rect 26293 16716 26327 16750
rect 26361 16716 26395 16750
rect 26429 16716 26463 16750
rect 26497 16716 26531 16750
rect 26565 16716 26599 16750
rect 26633 16716 26667 16750
rect 26701 16716 26735 16750
rect 26769 16716 26803 16750
rect 26837 16716 26871 16750
rect 26905 16716 26939 16750
rect 26973 16716 27007 16750
rect 27041 16716 27075 16750
rect 27109 16716 27143 16750
rect 27177 16716 27211 16750
rect 27245 16716 27279 16750
rect 27313 16716 27347 16750
rect 27381 16716 27415 16750
rect 27449 16716 27483 16750
rect 27517 16716 27551 16750
rect 27585 16716 27684 16750
rect 24460 16646 24494 16716
rect 27650 16646 27684 16716
rect 24460 16578 24494 16612
rect 27650 16578 27684 16612
rect 24460 16510 24494 16544
rect 24460 16442 24494 16476
rect 24460 16374 24494 16408
rect 24460 16306 24494 16340
rect 27650 16510 27684 16544
rect 27650 16442 27684 16476
rect 27650 16374 27684 16408
rect 27650 16306 27684 16340
rect 24460 16238 24494 16272
rect 27650 16238 27684 16272
rect 24460 16170 24494 16204
rect 24460 16102 24494 16136
rect 24460 16034 24494 16068
rect 24460 15966 24494 16000
rect 27650 16170 27684 16204
rect 27650 16102 27684 16136
rect 27650 16034 27684 16068
rect 24460 15898 24494 15932
rect 27650 15966 27684 16000
rect 23110 15817 24398 15852
rect 23110 15794 23240 15817
rect 23110 15760 23144 15794
rect 23178 15783 23240 15794
rect 23274 15783 23330 15817
rect 23364 15783 23420 15817
rect 23454 15783 23510 15817
rect 23544 15783 23600 15817
rect 23634 15783 23690 15817
rect 23724 15783 23780 15817
rect 23814 15783 23870 15817
rect 23904 15783 23960 15817
rect 23994 15783 24050 15817
rect 24084 15783 24140 15817
rect 24174 15783 24230 15817
rect 24264 15794 24398 15817
rect 24264 15783 24331 15794
rect 23178 15760 24331 15783
rect 24365 15760 24398 15794
rect 23110 15751 24398 15760
rect 23110 15704 23211 15751
rect 23110 15670 23144 15704
rect 23178 15670 23211 15704
rect 24297 15704 24398 15751
rect 23110 15614 23211 15670
rect 23110 15580 23144 15614
rect 23178 15580 23211 15614
rect 23110 15524 23211 15580
rect -7886 15466 -4427 15515
rect -7886 15432 -7630 15466
rect -7596 15432 -7562 15466
rect -7528 15432 -7494 15466
rect -7460 15432 -7426 15466
rect -7392 15432 -7358 15466
rect -7324 15432 -7290 15466
rect -7256 15432 -7222 15466
rect -7188 15432 -7154 15466
rect -7120 15432 -7086 15466
rect -7052 15432 -7018 15466
rect -6984 15432 -6950 15466
rect -6916 15432 -6882 15466
rect -6848 15432 -6814 15466
rect -6780 15432 -6746 15466
rect -6712 15432 -6678 15466
rect -6644 15432 -6610 15466
rect -6576 15432 -6542 15466
rect -6508 15432 -6474 15466
rect -6440 15432 -6406 15466
rect -6372 15432 -6338 15466
rect -6304 15432 -6270 15466
rect -6236 15432 -6202 15466
rect -6168 15432 -6134 15466
rect -6100 15432 -6066 15466
rect -6032 15432 -5998 15466
rect -5964 15432 -5930 15466
rect -5896 15432 -5862 15466
rect -5828 15432 -5794 15466
rect -5760 15432 -5726 15466
rect -5692 15432 -5658 15466
rect -5624 15432 -5590 15466
rect -5556 15432 -5522 15466
rect -5488 15432 -5454 15466
rect -5420 15432 -5386 15466
rect -5352 15432 -5318 15466
rect -5284 15432 -5250 15466
rect -5216 15432 -5182 15466
rect -5148 15432 -5114 15466
rect -5080 15432 -5046 15466
rect -5012 15432 -4978 15466
rect -4944 15432 -4910 15466
rect -4876 15432 -4842 15466
rect -4808 15432 -4774 15466
rect -4740 15432 -4706 15466
rect -4672 15432 -4427 15466
rect -7886 15381 -4427 15432
rect -7886 15308 -7753 15381
rect -7886 15274 -7843 15308
rect -7809 15274 -7753 15308
rect -7886 15240 -7753 15274
rect -7886 15206 -7843 15240
rect -7809 15206 -7753 15240
rect -7886 15172 -7753 15206
rect -7886 15138 -7843 15172
rect -7809 15138 -7753 15172
rect -7886 15104 -7753 15138
rect -7886 15070 -7843 15104
rect -7809 15070 -7753 15104
rect -7886 15036 -7753 15070
rect -7886 15002 -7843 15036
rect -7809 15002 -7753 15036
rect -7886 14968 -7753 15002
rect -4545 15268 -4427 15381
rect -4545 15234 -4503 15268
rect -4469 15234 -4427 15268
rect -4545 15200 -4427 15234
rect -4545 15166 -4503 15200
rect -4469 15166 -4427 15200
rect -4545 15132 -4427 15166
rect -4545 15098 -4503 15132
rect -4469 15098 -4427 15132
rect -4545 15064 -4427 15098
rect -4545 15030 -4503 15064
rect -4469 15030 -4427 15064
rect 23110 15490 23144 15524
rect 23178 15490 23211 15524
rect 23110 15434 23211 15490
rect 23110 15400 23144 15434
rect 23178 15400 23211 15434
rect 23110 15344 23211 15400
rect 23110 15310 23144 15344
rect 23178 15310 23211 15344
rect 23110 15254 23211 15310
rect 23110 15220 23144 15254
rect 23178 15220 23211 15254
rect 23110 15164 23211 15220
rect 23110 15130 23144 15164
rect 23178 15130 23211 15164
rect 23110 15074 23211 15130
rect 23110 15040 23144 15074
rect 23178 15040 23211 15074
rect -7886 14934 -7843 14968
rect -7809 14934 -7753 14968
rect -7886 14900 -7753 14934
rect -7886 14866 -7843 14900
rect -7809 14866 -7753 14900
rect -7886 14832 -7753 14866
rect -4545 14996 -4427 15030
rect -4545 14962 -4503 14996
rect -4469 14962 -4427 14996
rect -4545 14928 -4427 14962
rect -4545 14894 -4503 14928
rect -4469 14894 -4427 14928
rect -4545 14860 -4427 14894
rect -7886 14798 -7843 14832
rect -7809 14798 -7753 14832
rect -7886 14764 -7753 14798
rect -7886 14730 -7843 14764
rect -7809 14730 -7753 14764
rect -7886 14696 -7753 14730
rect -7886 14662 -7843 14696
rect -7809 14662 -7753 14696
rect -7886 14628 -7753 14662
rect -7886 14594 -7843 14628
rect -7809 14594 -7753 14628
rect -7886 14560 -7753 14594
rect -7886 14526 -7843 14560
rect -7809 14526 -7753 14560
rect -7886 14492 -7753 14526
rect -7886 14458 -7843 14492
rect -7809 14458 -7753 14492
rect -7886 14424 -7753 14458
rect -7886 14390 -7843 14424
rect -7809 14390 -7753 14424
rect -7886 14356 -7753 14390
rect -7886 14322 -7843 14356
rect -7809 14322 -7753 14356
rect -7886 14288 -7753 14322
rect -7886 14254 -7843 14288
rect -7809 14254 -7753 14288
rect -7886 14220 -7753 14254
rect -7886 14186 -7843 14220
rect -7809 14186 -7753 14220
rect -7886 14152 -7753 14186
rect -7886 14118 -7843 14152
rect -7809 14118 -7753 14152
rect -7886 14084 -7753 14118
rect -7886 14050 -7843 14084
rect -7809 14050 -7753 14084
rect -7886 14016 -7753 14050
rect -7886 13982 -7843 14016
rect -7809 13982 -7753 14016
rect -7886 13948 -7753 13982
rect -7886 13914 -7843 13948
rect -7809 13914 -7753 13948
rect -7886 13880 -7753 13914
rect -7886 13846 -7843 13880
rect -7809 13846 -7753 13880
rect -7886 13812 -7753 13846
rect -7886 13778 -7843 13812
rect -7809 13778 -7753 13812
rect -7886 13744 -7753 13778
rect -7886 13710 -7843 13744
rect -7809 13710 -7753 13744
rect -7886 13676 -7753 13710
rect -7886 13642 -7843 13676
rect -7809 13642 -7753 13676
rect -7886 13608 -7753 13642
rect -7886 13574 -7843 13608
rect -7809 13574 -7753 13608
rect -7886 13540 -7753 13574
rect -7886 13506 -7843 13540
rect -7809 13506 -7753 13540
rect -7886 13472 -7753 13506
rect -7886 13438 -7843 13472
rect -7809 13438 -7753 13472
rect -7886 13404 -7753 13438
rect -7886 13370 -7843 13404
rect -7809 13370 -7753 13404
rect -7886 13336 -7753 13370
rect -7886 13302 -7843 13336
rect -7809 13302 -7753 13336
rect -7886 13268 -7753 13302
rect -7886 13234 -7843 13268
rect -7809 13234 -7753 13268
rect -7886 13200 -7753 13234
rect -7886 13166 -7843 13200
rect -7809 13166 -7753 13200
rect -7886 13132 -7753 13166
rect -7886 13098 -7843 13132
rect -7809 13098 -7753 13132
rect -7886 13064 -7753 13098
rect -7886 13030 -7843 13064
rect -7809 13030 -7753 13064
rect -7886 12996 -7753 13030
rect -7886 12962 -7843 12996
rect -7809 12962 -7753 12996
rect -7886 12928 -7753 12962
rect -7886 12894 -7843 12928
rect -7809 12894 -7753 12928
rect -7886 12860 -7753 12894
rect -7886 12826 -7843 12860
rect -7809 12826 -7753 12860
rect -4545 14826 -4503 14860
rect -4469 14826 -4427 14860
rect -4545 14792 -4427 14826
rect -4545 14758 -4503 14792
rect -4469 14758 -4427 14792
rect -4545 14724 -4427 14758
rect -4545 14690 -4503 14724
rect -4469 14690 -4427 14724
rect -4545 14656 -4427 14690
rect -4545 14622 -4503 14656
rect -4469 14622 -4427 14656
rect -4545 14588 -4427 14622
rect -4545 14554 -4503 14588
rect -4469 14554 -4427 14588
rect -4545 14520 -4427 14554
rect -4545 14486 -4503 14520
rect -4469 14486 -4427 14520
rect -4545 14452 -4427 14486
rect -4545 14418 -4503 14452
rect -4469 14418 -4427 14452
rect -4545 14384 -4427 14418
rect -4545 14350 -4503 14384
rect -4469 14350 -4427 14384
rect -4545 14316 -4427 14350
rect -4545 14282 -4503 14316
rect -4469 14282 -4427 14316
rect -4545 14248 -4427 14282
rect -4545 14214 -4503 14248
rect -4469 14214 -4427 14248
rect -4545 14180 -4427 14214
rect -4545 14146 -4503 14180
rect -4469 14146 -4427 14180
rect -4545 14112 -4427 14146
rect -4545 14078 -4503 14112
rect -4469 14078 -4427 14112
rect -4545 14044 -4427 14078
rect -4545 14010 -4503 14044
rect -4469 14010 -4427 14044
rect -4545 13976 -4427 14010
rect -4545 13942 -4503 13976
rect -4469 13942 -4427 13976
rect -4545 13908 -4427 13942
rect -4545 13874 -4503 13908
rect -4469 13874 -4427 13908
rect -4545 13840 -4427 13874
rect -4545 13806 -4503 13840
rect -4469 13806 -4427 13840
rect -4545 13772 -4427 13806
rect -4545 13738 -4503 13772
rect -4469 13738 -4427 13772
rect -4545 13704 -4427 13738
rect -4545 13670 -4503 13704
rect -4469 13670 -4427 13704
rect -4545 13636 -4427 13670
rect -4545 13602 -4503 13636
rect -4469 13602 -4427 13636
rect -4545 13568 -4427 13602
rect -4545 13534 -4503 13568
rect -4469 13534 -4427 13568
rect -4545 13500 -4427 13534
rect -4545 13466 -4503 13500
rect -4469 13466 -4427 13500
rect -4545 13432 -4427 13466
rect -4545 13398 -4503 13432
rect -4469 13398 -4427 13432
rect -4545 13364 -4427 13398
rect -4545 13330 -4503 13364
rect -4469 13330 -4427 13364
rect -4545 13296 -4427 13330
rect -4545 13262 -4503 13296
rect -4469 13262 -4427 13296
rect -4545 13228 -4427 13262
rect -4545 13194 -4503 13228
rect -4469 13194 -4427 13228
rect -4545 13160 -4427 13194
rect -4545 13126 -4503 13160
rect -4469 13126 -4427 13160
rect -4545 13092 -4427 13126
rect -4545 13058 -4503 13092
rect -4469 13058 -4427 13092
rect -4545 13024 -4427 13058
rect -4545 12990 -4503 13024
rect -4469 12990 -4427 13024
rect -4545 12956 -4427 12990
rect -4545 12922 -4503 12956
rect -4469 12922 -4427 12956
rect -4545 12888 -4427 12922
rect -4545 12854 -4503 12888
rect -4469 12854 -4427 12888
rect -7886 12792 -7753 12826
rect -4545 12820 -4427 12854
rect -7886 12758 -7843 12792
rect -7809 12758 -7753 12792
rect -7886 12724 -7753 12758
rect -7886 12690 -7843 12724
rect -7809 12690 -7753 12724
rect -7886 12656 -7753 12690
rect -7886 12622 -7843 12656
rect -7809 12622 -7753 12656
rect -4545 12786 -4503 12820
rect -4469 12786 -4427 12820
rect -4545 12752 -4427 12786
rect -4545 12718 -4503 12752
rect -4469 12718 -4427 12752
rect -4545 12684 -4427 12718
rect -4545 12650 -4503 12684
rect -4469 12650 -4427 12684
rect -7886 12588 -7753 12622
rect -7886 12554 -7843 12588
rect -7809 12554 -7753 12588
rect -7886 12520 -7753 12554
rect -7886 12486 -7843 12520
rect -7809 12486 -7753 12520
rect -7886 12452 -7753 12486
rect -7886 12418 -7843 12452
rect -7809 12418 -7753 12452
rect -7886 12384 -7753 12418
rect -7886 12350 -7843 12384
rect -7809 12350 -7753 12384
rect -7886 12276 -7753 12350
rect -4545 12616 -4427 12650
rect -4545 12582 -4503 12616
rect -4469 12582 -4427 12616
rect -4545 12548 -4427 12582
rect -4545 12514 -4503 12548
rect -4469 12514 -4427 12548
rect -4545 12480 -4427 12514
rect -4545 12446 -4503 12480
rect -4469 12446 -4427 12480
rect -4545 12412 -4427 12446
rect -4545 12378 -4503 12412
rect -4469 12378 -4427 12412
rect -4545 12344 -4427 12378
rect -4545 12310 -4503 12344
rect -4469 12310 -4427 12344
rect -4010 15001 -3896 15035
rect -3862 15001 -3828 15035
rect -3794 15001 -3680 15035
rect -4010 14914 -3976 15001
rect -3714 14914 -3680 15001
rect -4010 14846 -3976 14880
rect -4010 14778 -3976 14812
rect -4010 14710 -3976 14744
rect -4010 14642 -3976 14676
rect -4010 14574 -3976 14608
rect -4010 14506 -3976 14540
rect -4010 14438 -3976 14472
rect -4010 14370 -3976 14404
rect -4010 14302 -3976 14336
rect -4010 14234 -3976 14268
rect -4010 14166 -3976 14200
rect -4010 14098 -3976 14132
rect -4010 14030 -3976 14064
rect -4010 13962 -3976 13996
rect -4010 13894 -3976 13928
rect -4010 13826 -3976 13860
rect -4010 13758 -3976 13792
rect -4010 13690 -3976 13724
rect -4010 13622 -3976 13656
rect -4010 13554 -3976 13588
rect -4010 13486 -3976 13520
rect -4010 13418 -3976 13452
rect -4010 13350 -3976 13384
rect -4010 13282 -3976 13316
rect -4010 13214 -3976 13248
rect -4010 13146 -3976 13180
rect -4010 13078 -3976 13112
rect -4010 13010 -3976 13044
rect -4010 12942 -3976 12976
rect -4010 12874 -3976 12908
rect -4010 12806 -3976 12840
rect -4010 12738 -3976 12772
rect -4010 12670 -3976 12704
rect -4010 12602 -3976 12636
rect -4010 12534 -3976 12568
rect -4010 12466 -3976 12500
rect -3714 14846 -3680 14880
rect -3714 14778 -3680 14812
rect -3714 14710 -3680 14744
rect -3714 14642 -3680 14676
rect -3714 14574 -3680 14608
rect -3714 14506 -3680 14540
rect -3714 14438 -3680 14472
rect -3714 14370 -3680 14404
rect -3714 14302 -3680 14336
rect -3714 14234 -3680 14268
rect -3714 14166 -3680 14200
rect -3714 14098 -3680 14132
rect -3714 14030 -3680 14064
rect -3714 13962 -3680 13996
rect -3714 13894 -3680 13928
rect -3714 13826 -3680 13860
rect -3714 13758 -3680 13792
rect -3714 13690 -3680 13724
rect -3714 13622 -3680 13656
rect -3714 13554 -3680 13588
rect -3714 13486 -3680 13520
rect -3714 13418 -3680 13452
rect -3714 13350 -3680 13384
rect -3714 13282 -3680 13316
rect -3714 13214 -3680 13248
rect -3714 13146 -3680 13180
rect -3714 13078 -3680 13112
rect -3714 13010 -3680 13044
rect -3714 12942 -3680 12976
rect -3714 12874 -3680 12908
rect -3714 12806 -3680 12840
rect -3714 12738 -3680 12772
rect -3714 12670 -3680 12704
rect -3714 12602 -3680 12636
rect -3714 12534 -3680 12568
rect -3714 12466 -3680 12500
rect -4010 12345 -3976 12432
rect -3714 12345 -3680 12432
rect -4010 12311 -3896 12345
rect -3862 12311 -3828 12345
rect -3794 12311 -3680 12345
rect -4545 12276 -4427 12310
rect -7886 12236 -4427 12276
rect -7886 12202 -7570 12236
rect -7536 12202 -7502 12236
rect -7468 12202 -7434 12236
rect -7400 12202 -7366 12236
rect -7332 12202 -7298 12236
rect -7264 12202 -7230 12236
rect -7196 12202 -7162 12236
rect -7128 12202 -7094 12236
rect -7060 12202 -7026 12236
rect -6992 12202 -6958 12236
rect -6924 12202 -6890 12236
rect -6856 12202 -6822 12236
rect -6788 12202 -6754 12236
rect -6720 12202 -6686 12236
rect -6652 12202 -6618 12236
rect -6584 12202 -6550 12236
rect -6516 12202 -6482 12236
rect -6448 12202 -6414 12236
rect -6380 12202 -6346 12236
rect -6312 12202 -6278 12236
rect -6244 12202 -6210 12236
rect -6176 12202 -6142 12236
rect -6108 12202 -6074 12236
rect -6040 12202 -6006 12236
rect -5972 12202 -5938 12236
rect -5904 12202 -5870 12236
rect -5836 12202 -5802 12236
rect -5768 12202 -5734 12236
rect -5700 12202 -5666 12236
rect -5632 12202 -5598 12236
rect -5564 12202 -5530 12236
rect -5496 12202 -5462 12236
rect -5428 12202 -5394 12236
rect -5360 12202 -5326 12236
rect -5292 12202 -5258 12236
rect -5224 12202 -5190 12236
rect -5156 12202 -5122 12236
rect -5088 12202 -5054 12236
rect -5020 12202 -4986 12236
rect -4952 12202 -4918 12236
rect -4884 12202 -4850 12236
rect -4816 12202 -4782 12236
rect -4748 12202 -4714 12236
rect -4680 12202 -4646 12236
rect -4612 12202 -4427 12236
rect -7886 12134 -4427 12202
rect 23110 14984 23211 15040
rect 23110 14950 23144 14984
rect 23178 14950 23211 14984
rect 23110 14894 23211 14950
rect 23110 14860 23144 14894
rect 23178 14860 23211 14894
rect 23110 14804 23211 14860
rect 23110 14770 23144 14804
rect 23178 14770 23211 14804
rect 23110 14714 23211 14770
rect 24297 15670 24331 15704
rect 24365 15670 24398 15704
rect 24297 15614 24398 15670
rect 24297 15580 24331 15614
rect 24365 15580 24398 15614
rect 24297 15524 24398 15580
rect 24297 15490 24331 15524
rect 24365 15490 24398 15524
rect 24297 15434 24398 15490
rect 24297 15400 24331 15434
rect 24365 15400 24398 15434
rect 24297 15344 24398 15400
rect 24297 15310 24331 15344
rect 24365 15310 24398 15344
rect 24297 15254 24398 15310
rect 24297 15220 24331 15254
rect 24365 15220 24398 15254
rect 24297 15164 24398 15220
rect 24297 15130 24331 15164
rect 24365 15130 24398 15164
rect 24460 15830 24494 15864
rect 24460 15762 24494 15796
rect 24460 15694 24494 15728
rect 27650 15898 27684 15932
rect 27650 15830 27684 15864
rect 27650 15762 27684 15796
rect 27650 15694 27684 15728
rect 24460 15626 24494 15660
rect 27650 15626 27684 15660
rect 24460 15558 24494 15592
rect 24460 15490 24494 15524
rect 24460 15422 24494 15456
rect 24460 15354 24494 15388
rect 27650 15558 27684 15592
rect 27650 15490 27684 15524
rect 27650 15422 27684 15456
rect 37706 16216 41165 16265
rect 37706 16182 37962 16216
rect 37996 16182 38030 16216
rect 38064 16182 38098 16216
rect 38132 16182 38166 16216
rect 38200 16182 38234 16216
rect 38268 16182 38302 16216
rect 38336 16182 38370 16216
rect 38404 16182 38438 16216
rect 38472 16182 38506 16216
rect 38540 16182 38574 16216
rect 38608 16182 38642 16216
rect 38676 16182 38710 16216
rect 38744 16182 38778 16216
rect 38812 16182 38846 16216
rect 38880 16182 38914 16216
rect 38948 16182 38982 16216
rect 39016 16182 39050 16216
rect 39084 16182 39118 16216
rect 39152 16182 39186 16216
rect 39220 16182 39254 16216
rect 39288 16182 39322 16216
rect 39356 16182 39390 16216
rect 39424 16182 39458 16216
rect 39492 16182 39526 16216
rect 39560 16182 39594 16216
rect 39628 16182 39662 16216
rect 39696 16182 39730 16216
rect 39764 16182 39798 16216
rect 39832 16182 39866 16216
rect 39900 16182 39934 16216
rect 39968 16182 40002 16216
rect 40036 16182 40070 16216
rect 40104 16182 40138 16216
rect 40172 16182 40206 16216
rect 40240 16182 40274 16216
rect 40308 16182 40342 16216
rect 40376 16182 40410 16216
rect 40444 16182 40478 16216
rect 40512 16182 40546 16216
rect 40580 16182 40614 16216
rect 40648 16182 40682 16216
rect 40716 16182 40750 16216
rect 40784 16182 40818 16216
rect 40852 16182 40886 16216
rect 40920 16182 41165 16216
rect 37706 16131 41165 16182
rect 37706 16058 37839 16131
rect 37706 16024 37749 16058
rect 37783 16024 37839 16058
rect 37706 15990 37839 16024
rect 37706 15956 37749 15990
rect 37783 15956 37839 15990
rect 37706 15922 37839 15956
rect 37706 15888 37749 15922
rect 37783 15888 37839 15922
rect 37706 15854 37839 15888
rect 37706 15820 37749 15854
rect 37783 15820 37839 15854
rect 37706 15786 37839 15820
rect 37706 15752 37749 15786
rect 37783 15752 37839 15786
rect 37706 15718 37839 15752
rect 41047 16018 41165 16131
rect 41047 15984 41089 16018
rect 41123 15984 41165 16018
rect 41047 15950 41165 15984
rect 41047 15916 41089 15950
rect 41123 15916 41165 15950
rect 41047 15882 41165 15916
rect 41047 15848 41089 15882
rect 41123 15848 41165 15882
rect 41047 15814 41165 15848
rect 41047 15780 41089 15814
rect 41123 15780 41165 15814
rect 37706 15684 37749 15718
rect 37783 15684 37839 15718
rect 37706 15650 37839 15684
rect 37706 15616 37749 15650
rect 37783 15616 37839 15650
rect 37706 15582 37839 15616
rect 41047 15746 41165 15780
rect 41047 15712 41089 15746
rect 41123 15712 41165 15746
rect 41047 15678 41165 15712
rect 41047 15644 41089 15678
rect 41123 15644 41165 15678
rect 41047 15610 41165 15644
rect 37706 15548 37749 15582
rect 37783 15548 37839 15582
rect 37706 15514 37839 15548
rect 37706 15480 37749 15514
rect 37783 15480 37839 15514
rect 37706 15446 37839 15480
rect 37706 15412 37749 15446
rect 37783 15412 37839 15446
rect 27650 15354 27684 15388
rect 24460 15286 24494 15320
rect 27650 15286 27684 15320
rect 24460 15182 24494 15252
rect 27650 15182 27684 15252
rect 24460 15148 24559 15182
rect 24593 15148 24627 15182
rect 24661 15148 24695 15182
rect 24729 15148 24763 15182
rect 24797 15148 24831 15182
rect 24865 15148 24899 15182
rect 24933 15148 24967 15182
rect 25001 15148 25035 15182
rect 25069 15148 25103 15182
rect 25137 15148 25171 15182
rect 25205 15148 25239 15182
rect 25273 15148 25307 15182
rect 25341 15148 25375 15182
rect 25409 15148 25443 15182
rect 25477 15148 25511 15182
rect 25545 15148 25579 15182
rect 25613 15148 25647 15182
rect 25681 15148 25715 15182
rect 25749 15148 25783 15182
rect 25817 15148 25851 15182
rect 25885 15148 25919 15182
rect 25953 15148 25987 15182
rect 26021 15148 26055 15182
rect 26089 15148 26123 15182
rect 26157 15148 26191 15182
rect 26225 15148 26259 15182
rect 26293 15148 26327 15182
rect 26361 15148 26395 15182
rect 26429 15148 26463 15182
rect 26497 15148 26531 15182
rect 26565 15148 26599 15182
rect 26633 15148 26667 15182
rect 26701 15148 26735 15182
rect 26769 15148 26803 15182
rect 26837 15148 26871 15182
rect 26905 15148 26939 15182
rect 26973 15148 27007 15182
rect 27041 15148 27075 15182
rect 27109 15148 27143 15182
rect 27177 15148 27211 15182
rect 27245 15148 27279 15182
rect 27313 15148 27347 15182
rect 27381 15148 27415 15182
rect 27449 15148 27483 15182
rect 27517 15148 27551 15182
rect 27585 15148 27684 15182
rect 28834 15358 28960 15392
rect 28994 15358 29028 15392
rect 29062 15358 29096 15392
rect 29130 15358 29164 15392
rect 29198 15358 29232 15392
rect 29266 15358 29300 15392
rect 29334 15358 29368 15392
rect 29402 15358 29436 15392
rect 29470 15358 29504 15392
rect 29538 15358 29572 15392
rect 29606 15358 29640 15392
rect 29674 15358 29800 15392
rect 28834 15275 28868 15358
rect 29766 15275 29800 15358
rect 28834 15207 28868 15241
rect 24297 15074 24398 15130
rect 24297 15040 24331 15074
rect 24365 15040 24398 15074
rect 24297 14984 24398 15040
rect 24297 14950 24331 14984
rect 24365 14950 24398 14984
rect 24297 14894 24398 14950
rect 24297 14860 24331 14894
rect 24365 14860 24398 14894
rect 24297 14804 24398 14860
rect 24297 14770 24331 14804
rect 24365 14770 24398 14804
rect 23110 14680 23144 14714
rect 23178 14680 23211 14714
rect 23110 14665 23211 14680
rect 24297 14714 24398 14770
rect 24297 14680 24331 14714
rect 24365 14680 24398 14714
rect 24297 14665 24398 14680
rect 23110 14630 24398 14665
rect 20382 14566 20497 14600
rect 20531 14566 20565 14600
rect 20599 14566 20633 14600
rect 20667 14566 20701 14600
rect 20735 14566 20769 14600
rect 20803 14566 20837 14600
rect 20871 14566 20905 14600
rect 20939 14566 20973 14600
rect 21007 14566 21041 14600
rect 21075 14566 21109 14600
rect 21143 14566 21177 14600
rect 21211 14566 21245 14600
rect 21279 14566 21313 14600
rect 21347 14566 21381 14600
rect 21415 14566 21449 14600
rect 21483 14566 21517 14600
rect 21551 14566 21666 14600
rect 20382 14474 20416 14566
rect 21632 14474 21666 14566
rect 23110 14596 23240 14630
rect 23274 14596 23330 14630
rect 23364 14596 23420 14630
rect 23454 14596 23510 14630
rect 23544 14596 23600 14630
rect 23634 14596 23690 14630
rect 23724 14596 23780 14630
rect 23814 14596 23870 14630
rect 23904 14596 23960 14630
rect 23994 14596 24050 14630
rect 24084 14596 24140 14630
rect 24174 14596 24230 14630
rect 24264 14596 24398 14630
rect 23110 14564 24398 14596
rect 28834 15139 28868 15173
rect 28834 15071 28868 15105
rect 28834 15003 28868 15037
rect 28834 14935 28868 14969
rect 28834 14867 28868 14901
rect 28834 14799 28868 14833
rect 28834 14731 28868 14765
rect 28834 14663 28868 14697
rect 28834 14595 28868 14629
rect 20382 14406 20416 14440
rect 20382 14338 20416 14372
rect 20382 14270 20416 14304
rect 20382 14202 20416 14236
rect 20382 14134 20416 14168
rect 20382 14066 20416 14100
rect 20382 13998 20416 14032
rect 20382 13930 20416 13964
rect 20382 13862 20416 13896
rect 20382 13794 20416 13828
rect 20382 13726 20416 13760
rect 20382 13658 20416 13692
rect 20382 13590 20416 13624
rect 20382 13522 20416 13556
rect 20382 13454 20416 13488
rect 20382 13386 20416 13420
rect 20382 13318 20416 13352
rect 20382 13250 20416 13284
rect 20382 13182 20416 13216
rect 20382 13114 20416 13148
rect 20382 13046 20416 13080
rect 20382 12978 20416 13012
rect 20382 12910 20416 12944
rect 20382 12842 20416 12876
rect 20382 12774 20416 12808
rect 20382 12706 20416 12740
rect 20382 12638 20416 12672
rect 20382 12570 20416 12604
rect 20382 12502 20416 12536
rect 20382 12434 20416 12468
rect 20382 12366 20416 12400
rect 20382 12298 20416 12332
rect 20382 12230 20416 12264
rect 20382 12162 20416 12196
rect 20382 12094 20416 12128
rect 20382 12026 20416 12060
rect 20382 11958 20416 11992
rect 20382 11890 20416 11924
rect 20382 11822 20416 11856
rect 20382 11754 20416 11788
rect 20382 11686 20416 11720
rect 20382 11618 20416 11652
rect 20382 11550 20416 11584
rect 20382 11482 20416 11516
rect 12782 11299 14070 11334
rect 12782 11276 12912 11299
rect 12782 11242 12816 11276
rect 12850 11265 12912 11276
rect 12946 11265 13002 11299
rect 13036 11265 13092 11299
rect 13126 11265 13182 11299
rect 13216 11265 13272 11299
rect 13306 11265 13362 11299
rect 13396 11265 13452 11299
rect 13486 11265 13542 11299
rect 13576 11265 13632 11299
rect 13666 11265 13722 11299
rect 13756 11265 13812 11299
rect 13846 11265 13902 11299
rect 13936 11276 14070 11299
rect 13936 11265 14003 11276
rect 12850 11242 14003 11265
rect 14037 11242 14070 11276
rect 12782 11233 14070 11242
rect 12782 11186 12883 11233
rect 12782 11152 12816 11186
rect 12850 11152 12883 11186
rect 13969 11186 14070 11233
rect 12782 11096 12883 11152
rect 12782 11062 12816 11096
rect 12850 11062 12883 11096
rect 12782 11006 12883 11062
rect 12782 10972 12816 11006
rect 12850 10972 12883 11006
rect 12782 10916 12883 10972
rect 12782 10882 12816 10916
rect 12850 10882 12883 10916
rect 12782 10826 12883 10882
rect 12782 10792 12816 10826
rect 12850 10792 12883 10826
rect 12782 10736 12883 10792
rect 12782 10702 12816 10736
rect 12850 10702 12883 10736
rect 12782 10646 12883 10702
rect 12782 10612 12816 10646
rect 12850 10612 12883 10646
rect 12782 10556 12883 10612
rect 12782 10522 12816 10556
rect 12850 10522 12883 10556
rect 12782 10466 12883 10522
rect 12782 10432 12816 10466
rect 12850 10432 12883 10466
rect 12782 10376 12883 10432
rect 12782 10342 12816 10376
rect 12850 10342 12883 10376
rect 12782 10286 12883 10342
rect 12782 10252 12816 10286
rect 12850 10252 12883 10286
rect 12782 10196 12883 10252
rect 13969 11152 14003 11186
rect 14037 11152 14070 11186
rect 13969 11096 14070 11152
rect 13969 11062 14003 11096
rect 14037 11062 14070 11096
rect 13969 11006 14070 11062
rect 13969 10972 14003 11006
rect 14037 10972 14070 11006
rect 13969 10916 14070 10972
rect 13969 10882 14003 10916
rect 14037 10882 14070 10916
rect 13969 10826 14070 10882
rect 13969 10792 14003 10826
rect 14037 10792 14070 10826
rect 13969 10736 14070 10792
rect 13969 10702 14003 10736
rect 14037 10702 14070 10736
rect 13969 10646 14070 10702
rect 13969 10612 14003 10646
rect 14037 10612 14070 10646
rect 13969 10556 14070 10612
rect 13969 10522 14003 10556
rect 14037 10522 14070 10556
rect 13969 10466 14070 10522
rect 13969 10432 14003 10466
rect 14037 10432 14070 10466
rect 13969 10376 14070 10432
rect 13969 10342 14003 10376
rect 14037 10342 14070 10376
rect 13969 10286 14070 10342
rect 13969 10252 14003 10286
rect 14037 10252 14070 10286
rect 12782 10162 12816 10196
rect 12850 10162 12883 10196
rect 12782 10147 12883 10162
rect 13969 10196 14070 10252
rect 13969 10162 14003 10196
rect 14037 10162 14070 10196
rect 13969 10147 14070 10162
rect 12782 10112 14070 10147
rect 12782 10078 12912 10112
rect 12946 10078 13002 10112
rect 13036 10078 13092 10112
rect 13126 10078 13182 10112
rect 13216 10078 13272 10112
rect 13306 10078 13362 10112
rect 13396 10078 13452 10112
rect 13486 10078 13542 10112
rect 13576 10078 13632 10112
rect 13666 10078 13722 10112
rect 13756 10078 13812 10112
rect 13846 10078 13902 10112
rect 13936 10078 14070 10112
rect 12782 10046 14070 10078
rect 12782 9809 14070 9844
rect 12782 9786 12912 9809
rect 12782 9752 12816 9786
rect 12850 9775 12912 9786
rect 12946 9775 13002 9809
rect 13036 9775 13092 9809
rect 13126 9775 13182 9809
rect 13216 9775 13272 9809
rect 13306 9775 13362 9809
rect 13396 9775 13452 9809
rect 13486 9775 13542 9809
rect 13576 9775 13632 9809
rect 13666 9775 13722 9809
rect 13756 9775 13812 9809
rect 13846 9775 13902 9809
rect 13936 9786 14070 9809
rect 13936 9775 14003 9786
rect 12850 9752 14003 9775
rect 14037 9752 14070 9786
rect 12782 9743 14070 9752
rect 12782 9696 12883 9743
rect 12782 9662 12816 9696
rect 12850 9662 12883 9696
rect 13969 9696 14070 9743
rect 12782 9606 12883 9662
rect 12782 9572 12816 9606
rect 12850 9572 12883 9606
rect 12782 9516 12883 9572
rect 12782 9482 12816 9516
rect 12850 9482 12883 9516
rect 12782 9426 12883 9482
rect 12782 9392 12816 9426
rect 12850 9392 12883 9426
rect 12782 9336 12883 9392
rect 12782 9302 12816 9336
rect 12850 9302 12883 9336
rect 12782 9246 12883 9302
rect 12782 9212 12816 9246
rect 12850 9212 12883 9246
rect 12782 9156 12883 9212
rect 12782 9122 12816 9156
rect 12850 9122 12883 9156
rect 12782 9066 12883 9122
rect 12782 9032 12816 9066
rect 12850 9032 12883 9066
rect 12782 8976 12883 9032
rect 12782 8942 12816 8976
rect 12850 8942 12883 8976
rect 12782 8886 12883 8942
rect 12782 8852 12816 8886
rect 12850 8852 12883 8886
rect 12782 8796 12883 8852
rect 12782 8762 12816 8796
rect 12850 8762 12883 8796
rect 12782 8706 12883 8762
rect 13969 9662 14003 9696
rect 14037 9662 14070 9696
rect 13969 9606 14070 9662
rect 13969 9572 14003 9606
rect 14037 9572 14070 9606
rect 13969 9516 14070 9572
rect 13969 9482 14003 9516
rect 14037 9482 14070 9516
rect 13969 9426 14070 9482
rect 13969 9392 14003 9426
rect 14037 9392 14070 9426
rect 13969 9336 14070 9392
rect 13969 9302 14003 9336
rect 14037 9302 14070 9336
rect 13969 9246 14070 9302
rect 13969 9212 14003 9246
rect 14037 9212 14070 9246
rect 13969 9156 14070 9212
rect 13969 9122 14003 9156
rect 14037 9122 14070 9156
rect 13969 9066 14070 9122
rect 13969 9032 14003 9066
rect 14037 9032 14070 9066
rect 13969 8976 14070 9032
rect 13969 8942 14003 8976
rect 14037 8942 14070 8976
rect 13969 8886 14070 8942
rect 13969 8852 14003 8886
rect 14037 8852 14070 8886
rect 13969 8796 14070 8852
rect 13969 8762 14003 8796
rect 14037 8762 14070 8796
rect 12782 8672 12816 8706
rect 12850 8672 12883 8706
rect 12782 8657 12883 8672
rect 13969 8706 14070 8762
rect 13969 8672 14003 8706
rect 14037 8672 14070 8706
rect 13969 8657 14070 8672
rect 12782 8622 14070 8657
rect 12782 8588 12912 8622
rect 12946 8588 13002 8622
rect 13036 8588 13092 8622
rect 13126 8588 13182 8622
rect 13216 8588 13272 8622
rect 13306 8588 13362 8622
rect 13396 8588 13452 8622
rect 13486 8588 13542 8622
rect 13576 8588 13632 8622
rect 13666 8588 13722 8622
rect 13756 8588 13812 8622
rect 13846 8588 13902 8622
rect 13936 8588 14070 8622
rect 12782 8556 14070 8588
rect 12772 8399 14060 8434
rect 12772 8376 12902 8399
rect 12772 8342 12806 8376
rect 12840 8365 12902 8376
rect 12936 8365 12992 8399
rect 13026 8365 13082 8399
rect 13116 8365 13172 8399
rect 13206 8365 13262 8399
rect 13296 8365 13352 8399
rect 13386 8365 13442 8399
rect 13476 8365 13532 8399
rect 13566 8365 13622 8399
rect 13656 8365 13712 8399
rect 13746 8365 13802 8399
rect 13836 8365 13892 8399
rect 13926 8376 14060 8399
rect 13926 8365 13993 8376
rect 12840 8342 13993 8365
rect 14027 8342 14060 8376
rect 12772 8333 14060 8342
rect 12772 8286 12873 8333
rect 12772 8252 12806 8286
rect 12840 8252 12873 8286
rect 13959 8286 14060 8333
rect 12772 8196 12873 8252
rect 12772 8162 12806 8196
rect 12840 8162 12873 8196
rect 12772 8106 12873 8162
rect 12772 8072 12806 8106
rect 12840 8072 12873 8106
rect 12772 8016 12873 8072
rect 12772 7982 12806 8016
rect 12840 7982 12873 8016
rect 12772 7926 12873 7982
rect 12772 7892 12806 7926
rect 12840 7892 12873 7926
rect 12772 7836 12873 7892
rect 12772 7802 12806 7836
rect 12840 7802 12873 7836
rect 12772 7746 12873 7802
rect 12772 7712 12806 7746
rect 12840 7712 12873 7746
rect 12772 7656 12873 7712
rect 12772 7622 12806 7656
rect 12840 7622 12873 7656
rect 12772 7566 12873 7622
rect 12772 7532 12806 7566
rect 12840 7532 12873 7566
rect 12772 7476 12873 7532
rect 12772 7442 12806 7476
rect 12840 7442 12873 7476
rect 12772 7386 12873 7442
rect 12772 7352 12806 7386
rect 12840 7352 12873 7386
rect 12772 7296 12873 7352
rect 13959 8252 13993 8286
rect 14027 8252 14060 8286
rect 13959 8196 14060 8252
rect 13959 8162 13993 8196
rect 14027 8162 14060 8196
rect 13959 8106 14060 8162
rect 13959 8072 13993 8106
rect 14027 8072 14060 8106
rect 13959 8016 14060 8072
rect 13959 7982 13993 8016
rect 14027 7982 14060 8016
rect 20382 11414 20416 11448
rect 20382 11346 20416 11380
rect 20382 11278 20416 11312
rect 20382 11210 20416 11244
rect 20382 11142 20416 11176
rect 20382 11074 20416 11108
rect 20382 11006 20416 11040
rect 20382 10938 20416 10972
rect 20382 10870 20416 10904
rect 20382 10802 20416 10836
rect 20382 10734 20416 10768
rect 20382 10666 20416 10700
rect 20382 10598 20416 10632
rect 20382 10530 20416 10564
rect 20382 10462 20416 10496
rect 20382 10394 20416 10428
rect 20382 10326 20416 10360
rect 20382 10258 20416 10292
rect 20382 10190 20416 10224
rect 20382 10122 20416 10156
rect 20382 10054 20416 10088
rect 20382 9986 20416 10020
rect 20382 9918 20416 9952
rect 20382 9850 20416 9884
rect 20382 9782 20416 9816
rect 20382 9714 20416 9748
rect 20382 9646 20416 9680
rect 20382 9578 20416 9612
rect 20382 9510 20416 9544
rect 20382 9442 20416 9476
rect 20382 9374 20416 9408
rect 20382 9306 20416 9340
rect 20382 9238 20416 9272
rect 20382 9170 20416 9204
rect 20382 9102 20416 9136
rect 20382 9034 20416 9068
rect 20382 8966 20416 9000
rect 20382 8898 20416 8932
rect 20382 8830 20416 8864
rect 20382 8762 20416 8796
rect 20382 8694 20416 8728
rect 20382 8626 20416 8660
rect 20382 8558 20416 8592
rect 20382 8490 20416 8524
rect 20382 8422 20416 8456
rect 20382 8354 20416 8388
rect 20382 8286 20416 8320
rect 20382 8218 20416 8252
rect 20382 8150 20416 8184
rect 20382 8082 20416 8116
rect 20382 8014 20416 8048
rect 13959 7926 14060 7982
rect 13959 7892 13993 7926
rect 14027 7892 14060 7926
rect 13959 7836 14060 7892
rect 13959 7802 13993 7836
rect 14027 7802 14060 7836
rect 13959 7746 14060 7802
rect 20382 7946 20416 7980
rect 20382 7878 20416 7912
rect 20382 7810 20416 7844
rect 13959 7712 13993 7746
rect 14027 7712 14060 7746
rect 13959 7656 14060 7712
rect 13959 7622 13993 7656
rect 14027 7622 14060 7656
rect 13959 7566 14060 7622
rect 13959 7532 13993 7566
rect 14027 7532 14060 7566
rect 13959 7476 14060 7532
rect 13959 7442 13993 7476
rect 14027 7442 14060 7476
rect 13959 7386 14060 7442
rect 13959 7352 13993 7386
rect 14027 7352 14060 7386
rect 12772 7262 12806 7296
rect 12840 7262 12873 7296
rect 12772 7247 12873 7262
rect 13959 7296 14060 7352
rect 13959 7262 13993 7296
rect 14027 7262 14060 7296
rect 13959 7247 14060 7262
rect 12772 7212 14060 7247
rect 12772 7178 12902 7212
rect 12936 7178 12992 7212
rect 13026 7178 13082 7212
rect 13116 7178 13172 7212
rect 13206 7178 13262 7212
rect 13296 7178 13352 7212
rect 13386 7178 13442 7212
rect 13476 7178 13532 7212
rect 13566 7178 13622 7212
rect 13656 7178 13712 7212
rect 13746 7178 13802 7212
rect 13836 7178 13892 7212
rect 13926 7178 14060 7212
rect 12772 7146 14060 7178
rect 16080 7206 16206 7240
rect 16240 7206 16274 7240
rect 16308 7206 16342 7240
rect 16376 7206 16410 7240
rect 16444 7206 16478 7240
rect 16512 7206 16546 7240
rect 16580 7206 16614 7240
rect 16648 7206 16682 7240
rect 16716 7206 16750 7240
rect 16784 7206 16818 7240
rect 16852 7206 16886 7240
rect 16920 7206 17046 7240
rect 16080 7119 16114 7206
rect 12772 7049 14060 7084
rect 12772 7026 12902 7049
rect 12772 6992 12806 7026
rect 12840 7015 12902 7026
rect 12936 7015 12992 7049
rect 13026 7015 13082 7049
rect 13116 7015 13172 7049
rect 13206 7015 13262 7049
rect 13296 7015 13352 7049
rect 13386 7015 13442 7049
rect 13476 7015 13532 7049
rect 13566 7015 13622 7049
rect 13656 7015 13712 7049
rect 13746 7015 13802 7049
rect 13836 7015 13892 7049
rect 13926 7026 14060 7049
rect 13926 7015 13993 7026
rect 12840 6992 13993 7015
rect 14027 6992 14060 7026
rect 12772 6983 14060 6992
rect 12772 6936 12873 6983
rect 12772 6902 12806 6936
rect 12840 6902 12873 6936
rect 13959 6936 14060 6983
rect 12772 6846 12873 6902
rect 12772 6812 12806 6846
rect 12840 6812 12873 6846
rect 12772 6756 12873 6812
rect 12772 6722 12806 6756
rect 12840 6722 12873 6756
rect 12772 6666 12873 6722
rect 12772 6632 12806 6666
rect 12840 6632 12873 6666
rect 12772 6576 12873 6632
rect 12772 6542 12806 6576
rect 12840 6542 12873 6576
rect 12772 6486 12873 6542
rect 12772 6452 12806 6486
rect 12840 6452 12873 6486
rect 12772 6396 12873 6452
rect 12772 6362 12806 6396
rect 12840 6362 12873 6396
rect 12772 6306 12873 6362
rect 12772 6272 12806 6306
rect 12840 6272 12873 6306
rect 12772 6216 12873 6272
rect 12772 6182 12806 6216
rect 12840 6182 12873 6216
rect 12772 6126 12873 6182
rect 12772 6092 12806 6126
rect 12840 6092 12873 6126
rect 12772 6036 12873 6092
rect 12772 6002 12806 6036
rect 12840 6002 12873 6036
rect 12772 5946 12873 6002
rect 13959 6902 13993 6936
rect 14027 6902 14060 6936
rect 13959 6846 14060 6902
rect 13959 6812 13993 6846
rect 14027 6812 14060 6846
rect 13959 6756 14060 6812
rect 13959 6722 13993 6756
rect 14027 6722 14060 6756
rect 13959 6666 14060 6722
rect 13959 6632 13993 6666
rect 14027 6632 14060 6666
rect 13959 6576 14060 6632
rect 13959 6542 13993 6576
rect 14027 6542 14060 6576
rect 13959 6486 14060 6542
rect 13959 6452 13993 6486
rect 14027 6452 14060 6486
rect 13959 6396 14060 6452
rect 13959 6362 13993 6396
rect 14027 6362 14060 6396
rect 13959 6306 14060 6362
rect 13959 6272 13993 6306
rect 14027 6272 14060 6306
rect 13959 6216 14060 6272
rect 13959 6182 13993 6216
rect 14027 6182 14060 6216
rect 13959 6126 14060 6182
rect 13959 6092 13993 6126
rect 14027 6092 14060 6126
rect 13959 6036 14060 6092
rect 13959 6002 13993 6036
rect 14027 6002 14060 6036
rect 12772 5912 12806 5946
rect 12840 5912 12873 5946
rect 12772 5897 12873 5912
rect 13959 5946 14060 6002
rect 13959 5912 13993 5946
rect 14027 5912 14060 5946
rect 13959 5897 14060 5912
rect 12772 5862 14060 5897
rect 12772 5828 12902 5862
rect 12936 5828 12992 5862
rect 13026 5828 13082 5862
rect 13116 5828 13172 5862
rect 13206 5828 13262 5862
rect 13296 5828 13352 5862
rect 13386 5828 13442 5862
rect 13476 5828 13532 5862
rect 13566 5828 13622 5862
rect 13656 5828 13712 5862
rect 13746 5828 13802 5862
rect 13836 5828 13892 5862
rect 13926 5828 14060 5862
rect 12772 5796 14060 5828
rect 14422 7079 15710 7114
rect 14422 7056 14552 7079
rect 14422 7022 14456 7056
rect 14490 7045 14552 7056
rect 14586 7045 14642 7079
rect 14676 7045 14732 7079
rect 14766 7045 14822 7079
rect 14856 7045 14912 7079
rect 14946 7045 15002 7079
rect 15036 7045 15092 7079
rect 15126 7045 15182 7079
rect 15216 7045 15272 7079
rect 15306 7045 15362 7079
rect 15396 7045 15452 7079
rect 15486 7045 15542 7079
rect 15576 7056 15710 7079
rect 15576 7045 15643 7056
rect 14490 7022 15643 7045
rect 15677 7022 15710 7056
rect 14422 7013 15710 7022
rect 14422 6966 14523 7013
rect 14422 6932 14456 6966
rect 14490 6932 14523 6966
rect 15609 6966 15710 7013
rect 14422 6876 14523 6932
rect 14422 6842 14456 6876
rect 14490 6842 14523 6876
rect 14422 6786 14523 6842
rect 14422 6752 14456 6786
rect 14490 6752 14523 6786
rect 14422 6696 14523 6752
rect 14422 6662 14456 6696
rect 14490 6662 14523 6696
rect 14422 6606 14523 6662
rect 14422 6572 14456 6606
rect 14490 6572 14523 6606
rect 14422 6516 14523 6572
rect 14422 6482 14456 6516
rect 14490 6482 14523 6516
rect 14422 6426 14523 6482
rect 14422 6392 14456 6426
rect 14490 6392 14523 6426
rect 14422 6336 14523 6392
rect 14422 6302 14456 6336
rect 14490 6302 14523 6336
rect 14422 6246 14523 6302
rect 14422 6212 14456 6246
rect 14490 6212 14523 6246
rect 14422 6156 14523 6212
rect 14422 6122 14456 6156
rect 14490 6122 14523 6156
rect 14422 6066 14523 6122
rect 14422 6032 14456 6066
rect 14490 6032 14523 6066
rect 14422 5976 14523 6032
rect 15609 6932 15643 6966
rect 15677 6932 15710 6966
rect 15609 6876 15710 6932
rect 15609 6842 15643 6876
rect 15677 6842 15710 6876
rect 15609 6786 15710 6842
rect 15609 6752 15643 6786
rect 15677 6752 15710 6786
rect 15609 6696 15710 6752
rect 15609 6662 15643 6696
rect 15677 6662 15710 6696
rect 15609 6606 15710 6662
rect 15609 6572 15643 6606
rect 15677 6572 15710 6606
rect 15609 6516 15710 6572
rect 15609 6482 15643 6516
rect 15677 6482 15710 6516
rect 15609 6426 15710 6482
rect 15609 6392 15643 6426
rect 15677 6392 15710 6426
rect 15609 6336 15710 6392
rect 15609 6302 15643 6336
rect 15677 6302 15710 6336
rect 15609 6246 15710 6302
rect 15609 6212 15643 6246
rect 15677 6212 15710 6246
rect 15609 6156 15710 6212
rect 15609 6122 15643 6156
rect 15677 6122 15710 6156
rect 15609 6066 15710 6122
rect 15609 6032 15643 6066
rect 15677 6032 15710 6066
rect 14422 5942 14456 5976
rect 14490 5942 14523 5976
rect 14422 5927 14523 5942
rect 15609 5976 15710 6032
rect 15609 5942 15643 5976
rect 15677 5942 15710 5976
rect 15609 5927 15710 5942
rect 14422 5892 15710 5927
rect 14422 5858 14552 5892
rect 14586 5858 14642 5892
rect 14676 5858 14732 5892
rect 14766 5858 14822 5892
rect 14856 5858 14912 5892
rect 14946 5858 15002 5892
rect 15036 5858 15092 5892
rect 15126 5858 15182 5892
rect 15216 5858 15272 5892
rect 15306 5858 15362 5892
rect 15396 5858 15452 5892
rect 15486 5858 15542 5892
rect 15576 5858 15710 5892
rect 14422 5826 15710 5858
rect 17012 7119 17046 7206
rect 16080 7051 16114 7085
rect 16080 6983 16114 7017
rect 16080 6915 16114 6949
rect 16080 6847 16114 6881
rect 16080 6779 16114 6813
rect 16080 6711 16114 6745
rect 16080 6643 16114 6677
rect 16080 6575 16114 6609
rect 16080 6507 16114 6541
rect 16080 6439 16114 6473
rect 16080 6371 16114 6405
rect 16080 6303 16114 6337
rect 16080 6235 16114 6269
rect 16080 6167 16114 6201
rect 16080 6099 16114 6133
rect 16080 6031 16114 6065
rect 16080 5963 16114 5997
rect 16080 5895 16114 5929
rect 16080 5827 16114 5861
rect 16080 5759 16114 5793
rect 12772 5699 14060 5734
rect 12772 5676 12902 5699
rect 12772 5642 12806 5676
rect 12840 5665 12902 5676
rect 12936 5665 12992 5699
rect 13026 5665 13082 5699
rect 13116 5665 13172 5699
rect 13206 5665 13262 5699
rect 13296 5665 13352 5699
rect 13386 5665 13442 5699
rect 13476 5665 13532 5699
rect 13566 5665 13622 5699
rect 13656 5665 13712 5699
rect 13746 5665 13802 5699
rect 13836 5665 13892 5699
rect 13926 5676 14060 5699
rect 13926 5665 13993 5676
rect 12840 5642 13993 5665
rect 14027 5642 14060 5676
rect 12772 5633 14060 5642
rect 12772 5586 12873 5633
rect 12772 5552 12806 5586
rect 12840 5552 12873 5586
rect 13959 5586 14060 5633
rect 12772 5496 12873 5552
rect 12772 5462 12806 5496
rect 12840 5462 12873 5496
rect 12772 5406 12873 5462
rect 12772 5372 12806 5406
rect 12840 5372 12873 5406
rect 12772 5316 12873 5372
rect 12772 5282 12806 5316
rect 12840 5282 12873 5316
rect 12772 5226 12873 5282
rect 12772 5192 12806 5226
rect 12840 5192 12873 5226
rect 12772 5136 12873 5192
rect 12772 5102 12806 5136
rect 12840 5102 12873 5136
rect 12772 5046 12873 5102
rect 12772 5012 12806 5046
rect 12840 5012 12873 5046
rect 12772 4956 12873 5012
rect 12772 4922 12806 4956
rect 12840 4922 12873 4956
rect 12772 4866 12873 4922
rect 12772 4832 12806 4866
rect 12840 4832 12873 4866
rect 12772 4776 12873 4832
rect 12772 4742 12806 4776
rect 12840 4742 12873 4776
rect 12772 4686 12873 4742
rect 12772 4652 12806 4686
rect 12840 4652 12873 4686
rect 12772 4596 12873 4652
rect 13959 5552 13993 5586
rect 14027 5552 14060 5586
rect 13959 5496 14060 5552
rect 13959 5462 13993 5496
rect 14027 5462 14060 5496
rect 13959 5406 14060 5462
rect 13959 5372 13993 5406
rect 14027 5372 14060 5406
rect 13959 5316 14060 5372
rect 13959 5282 13993 5316
rect 14027 5282 14060 5316
rect 13959 5226 14060 5282
rect 13959 5192 13993 5226
rect 14027 5192 14060 5226
rect 13959 5136 14060 5192
rect 13959 5102 13993 5136
rect 14027 5102 14060 5136
rect 13959 5046 14060 5102
rect 13959 5012 13993 5046
rect 14027 5012 14060 5046
rect 13959 4956 14060 5012
rect 13959 4922 13993 4956
rect 14027 4922 14060 4956
rect 13959 4866 14060 4922
rect 13959 4832 13993 4866
rect 14027 4832 14060 4866
rect 13959 4776 14060 4832
rect 13959 4742 13993 4776
rect 14027 4742 14060 4776
rect 13959 4686 14060 4742
rect 13959 4652 13993 4686
rect 14027 4652 14060 4686
rect 12772 4562 12806 4596
rect 12840 4562 12873 4596
rect 12772 4547 12873 4562
rect 13959 4596 14060 4652
rect 13959 4562 13993 4596
rect 14027 4562 14060 4596
rect 13959 4547 14060 4562
rect 12772 4512 14060 4547
rect 12772 4478 12902 4512
rect 12936 4478 12992 4512
rect 13026 4478 13082 4512
rect 13116 4478 13172 4512
rect 13206 4478 13262 4512
rect 13296 4478 13352 4512
rect 13386 4478 13442 4512
rect 13476 4478 13532 4512
rect 13566 4478 13622 4512
rect 13656 4478 13712 4512
rect 13746 4478 13802 4512
rect 13836 4478 13892 4512
rect 13926 4478 14060 4512
rect 12772 4446 14060 4478
rect 14422 5719 15710 5754
rect 14422 5696 14552 5719
rect 14422 5662 14456 5696
rect 14490 5685 14552 5696
rect 14586 5685 14642 5719
rect 14676 5685 14732 5719
rect 14766 5685 14822 5719
rect 14856 5685 14912 5719
rect 14946 5685 15002 5719
rect 15036 5685 15092 5719
rect 15126 5685 15182 5719
rect 15216 5685 15272 5719
rect 15306 5685 15362 5719
rect 15396 5685 15452 5719
rect 15486 5685 15542 5719
rect 15576 5696 15710 5719
rect 15576 5685 15643 5696
rect 14490 5662 15643 5685
rect 15677 5662 15710 5696
rect 14422 5653 15710 5662
rect 14422 5606 14523 5653
rect 14422 5572 14456 5606
rect 14490 5572 14523 5606
rect 15609 5606 15710 5653
rect 14422 5516 14523 5572
rect 14422 5482 14456 5516
rect 14490 5482 14523 5516
rect 14422 5426 14523 5482
rect 14422 5392 14456 5426
rect 14490 5392 14523 5426
rect 14422 5336 14523 5392
rect 14422 5302 14456 5336
rect 14490 5302 14523 5336
rect 14422 5246 14523 5302
rect 14422 5212 14456 5246
rect 14490 5212 14523 5246
rect 14422 5156 14523 5212
rect 14422 5122 14456 5156
rect 14490 5122 14523 5156
rect 14422 5066 14523 5122
rect 14422 5032 14456 5066
rect 14490 5032 14523 5066
rect 14422 4976 14523 5032
rect 14422 4942 14456 4976
rect 14490 4942 14523 4976
rect 14422 4886 14523 4942
rect 14422 4852 14456 4886
rect 14490 4852 14523 4886
rect 14422 4796 14523 4852
rect 14422 4762 14456 4796
rect 14490 4762 14523 4796
rect 14422 4706 14523 4762
rect 14422 4672 14456 4706
rect 14490 4672 14523 4706
rect 14422 4616 14523 4672
rect 15609 5572 15643 5606
rect 15677 5572 15710 5606
rect 15609 5516 15710 5572
rect 15609 5482 15643 5516
rect 15677 5482 15710 5516
rect 15609 5426 15710 5482
rect 15609 5392 15643 5426
rect 15677 5392 15710 5426
rect 15609 5336 15710 5392
rect 15609 5302 15643 5336
rect 15677 5302 15710 5336
rect 15609 5246 15710 5302
rect 15609 5212 15643 5246
rect 15677 5212 15710 5246
rect 15609 5156 15710 5212
rect 15609 5122 15643 5156
rect 15677 5122 15710 5156
rect 15609 5066 15710 5122
rect 15609 5032 15643 5066
rect 15677 5032 15710 5066
rect 15609 4976 15710 5032
rect 15609 4942 15643 4976
rect 15677 4942 15710 4976
rect 15609 4886 15710 4942
rect 15609 4852 15643 4886
rect 15677 4852 15710 4886
rect 15609 4796 15710 4852
rect 15609 4762 15643 4796
rect 15677 4762 15710 4796
rect 15609 4706 15710 4762
rect 15609 4672 15643 4706
rect 15677 4672 15710 4706
rect 14422 4582 14456 4616
rect 14490 4582 14523 4616
rect 14422 4567 14523 4582
rect 15609 4616 15710 4672
rect 15609 4582 15643 4616
rect 15677 4582 15710 4616
rect 15609 4567 15710 4582
rect 14422 4532 15710 4567
rect 14422 4498 14552 4532
rect 14586 4498 14642 4532
rect 14676 4498 14732 4532
rect 14766 4498 14822 4532
rect 14856 4498 14912 4532
rect 14946 4498 15002 4532
rect 15036 4498 15092 4532
rect 15126 4498 15182 4532
rect 15216 4498 15272 4532
rect 15306 4498 15362 4532
rect 15396 4498 15452 4532
rect 15486 4498 15542 4532
rect 15576 4498 15710 4532
rect 16080 5691 16114 5725
rect 16080 5623 16114 5657
rect 16080 5555 16114 5589
rect 16080 5487 16114 5521
rect 16080 5419 16114 5453
rect 16080 5351 16114 5385
rect 16080 5283 16114 5317
rect 16080 5215 16114 5249
rect 16080 5147 16114 5181
rect 16080 5079 16114 5113
rect 16080 5011 16114 5045
rect 16080 4943 16114 4977
rect 16080 4875 16114 4909
rect 16080 4807 16114 4841
rect 16080 4739 16114 4773
rect 16080 4671 16114 4705
rect 17012 7051 17046 7085
rect 17012 6983 17046 7017
rect 17012 6915 17046 6949
rect 17012 6847 17046 6881
rect 17012 6779 17046 6813
rect 17012 6711 17046 6745
rect 17012 6643 17046 6677
rect 17012 6575 17046 6609
rect 17012 6507 17046 6541
rect 17012 6439 17046 6473
rect 17012 6371 17046 6405
rect 17012 6303 17046 6337
rect 17012 6235 17046 6269
rect 17012 6167 17046 6201
rect 17012 6099 17046 6133
rect 17012 6031 17046 6065
rect 17012 5963 17046 5997
rect 17012 5895 17046 5929
rect 17012 5827 17046 5861
rect 17012 5759 17046 5793
rect 17012 5691 17046 5725
rect 17012 5623 17046 5657
rect 17012 5555 17046 5589
rect 17012 5487 17046 5521
rect 17012 5419 17046 5453
rect 17012 5351 17046 5385
rect 17012 5283 17046 5317
rect 17012 5215 17046 5249
rect 17012 5147 17046 5181
rect 17012 5079 17046 5113
rect 17012 5011 17046 5045
rect 17012 4943 17046 4977
rect 17012 4875 17046 4909
rect 17012 4807 17046 4841
rect 17012 4739 17046 4773
rect 17012 4671 17046 4705
rect 16080 4550 16114 4637
rect 17012 4550 17046 4637
rect 16080 4516 16206 4550
rect 16240 4516 16274 4550
rect 16308 4516 16342 4550
rect 16376 4516 16410 4550
rect 16444 4516 16478 4550
rect 16512 4516 16546 4550
rect 16580 4516 16614 4550
rect 16648 4516 16682 4550
rect 16716 4516 16750 4550
rect 16784 4516 16818 4550
rect 16852 4516 16886 4550
rect 16920 4516 17046 4550
rect 14422 4466 15710 4498
rect 20382 7742 20416 7776
rect 20382 7674 20416 7708
rect 20382 7606 20416 7640
rect 20382 7538 20416 7572
rect 20382 7470 20416 7504
rect 20382 7402 20416 7436
rect 20382 7334 20416 7368
rect 20382 7266 20416 7300
rect 20382 7198 20416 7232
rect 20382 7130 20416 7164
rect 20382 7062 20416 7096
rect 20382 6994 20416 7028
rect 20382 6926 20416 6960
rect 20382 6858 20416 6892
rect 20382 6790 20416 6824
rect 20382 6722 20416 6756
rect 20382 6654 20416 6688
rect 20382 6586 20416 6620
rect 20382 6518 20416 6552
rect 20382 6450 20416 6484
rect 20382 6382 20416 6416
rect 20382 6314 20416 6348
rect 20382 6246 20416 6280
rect 20382 6178 20416 6212
rect 20382 6110 20416 6144
rect 20382 6042 20416 6076
rect 20382 5974 20416 6008
rect 20382 5906 20416 5940
rect 20382 5838 20416 5872
rect 20382 5770 20416 5804
rect 20382 5702 20416 5736
rect 20382 5634 20416 5668
rect 20382 5566 20416 5600
rect 20382 5498 20416 5532
rect 20382 5430 20416 5464
rect 20382 5362 20416 5396
rect 20382 5294 20416 5328
rect 20382 5226 20416 5260
rect 20382 5158 20416 5192
rect 20382 5090 20416 5124
rect 20382 5022 20416 5056
rect 20382 4954 20416 4988
rect 20382 4886 20416 4920
rect 20382 4818 20416 4852
rect 20382 4750 20416 4784
rect 21632 14406 21666 14440
rect 21632 14338 21666 14372
rect 21632 14270 21666 14304
rect 21632 14202 21666 14236
rect 21632 14134 21666 14168
rect 21632 14066 21666 14100
rect 21632 13998 21666 14032
rect 21632 13930 21666 13964
rect 21632 13862 21666 13896
rect 21632 13794 21666 13828
rect 21632 13726 21666 13760
rect 21632 13658 21666 13692
rect 28834 14527 28868 14561
rect 28834 14459 28868 14493
rect 28834 14391 28868 14425
rect 28834 14323 28868 14357
rect 28834 14255 28868 14289
rect 28834 14187 28868 14221
rect 28834 14119 28868 14153
rect 28834 14051 28868 14085
rect 28834 13983 28868 14017
rect 28834 13915 28868 13949
rect 28834 13847 28868 13881
rect 28834 13779 28868 13813
rect 29766 15207 29800 15241
rect 29766 15139 29800 15173
rect 29766 15071 29800 15105
rect 29766 15003 29800 15037
rect 29766 14935 29800 14969
rect 29766 14867 29800 14901
rect 29766 14799 29800 14833
rect 29766 14731 29800 14765
rect 29766 14663 29800 14697
rect 29766 14595 29800 14629
rect 29766 14527 29800 14561
rect 29766 14459 29800 14493
rect 29766 14391 29800 14425
rect 29766 14323 29800 14357
rect 29766 14255 29800 14289
rect 29766 14187 29800 14221
rect 29766 14119 29800 14153
rect 29766 14051 29800 14085
rect 29766 13983 29800 14017
rect 29766 13915 29800 13949
rect 29766 13847 29800 13881
rect 29766 13779 29800 13813
rect 28834 13662 28868 13745
rect 29766 13662 29800 13745
rect 28834 13628 28960 13662
rect 28994 13628 29028 13662
rect 29062 13628 29096 13662
rect 29130 13628 29164 13662
rect 29198 13628 29232 13662
rect 29266 13628 29300 13662
rect 29334 13628 29368 13662
rect 29402 13628 29436 13662
rect 29470 13628 29504 13662
rect 29538 13628 29572 13662
rect 29606 13628 29640 13662
rect 29674 13628 29800 13662
rect 37706 15378 37839 15412
rect 37706 15344 37749 15378
rect 37783 15344 37839 15378
rect 37706 15310 37839 15344
rect 37706 15276 37749 15310
rect 37783 15276 37839 15310
rect 37706 15242 37839 15276
rect 37706 15208 37749 15242
rect 37783 15208 37839 15242
rect 37706 15174 37839 15208
rect 37706 15140 37749 15174
rect 37783 15140 37839 15174
rect 37706 15106 37839 15140
rect 37706 15072 37749 15106
rect 37783 15072 37839 15106
rect 37706 15038 37839 15072
rect 37706 15004 37749 15038
rect 37783 15004 37839 15038
rect 37706 14970 37839 15004
rect 37706 14936 37749 14970
rect 37783 14936 37839 14970
rect 37706 14902 37839 14936
rect 37706 14868 37749 14902
rect 37783 14868 37839 14902
rect 37706 14834 37839 14868
rect 37706 14800 37749 14834
rect 37783 14800 37839 14834
rect 37706 14766 37839 14800
rect 37706 14732 37749 14766
rect 37783 14732 37839 14766
rect 37706 14698 37839 14732
rect 37706 14664 37749 14698
rect 37783 14664 37839 14698
rect 37706 14630 37839 14664
rect 37706 14596 37749 14630
rect 37783 14596 37839 14630
rect 37706 14562 37839 14596
rect 37706 14528 37749 14562
rect 37783 14528 37839 14562
rect 37706 14494 37839 14528
rect 37706 14460 37749 14494
rect 37783 14460 37839 14494
rect 37706 14426 37839 14460
rect 37706 14392 37749 14426
rect 37783 14392 37839 14426
rect 37706 14358 37839 14392
rect 37706 14324 37749 14358
rect 37783 14324 37839 14358
rect 37706 14290 37839 14324
rect 37706 14256 37749 14290
rect 37783 14256 37839 14290
rect 37706 14222 37839 14256
rect 37706 14188 37749 14222
rect 37783 14188 37839 14222
rect 37706 14154 37839 14188
rect 37706 14120 37749 14154
rect 37783 14120 37839 14154
rect 37706 14086 37839 14120
rect 37706 14052 37749 14086
rect 37783 14052 37839 14086
rect 37706 14018 37839 14052
rect 37706 13984 37749 14018
rect 37783 13984 37839 14018
rect 37706 13950 37839 13984
rect 37706 13916 37749 13950
rect 37783 13916 37839 13950
rect 37706 13882 37839 13916
rect 37706 13848 37749 13882
rect 37783 13848 37839 13882
rect 37706 13814 37839 13848
rect 37706 13780 37749 13814
rect 37783 13780 37839 13814
rect 37706 13746 37839 13780
rect 37706 13712 37749 13746
rect 37783 13712 37839 13746
rect 37706 13678 37839 13712
rect 37706 13644 37749 13678
rect 37783 13644 37839 13678
rect 21632 13590 21666 13624
rect 21632 13522 21666 13556
rect 37706 13610 37839 13644
rect 37706 13576 37749 13610
rect 37783 13576 37839 13610
rect 41047 15576 41089 15610
rect 41123 15576 41165 15610
rect 41047 15542 41165 15576
rect 41047 15508 41089 15542
rect 41123 15508 41165 15542
rect 41047 15474 41165 15508
rect 41047 15440 41089 15474
rect 41123 15440 41165 15474
rect 41047 15406 41165 15440
rect 41047 15372 41089 15406
rect 41123 15372 41165 15406
rect 41047 15338 41165 15372
rect 41047 15304 41089 15338
rect 41123 15304 41165 15338
rect 41047 15270 41165 15304
rect 41047 15236 41089 15270
rect 41123 15236 41165 15270
rect 41047 15202 41165 15236
rect 41047 15168 41089 15202
rect 41123 15168 41165 15202
rect 41047 15134 41165 15168
rect 41047 15100 41089 15134
rect 41123 15100 41165 15134
rect 41047 15066 41165 15100
rect 41047 15032 41089 15066
rect 41123 15032 41165 15066
rect 41047 14998 41165 15032
rect 41047 14964 41089 14998
rect 41123 14964 41165 14998
rect 41047 14930 41165 14964
rect 41047 14896 41089 14930
rect 41123 14896 41165 14930
rect 41047 14862 41165 14896
rect 41047 14828 41089 14862
rect 41123 14828 41165 14862
rect 41047 14794 41165 14828
rect 41047 14760 41089 14794
rect 41123 14760 41165 14794
rect 41047 14726 41165 14760
rect 41047 14692 41089 14726
rect 41123 14692 41165 14726
rect 41047 14658 41165 14692
rect 41047 14624 41089 14658
rect 41123 14624 41165 14658
rect 41047 14590 41165 14624
rect 41047 14556 41089 14590
rect 41123 14556 41165 14590
rect 41047 14522 41165 14556
rect 41047 14488 41089 14522
rect 41123 14488 41165 14522
rect 41047 14454 41165 14488
rect 41047 14420 41089 14454
rect 41123 14420 41165 14454
rect 41047 14386 41165 14420
rect 41047 14352 41089 14386
rect 41123 14352 41165 14386
rect 41047 14318 41165 14352
rect 41047 14284 41089 14318
rect 41123 14284 41165 14318
rect 41047 14250 41165 14284
rect 41047 14216 41089 14250
rect 41123 14216 41165 14250
rect 41047 14182 41165 14216
rect 41047 14148 41089 14182
rect 41123 14148 41165 14182
rect 41047 14114 41165 14148
rect 41047 14080 41089 14114
rect 41123 14080 41165 14114
rect 41047 14046 41165 14080
rect 41047 14012 41089 14046
rect 41123 14012 41165 14046
rect 41047 13978 41165 14012
rect 41047 13944 41089 13978
rect 41123 13944 41165 13978
rect 41047 13910 41165 13944
rect 41047 13876 41089 13910
rect 41123 13876 41165 13910
rect 41047 13842 41165 13876
rect 41047 13808 41089 13842
rect 41123 13808 41165 13842
rect 41047 13774 41165 13808
rect 41047 13740 41089 13774
rect 41123 13740 41165 13774
rect 41047 13706 41165 13740
rect 41047 13672 41089 13706
rect 41123 13672 41165 13706
rect 41047 13638 41165 13672
rect 41047 13604 41089 13638
rect 41123 13604 41165 13638
rect 37706 13542 37839 13576
rect 41047 13570 41165 13604
rect 37706 13508 37749 13542
rect 37783 13508 37839 13542
rect 21632 13454 21666 13488
rect 21632 13386 21666 13420
rect 21632 13318 21666 13352
rect 21632 13250 21666 13284
rect 21632 13182 21666 13216
rect 21632 13114 21666 13148
rect 21632 13046 21666 13080
rect 21632 12978 21666 13012
rect 21632 12910 21666 12944
rect 21632 12842 21666 12876
rect 21632 12774 21666 12808
rect 21632 12706 21666 12740
rect 21632 12638 21666 12672
rect 21632 12570 21666 12604
rect 21632 12502 21666 12536
rect 21632 12434 21666 12468
rect 21632 12366 21666 12400
rect 21632 12298 21666 12332
rect 21632 12230 21666 12264
rect 21632 12162 21666 12196
rect 21632 12094 21666 12128
rect 37706 13474 37839 13508
rect 21632 12026 21666 12060
rect 21632 11958 21666 11992
rect 21632 11890 21666 11924
rect 21632 11822 21666 11856
rect 21632 11754 21666 11788
rect 21632 11686 21666 11720
rect 21632 11618 21666 11652
rect 21632 11550 21666 11584
rect 21632 11482 21666 11516
rect 21632 11414 21666 11448
rect 21632 11346 21666 11380
rect 21632 11278 21666 11312
rect 21632 11210 21666 11244
rect 21632 11142 21666 11176
rect 21632 11074 21666 11108
rect 21632 11006 21666 11040
rect 21632 10938 21666 10972
rect 21632 10870 21666 10904
rect 21632 10802 21666 10836
rect 21632 10734 21666 10768
rect 21632 10666 21666 10700
rect 21632 10598 21666 10632
rect 21632 10530 21666 10564
rect 21632 10462 21666 10496
rect 21632 10394 21666 10428
rect 21632 10326 21666 10360
rect 21632 10258 21666 10292
rect 21632 10190 21666 10224
rect 21632 10122 21666 10156
rect 21632 10054 21666 10088
rect 21632 9986 21666 10020
rect 21632 9918 21666 9952
rect 21632 9850 21666 9884
rect 21632 9782 21666 9816
rect 21632 9714 21666 9748
rect 21632 9646 21666 9680
rect 21632 9578 21666 9612
rect 21632 9510 21666 9544
rect 21632 9442 21666 9476
rect 21632 9374 21666 9408
rect 21632 9306 21666 9340
rect 21632 9238 21666 9272
rect 21632 9170 21666 9204
rect 21632 9102 21666 9136
rect 21632 9034 21666 9068
rect 21632 8966 21666 9000
rect 26398 13440 26524 13474
rect 26558 13440 26592 13474
rect 26626 13440 26660 13474
rect 26694 13440 26728 13474
rect 26762 13440 26796 13474
rect 26830 13440 26864 13474
rect 26898 13440 26932 13474
rect 26966 13440 27000 13474
rect 27034 13440 27068 13474
rect 27102 13440 27136 13474
rect 27170 13440 27204 13474
rect 27238 13440 27364 13474
rect 26398 13363 26432 13440
rect 27330 13363 27364 13440
rect 26398 13295 26432 13329
rect 26398 13227 26432 13261
rect 26398 13159 26432 13193
rect 26398 13091 26432 13125
rect 26398 13023 26432 13057
rect 26398 12955 26432 12989
rect 26398 12887 26432 12921
rect 26398 12819 26432 12853
rect 26398 12751 26432 12785
rect 26398 12683 26432 12717
rect 26398 12615 26432 12649
rect 26398 12547 26432 12581
rect 26398 12479 26432 12513
rect 26398 12411 26432 12445
rect 26398 12343 26432 12377
rect 26398 12275 26432 12309
rect 26398 12207 26432 12241
rect 26398 12139 26432 12173
rect 26398 12071 26432 12105
rect 26398 12003 26432 12037
rect 26398 11935 26432 11969
rect 26398 11867 26432 11901
rect 26398 11799 26432 11833
rect 26398 11731 26432 11765
rect 26398 11663 26432 11697
rect 26398 11595 26432 11629
rect 26398 11527 26432 11561
rect 26398 11459 26432 11493
rect 26398 11391 26432 11425
rect 26398 11323 26432 11357
rect 26398 11255 26432 11289
rect 26398 11187 26432 11221
rect 26398 11119 26432 11153
rect 26398 11051 26432 11085
rect 26398 10983 26432 11017
rect 26398 10915 26432 10949
rect 26398 10847 26432 10881
rect 26398 10779 26432 10813
rect 26398 10711 26432 10745
rect 26398 10643 26432 10677
rect 26398 10575 26432 10609
rect 26398 10507 26432 10541
rect 26398 10439 26432 10473
rect 26398 10371 26432 10405
rect 26398 10303 26432 10337
rect 26398 10235 26432 10269
rect 26398 10167 26432 10201
rect 26398 10099 26432 10133
rect 26398 10031 26432 10065
rect 26398 9963 26432 9997
rect 26398 9895 26432 9929
rect 26398 9827 26432 9861
rect 26398 9759 26432 9793
rect 26398 9691 26432 9725
rect 26398 9623 26432 9657
rect 26398 9555 26432 9589
rect 26398 9487 26432 9521
rect 26398 9419 26432 9453
rect 26398 9351 26432 9385
rect 26398 9283 26432 9317
rect 26398 9215 26432 9249
rect 26398 9147 26432 9181
rect 26398 9079 26432 9113
rect 26398 9011 26432 9045
rect 26398 8943 26432 8977
rect 21632 8898 21666 8932
rect 21632 8830 21666 8864
rect 21632 8762 21666 8796
rect 21632 8694 21666 8728
rect 21632 8626 21666 8660
rect 21632 8558 21666 8592
rect 21632 8490 21666 8524
rect 21632 8422 21666 8456
rect 21632 8354 21666 8388
rect 21632 8286 21666 8320
rect 21632 8218 21666 8252
rect 21632 8150 21666 8184
rect 21632 8082 21666 8116
rect 21632 8014 21666 8048
rect 26398 8875 26432 8909
rect 26398 8807 26432 8841
rect 26398 8739 26432 8773
rect 26398 8671 26432 8705
rect 26398 8603 26432 8637
rect 26398 8535 26432 8569
rect 26398 8467 26432 8501
rect 26398 8399 26432 8433
rect 26398 8331 26432 8365
rect 26398 8263 26432 8297
rect 26398 8195 26432 8229
rect 26398 8127 26432 8161
rect 26398 8059 26432 8093
rect 21632 7946 21666 7980
rect 21632 7878 21666 7912
rect 21632 7810 21666 7844
rect 21632 7742 21666 7776
rect 21632 7674 21666 7708
rect 21632 7606 21666 7640
rect 21632 7538 21666 7572
rect 21632 7470 21666 7504
rect 21632 7402 21666 7436
rect 21632 7334 21666 7368
rect 21632 7266 21666 7300
rect 21632 7198 21666 7232
rect 21632 7130 21666 7164
rect 21632 7062 21666 7096
rect 21632 6994 21666 7028
rect 21632 6926 21666 6960
rect 21632 6858 21666 6892
rect 21632 6790 21666 6824
rect 21632 6722 21666 6756
rect 21632 6654 21666 6688
rect 21632 6586 21666 6620
rect 21632 6518 21666 6552
rect 21632 6450 21666 6484
rect 21632 6382 21666 6416
rect 21632 6314 21666 6348
rect 21632 6246 21666 6280
rect 21632 6178 21666 6212
rect 21632 6110 21666 6144
rect 21632 6042 21666 6076
rect 21632 5974 21666 6008
rect 21632 5906 21666 5940
rect 21632 5838 21666 5872
rect 21632 5770 21666 5804
rect 21632 5702 21666 5736
rect 21632 5634 21666 5668
rect 21632 5566 21666 5600
rect 21632 5498 21666 5532
rect 21632 5430 21666 5464
rect 21632 5362 21666 5396
rect 21632 5294 21666 5328
rect 21632 5226 21666 5260
rect 21632 5158 21666 5192
rect 21632 5090 21666 5124
rect 21632 5022 21666 5056
rect 21632 4954 21666 4988
rect 21632 4886 21666 4920
rect 21632 4818 21666 4852
rect 21632 4750 21666 4784
rect 20382 4624 20416 4716
rect 21632 4624 21666 4716
rect 20382 4590 20497 4624
rect 20531 4590 20565 4624
rect 20599 4590 20633 4624
rect 20667 4590 20701 4624
rect 20735 4590 20769 4624
rect 20803 4590 20837 4624
rect 20871 4590 20905 4624
rect 20939 4590 20973 4624
rect 21007 4590 21041 4624
rect 21075 4590 21109 4624
rect 21143 4590 21177 4624
rect 21211 4590 21245 4624
rect 21279 4590 21313 4624
rect 21347 4590 21381 4624
rect 21415 4590 21449 4624
rect 21483 4590 21517 4624
rect 21551 4590 21666 4624
rect 26398 7991 26432 8025
rect 26398 7923 26432 7957
rect 26398 7855 26432 7889
rect 26398 7787 26432 7821
rect 26398 7719 26432 7753
rect 26398 7651 26432 7685
rect 26398 7583 26432 7617
rect 26398 7515 26432 7549
rect 26398 7447 26432 7481
rect 26398 7379 26432 7413
rect 26398 7311 26432 7345
rect 26398 7243 26432 7277
rect 26398 7175 26432 7209
rect 26398 7107 26432 7141
rect 26398 7039 26432 7073
rect 26398 6971 26432 7005
rect 26398 6903 26432 6937
rect 26398 6835 26432 6869
rect 26398 6767 26432 6801
rect 26398 6699 26432 6733
rect 26398 6631 26432 6665
rect 26398 6563 26432 6597
rect 26398 6495 26432 6529
rect 26398 6427 26432 6461
rect 26398 6359 26432 6393
rect 26398 6291 26432 6325
rect 26398 6223 26432 6257
rect 26398 6155 26432 6189
rect 26398 6087 26432 6121
rect 26398 6019 26432 6053
rect 26398 5951 26432 5985
rect 26398 5883 26432 5917
rect 26398 5815 26432 5849
rect 26398 5747 26432 5781
rect 26398 5679 26432 5713
rect 26398 5611 26432 5645
rect 26398 5543 26432 5577
rect 26398 5475 26432 5509
rect 26398 5407 26432 5441
rect 26398 5339 26432 5373
rect 26398 5271 26432 5305
rect 26398 5203 26432 5237
rect 26398 5135 26432 5169
rect 26398 5067 26432 5101
rect 26398 4999 26432 5033
rect 26398 4931 26432 4965
rect 26398 4863 26432 4897
rect 26398 4795 26432 4829
rect 26398 4727 26432 4761
rect 26398 4659 26432 4693
rect 26398 4591 26432 4625
rect 26398 4523 26432 4557
rect 26398 4455 26432 4489
rect 26398 4387 26432 4421
rect 26398 4319 26432 4353
rect 26398 4251 26432 4285
rect 26398 4183 26432 4217
rect 26398 4115 26432 4149
rect 26398 4047 26432 4081
rect 26398 3979 26432 4013
rect 26398 3911 26432 3945
rect 26398 3843 26432 3877
rect 26398 3775 26432 3809
rect 26398 3707 26432 3741
rect 26398 3639 26432 3673
rect 26398 3571 26432 3605
rect 26398 3503 26432 3537
rect 26398 3435 26432 3469
rect 26398 3367 26432 3401
rect 26398 3299 26432 3333
rect 26398 3231 26432 3265
rect 26398 3163 26432 3197
rect 26398 3095 26432 3129
rect 27330 13295 27364 13329
rect 27330 13227 27364 13261
rect 27330 13159 27364 13193
rect 27330 13091 27364 13125
rect 27330 13023 27364 13057
rect 27330 12955 27364 12989
rect 27330 12887 27364 12921
rect 27330 12819 27364 12853
rect 27330 12751 27364 12785
rect 27330 12683 27364 12717
rect 27330 12615 27364 12649
rect 27330 12547 27364 12581
rect 27330 12479 27364 12513
rect 27330 12411 27364 12445
rect 27330 12343 27364 12377
rect 27330 12275 27364 12309
rect 27330 12207 27364 12241
rect 27330 12139 27364 12173
rect 27330 12071 27364 12105
rect 27330 12003 27364 12037
rect 27330 11935 27364 11969
rect 27330 11867 27364 11901
rect 27330 11799 27364 11833
rect 27330 11731 27364 11765
rect 27330 11663 27364 11697
rect 27330 11595 27364 11629
rect 27330 11527 27364 11561
rect 27330 11459 27364 11493
rect 27330 11391 27364 11425
rect 27330 11323 27364 11357
rect 27330 11255 27364 11289
rect 27330 11187 27364 11221
rect 27330 11119 27364 11153
rect 27330 11051 27364 11085
rect 27330 10983 27364 11017
rect 27330 10915 27364 10949
rect 27330 10847 27364 10881
rect 27330 10779 27364 10813
rect 27330 10711 27364 10745
rect 27330 10643 27364 10677
rect 27330 10575 27364 10609
rect 27330 10507 27364 10541
rect 27330 10439 27364 10473
rect 27330 10371 27364 10405
rect 27330 10303 27364 10337
rect 27330 10235 27364 10269
rect 27330 10167 27364 10201
rect 27330 10099 27364 10133
rect 27330 10031 27364 10065
rect 27330 9963 27364 9997
rect 27330 9895 27364 9929
rect 27330 9827 27364 9861
rect 27330 9759 27364 9793
rect 27330 9691 27364 9725
rect 27330 9623 27364 9657
rect 27330 9555 27364 9589
rect 27330 9487 27364 9521
rect 27330 9419 27364 9453
rect 27330 9351 27364 9385
rect 27330 9283 27364 9317
rect 27330 9215 27364 9249
rect 27330 9147 27364 9181
rect 27330 9079 27364 9113
rect 27330 9011 27364 9045
rect 27330 8943 27364 8977
rect 27330 8875 27364 8909
rect 27330 8807 27364 8841
rect 27330 8739 27364 8773
rect 27330 8671 27364 8705
rect 27330 8603 27364 8637
rect 27330 8535 27364 8569
rect 27330 8467 27364 8501
rect 27330 8399 27364 8433
rect 27330 8331 27364 8365
rect 27330 8263 27364 8297
rect 27330 8195 27364 8229
rect 27330 8127 27364 8161
rect 27330 8059 27364 8093
rect 27330 7991 27364 8025
rect 27330 7923 27364 7957
rect 27330 7855 27364 7889
rect 27330 7787 27364 7821
rect 27330 7719 27364 7753
rect 27330 7651 27364 7685
rect 27330 7583 27364 7617
rect 27330 7515 27364 7549
rect 27330 7447 27364 7481
rect 27330 7379 27364 7413
rect 27330 7311 27364 7345
rect 27330 7243 27364 7277
rect 27330 7175 27364 7209
rect 27330 7107 27364 7141
rect 27330 7039 27364 7073
rect 27330 6971 27364 7005
rect 27330 6903 27364 6937
rect 27330 6835 27364 6869
rect 27330 6767 27364 6801
rect 27330 6699 27364 6733
rect 27330 6631 27364 6665
rect 27330 6563 27364 6597
rect 27330 6495 27364 6529
rect 27330 6427 27364 6461
rect 27330 6359 27364 6393
rect 27570 13424 27686 13458
rect 27720 13424 27754 13458
rect 27788 13424 27822 13458
rect 27856 13424 27890 13458
rect 27924 13424 27958 13458
rect 27992 13424 28026 13458
rect 28060 13424 28094 13458
rect 28128 13424 28162 13458
rect 28196 13424 28230 13458
rect 28264 13424 28298 13458
rect 28332 13424 28366 13458
rect 28400 13424 28434 13458
rect 28468 13424 28502 13458
rect 28536 13424 28570 13458
rect 28604 13424 28638 13458
rect 28672 13424 28706 13458
rect 28740 13424 28774 13458
rect 28808 13424 28842 13458
rect 28876 13424 28910 13458
rect 28944 13424 28978 13458
rect 29012 13424 29046 13458
rect 29080 13424 29114 13458
rect 29148 13424 29182 13458
rect 29216 13424 29250 13458
rect 29284 13424 29318 13458
rect 29352 13424 29386 13458
rect 29420 13424 29454 13458
rect 29488 13424 29522 13458
rect 29556 13424 29590 13458
rect 29624 13424 29658 13458
rect 29692 13424 29808 13458
rect 27570 13347 27604 13424
rect 29774 13347 29808 13424
rect 27570 13279 27604 13313
rect 27570 13211 27604 13245
rect 27570 13143 27604 13177
rect 27570 13075 27604 13109
rect 27570 13007 27604 13041
rect 27570 12939 27604 12973
rect 27570 12871 27604 12905
rect 27570 12803 27604 12837
rect 27570 12735 27604 12769
rect 27570 12667 27604 12701
rect 27570 12599 27604 12633
rect 27570 12531 27604 12565
rect 27570 12463 27604 12497
rect 27570 12395 27604 12429
rect 27570 12327 27604 12361
rect 27570 12259 27604 12293
rect 27570 12191 27604 12225
rect 27570 12123 27604 12157
rect 27570 12055 27604 12089
rect 27570 11987 27604 12021
rect 27570 11919 27604 11953
rect 27570 11851 27604 11885
rect 27570 11783 27604 11817
rect 27570 11715 27604 11749
rect 27570 11647 27604 11681
rect 27570 11579 27604 11613
rect 27570 11511 27604 11545
rect 27570 11443 27604 11477
rect 27570 11375 27604 11409
rect 27570 11307 27604 11341
rect 27570 11239 27604 11273
rect 27570 11171 27604 11205
rect 27570 11103 27604 11137
rect 27570 11035 27604 11069
rect 27570 10967 27604 11001
rect 27570 10899 27604 10933
rect 27570 10831 27604 10865
rect 27570 10763 27604 10797
rect 27570 10695 27604 10729
rect 27570 10627 27604 10661
rect 27570 10559 27604 10593
rect 27570 10491 27604 10525
rect 27570 10423 27604 10457
rect 27570 10355 27604 10389
rect 27570 10287 27604 10321
rect 27570 10219 27604 10253
rect 27570 10151 27604 10185
rect 27570 10083 27604 10117
rect 27570 10015 27604 10049
rect 27570 9947 27604 9981
rect 27570 9879 27604 9913
rect 27570 9811 27604 9845
rect 27570 9743 27604 9777
rect 27570 9675 27604 9709
rect 27570 9607 27604 9641
rect 27570 9539 27604 9573
rect 27570 9471 27604 9505
rect 27570 9403 27604 9437
rect 27570 9335 27604 9369
rect 27570 9267 27604 9301
rect 27570 9199 27604 9233
rect 27570 9131 27604 9165
rect 27570 9063 27604 9097
rect 27570 8995 27604 9029
rect 27570 8927 27604 8961
rect 27570 8859 27604 8893
rect 27570 8791 27604 8825
rect 27570 8723 27604 8757
rect 27570 8655 27604 8689
rect 27570 8587 27604 8621
rect 27570 8519 27604 8553
rect 27570 8451 27604 8485
rect 27570 8383 27604 8417
rect 27570 8315 27604 8349
rect 27570 8247 27604 8281
rect 27570 8179 27604 8213
rect 27570 8111 27604 8145
rect 27570 8043 27604 8077
rect 27570 7975 27604 8009
rect 27570 7907 27604 7941
rect 27570 7839 27604 7873
rect 27570 7771 27604 7805
rect 27570 7703 27604 7737
rect 27570 7635 27604 7669
rect 27570 7567 27604 7601
rect 27570 7499 27604 7533
rect 27570 7431 27604 7465
rect 27570 7363 27604 7397
rect 27570 7295 27604 7329
rect 27570 7227 27604 7261
rect 27570 7159 27604 7193
rect 27570 7091 27604 7125
rect 27570 7023 27604 7057
rect 27570 6955 27604 6989
rect 27570 6887 27604 6921
rect 27570 6819 27604 6853
rect 27570 6751 27604 6785
rect 27570 6683 27604 6717
rect 27570 6615 27604 6649
rect 27570 6547 27604 6581
rect 27570 6479 27604 6513
rect 29774 13279 29808 13313
rect 29774 13211 29808 13245
rect 29774 13143 29808 13177
rect 29774 13075 29808 13109
rect 29774 13007 29808 13041
rect 29774 12939 29808 12973
rect 29774 12871 29808 12905
rect 37706 13440 37749 13474
rect 37783 13440 37839 13474
rect 37706 13406 37839 13440
rect 37706 13372 37749 13406
rect 37783 13372 37839 13406
rect 41047 13536 41089 13570
rect 41123 13536 41165 13570
rect 41047 13502 41165 13536
rect 41047 13468 41089 13502
rect 41123 13468 41165 13502
rect 41047 13434 41165 13468
rect 41047 13400 41089 13434
rect 41123 13400 41165 13434
rect 37706 13338 37839 13372
rect 37706 13304 37749 13338
rect 37783 13304 37839 13338
rect 37706 13270 37839 13304
rect 37706 13236 37749 13270
rect 37783 13236 37839 13270
rect 37706 13202 37839 13236
rect 37706 13168 37749 13202
rect 37783 13168 37839 13202
rect 37706 13134 37839 13168
rect 37706 13100 37749 13134
rect 37783 13100 37839 13134
rect 37706 13026 37839 13100
rect 41047 13366 41165 13400
rect 41047 13332 41089 13366
rect 41123 13332 41165 13366
rect 41047 13298 41165 13332
rect 41047 13264 41089 13298
rect 41123 13264 41165 13298
rect 41047 13230 41165 13264
rect 41047 13196 41089 13230
rect 41123 13196 41165 13230
rect 41047 13162 41165 13196
rect 41047 13128 41089 13162
rect 41123 13128 41165 13162
rect 41047 13094 41165 13128
rect 41047 13060 41089 13094
rect 41123 13060 41165 13094
rect 41582 15751 41696 15785
rect 41730 15751 41764 15785
rect 41798 15751 41912 15785
rect 41582 15664 41616 15751
rect 41878 15664 41912 15751
rect 41582 15596 41616 15630
rect 41582 15528 41616 15562
rect 41582 15460 41616 15494
rect 41582 15392 41616 15426
rect 41582 15324 41616 15358
rect 41582 15256 41616 15290
rect 41582 15188 41616 15222
rect 41582 15120 41616 15154
rect 41582 15052 41616 15086
rect 41582 14984 41616 15018
rect 41582 14916 41616 14950
rect 41582 14848 41616 14882
rect 41582 14780 41616 14814
rect 41582 14712 41616 14746
rect 41582 14644 41616 14678
rect 41582 14576 41616 14610
rect 41582 14508 41616 14542
rect 41582 14440 41616 14474
rect 41582 14372 41616 14406
rect 41582 14304 41616 14338
rect 41582 14236 41616 14270
rect 41582 14168 41616 14202
rect 41582 14100 41616 14134
rect 41582 14032 41616 14066
rect 41582 13964 41616 13998
rect 41582 13896 41616 13930
rect 41582 13828 41616 13862
rect 41582 13760 41616 13794
rect 41582 13692 41616 13726
rect 41582 13624 41616 13658
rect 41582 13556 41616 13590
rect 41582 13488 41616 13522
rect 41582 13420 41616 13454
rect 41582 13352 41616 13386
rect 41582 13284 41616 13318
rect 41582 13216 41616 13250
rect 41878 15596 41912 15630
rect 41878 15528 41912 15562
rect 41878 15460 41912 15494
rect 41878 15392 41912 15426
rect 41878 15324 41912 15358
rect 41878 15256 41912 15290
rect 41878 15188 41912 15222
rect 41878 15120 41912 15154
rect 41878 15052 41912 15086
rect 41878 14984 41912 15018
rect 41878 14916 41912 14950
rect 41878 14848 41912 14882
rect 41878 14780 41912 14814
rect 41878 14712 41912 14746
rect 41878 14644 41912 14678
rect 41878 14576 41912 14610
rect 41878 14508 41912 14542
rect 41878 14440 41912 14474
rect 41878 14372 41912 14406
rect 41878 14304 41912 14338
rect 41878 14236 41912 14270
rect 41878 14168 41912 14202
rect 41878 14100 41912 14134
rect 41878 14032 41912 14066
rect 41878 13964 41912 13998
rect 41878 13896 41912 13930
rect 41878 13828 41912 13862
rect 41878 13760 41912 13794
rect 41878 13692 41912 13726
rect 41878 13624 41912 13658
rect 41878 13556 41912 13590
rect 41878 13488 41912 13522
rect 41878 13420 41912 13454
rect 41878 13352 41912 13386
rect 41878 13284 41912 13318
rect 41878 13216 41912 13250
rect 41582 13095 41616 13182
rect 41878 13095 41912 13182
rect 41582 13061 41696 13095
rect 41730 13061 41764 13095
rect 41798 13061 41912 13095
rect 41047 13026 41165 13060
rect 37706 12986 41165 13026
rect 37706 12952 38022 12986
rect 38056 12952 38090 12986
rect 38124 12952 38158 12986
rect 38192 12952 38226 12986
rect 38260 12952 38294 12986
rect 38328 12952 38362 12986
rect 38396 12952 38430 12986
rect 38464 12952 38498 12986
rect 38532 12952 38566 12986
rect 38600 12952 38634 12986
rect 38668 12952 38702 12986
rect 38736 12952 38770 12986
rect 38804 12952 38838 12986
rect 38872 12952 38906 12986
rect 38940 12952 38974 12986
rect 39008 12952 39042 12986
rect 39076 12952 39110 12986
rect 39144 12952 39178 12986
rect 39212 12952 39246 12986
rect 39280 12952 39314 12986
rect 39348 12952 39382 12986
rect 39416 12952 39450 12986
rect 39484 12952 39518 12986
rect 39552 12952 39586 12986
rect 39620 12952 39654 12986
rect 39688 12952 39722 12986
rect 39756 12952 39790 12986
rect 39824 12952 39858 12986
rect 39892 12952 39926 12986
rect 39960 12952 39994 12986
rect 40028 12952 40062 12986
rect 40096 12952 40130 12986
rect 40164 12952 40198 12986
rect 40232 12952 40266 12986
rect 40300 12952 40334 12986
rect 40368 12952 40402 12986
rect 40436 12952 40470 12986
rect 40504 12952 40538 12986
rect 40572 12952 40606 12986
rect 40640 12952 40674 12986
rect 40708 12952 40742 12986
rect 40776 12952 40810 12986
rect 40844 12952 40878 12986
rect 40912 12952 40946 12986
rect 40980 12952 41165 12986
rect 37706 12884 41165 12952
rect 29774 12803 29808 12837
rect 29774 12735 29808 12769
rect 29774 12667 29808 12701
rect 29774 12599 29808 12633
rect 29774 12531 29808 12565
rect 29774 12463 29808 12497
rect 29774 12395 29808 12429
rect 29774 12327 29808 12361
rect 29774 12259 29808 12293
rect 29774 12191 29808 12225
rect 29774 12123 29808 12157
rect 29774 12055 29808 12089
rect 29774 11987 29808 12021
rect 29774 11919 29808 11953
rect 29774 11851 29808 11885
rect 29774 11783 29808 11817
rect 29774 11715 29808 11749
rect 29774 11647 29808 11681
rect 29774 11579 29808 11613
rect 29774 11511 29808 11545
rect 29774 11443 29808 11477
rect 29774 11375 29808 11409
rect 29774 11307 29808 11341
rect 29774 11239 29808 11273
rect 29774 11171 29808 11205
rect 29774 11103 29808 11137
rect 29774 11035 29808 11069
rect 29774 10967 29808 11001
rect 29774 10899 29808 10933
rect 29774 10831 29808 10865
rect 29774 10763 29808 10797
rect 29774 10695 29808 10729
rect 29774 10627 29808 10661
rect 29774 10559 29808 10593
rect 29774 10491 29808 10525
rect 29774 10423 29808 10457
rect 29774 10355 29808 10389
rect 29774 10287 29808 10321
rect 29774 10219 29808 10253
rect 29774 10151 29808 10185
rect 29774 10083 29808 10117
rect 29774 10015 29808 10049
rect 29774 9947 29808 9981
rect 29774 9879 29808 9913
rect 29774 9811 29808 9845
rect 29774 9743 29808 9777
rect 29774 9675 29808 9709
rect 29774 9607 29808 9641
rect 29774 9539 29808 9573
rect 29774 9471 29808 9505
rect 29774 9403 29808 9437
rect 29774 9335 29808 9369
rect 29774 9267 29808 9301
rect 29774 9199 29808 9233
rect 29774 9131 29808 9165
rect 29774 9063 29808 9097
rect 29774 8995 29808 9029
rect 29774 8927 29808 8961
rect 29774 8859 29808 8893
rect 29774 8791 29808 8825
rect 29774 8723 29808 8757
rect 29774 8655 29808 8689
rect 29774 8587 29808 8621
rect 29774 8519 29808 8553
rect 29774 8451 29808 8485
rect 29774 8383 29808 8417
rect 29774 8315 29808 8349
rect 29774 8247 29808 8281
rect 29774 8179 29808 8213
rect 29774 8111 29808 8145
rect 29774 8043 29808 8077
rect 29774 7975 29808 8009
rect 29774 7907 29808 7941
rect 29774 7839 29808 7873
rect 29774 7771 29808 7805
rect 29774 7703 29808 7737
rect 29774 7635 29808 7669
rect 29774 7567 29808 7601
rect 29774 7499 29808 7533
rect 29774 7431 29808 7465
rect 29774 7363 29808 7397
rect 29774 7295 29808 7329
rect 29774 7227 29808 7261
rect 29774 7159 29808 7193
rect 29774 7091 29808 7125
rect 29774 7023 29808 7057
rect 29774 6955 29808 6989
rect 29774 6887 29808 6921
rect 29774 6819 29808 6853
rect 29774 6751 29808 6785
rect 29774 6683 29808 6717
rect 29774 6615 29808 6649
rect 29774 6547 29808 6581
rect 29774 6479 29808 6513
rect 27570 6368 27604 6445
rect 29774 6368 29808 6445
rect 27570 6334 27686 6368
rect 27720 6334 27754 6368
rect 27788 6334 27822 6368
rect 27856 6334 27890 6368
rect 27924 6334 27958 6368
rect 27992 6334 28026 6368
rect 28060 6334 28094 6368
rect 28128 6334 28162 6368
rect 28196 6334 28230 6368
rect 28264 6334 28298 6368
rect 28332 6334 28366 6368
rect 28400 6334 28434 6368
rect 28468 6334 28502 6368
rect 28536 6334 28570 6368
rect 28604 6334 28638 6368
rect 28672 6334 28706 6368
rect 28740 6334 28774 6368
rect 28808 6334 28842 6368
rect 28876 6334 28910 6368
rect 28944 6334 28978 6368
rect 29012 6334 29046 6368
rect 29080 6334 29114 6368
rect 29148 6334 29182 6368
rect 29216 6334 29250 6368
rect 29284 6334 29318 6368
rect 29352 6334 29386 6368
rect 29420 6334 29454 6368
rect 29488 6334 29522 6368
rect 29556 6334 29590 6368
rect 29624 6334 29658 6368
rect 29692 6334 29808 6368
rect 27330 6291 27364 6325
rect 27330 6223 27364 6257
rect 27330 6155 27364 6189
rect 27330 6087 27364 6121
rect 27330 6019 27364 6053
rect 27330 5951 27364 5985
rect 27330 5883 27364 5917
rect 27330 5815 27364 5849
rect 27330 5747 27364 5781
rect 27330 5679 27364 5713
rect 27330 5611 27364 5645
rect 27330 5543 27364 5577
rect 27330 5475 27364 5509
rect 27330 5407 27364 5441
rect 27330 5339 27364 5373
rect 27330 5271 27364 5305
rect 27330 5203 27364 5237
rect 27330 5135 27364 5169
rect 27330 5067 27364 5101
rect 27330 4999 27364 5033
rect 27330 4931 27364 4965
rect 27330 4863 27364 4897
rect 27330 4795 27364 4829
rect 27330 4727 27364 4761
rect 27330 4659 27364 4693
rect 27330 4591 27364 4625
rect 27330 4523 27364 4557
rect 27330 4455 27364 4489
rect 27330 4387 27364 4421
rect 27330 4319 27364 4353
rect 27330 4251 27364 4285
rect 27330 4183 27364 4217
rect 27330 4115 27364 4149
rect 27330 4047 27364 4081
rect 27330 3979 27364 4013
rect 27330 3911 27364 3945
rect 27330 3843 27364 3877
rect 27330 3775 27364 3809
rect 27330 3707 27364 3741
rect 27330 3639 27364 3673
rect 27330 3571 27364 3605
rect 27330 3503 27364 3537
rect 27330 3435 27364 3469
rect 27330 3367 27364 3401
rect 27330 3299 27364 3333
rect 27330 3231 27364 3265
rect 27330 3163 27364 3197
rect 27330 3095 27364 3129
rect 26398 2984 26432 3061
rect 27330 2984 27364 3061
rect 26398 2950 26524 2984
rect 26558 2950 26592 2984
rect 26626 2950 26660 2984
rect 26694 2950 26728 2984
rect 26762 2950 26796 2984
rect 26830 2950 26864 2984
rect 26898 2950 26932 2984
rect 26966 2950 27000 2984
rect 27034 2950 27068 2984
rect 27102 2950 27136 2984
rect 27170 2950 27204 2984
rect 27238 2950 27364 2984
<< nsubdiff >>
rect 23273 15670 24235 15689
rect 23273 15636 23404 15670
rect 23438 15636 23494 15670
rect 23528 15636 23584 15670
rect 23618 15636 23674 15670
rect 23708 15636 23764 15670
rect 23798 15636 23854 15670
rect 23888 15636 23944 15670
rect 23978 15636 24034 15670
rect 24068 15636 24124 15670
rect 24158 15636 24235 15670
rect 23273 15617 24235 15636
rect 23273 15613 23345 15617
rect 23273 15579 23292 15613
rect 23326 15579 23345 15613
rect 23273 15523 23345 15579
rect 24163 15594 24235 15617
rect 24163 15560 24182 15594
rect 24216 15560 24235 15594
rect 23273 15489 23292 15523
rect 23326 15489 23345 15523
rect 23273 15433 23345 15489
rect 23273 15399 23292 15433
rect 23326 15399 23345 15433
rect 23273 15343 23345 15399
rect 23273 15309 23292 15343
rect 23326 15309 23345 15343
rect 23273 15253 23345 15309
rect 23273 15219 23292 15253
rect 23326 15219 23345 15253
rect 23273 15163 23345 15219
rect 23273 15129 23292 15163
rect 23326 15129 23345 15163
rect 23273 15073 23345 15129
rect 23273 15039 23292 15073
rect 23326 15039 23345 15073
rect 23273 14983 23345 15039
rect 23273 14949 23292 14983
rect 23326 14949 23345 14983
rect 23273 14893 23345 14949
rect 23273 14859 23292 14893
rect 23326 14859 23345 14893
rect 24163 15504 24235 15560
rect 24163 15470 24182 15504
rect 24216 15470 24235 15504
rect 24163 15414 24235 15470
rect 24163 15380 24182 15414
rect 24216 15380 24235 15414
rect 24163 15324 24235 15380
rect 24163 15290 24182 15324
rect 24216 15290 24235 15324
rect 24163 15234 24235 15290
rect 24163 15200 24182 15234
rect 24216 15200 24235 15234
rect 24163 15144 24235 15200
rect 24163 15110 24182 15144
rect 24216 15110 24235 15144
rect 24163 15054 24235 15110
rect 24163 15020 24182 15054
rect 24216 15020 24235 15054
rect 24163 14964 24235 15020
rect 24163 14930 24182 14964
rect 24216 14930 24235 14964
rect 24163 14874 24235 14930
rect 23273 14799 23345 14859
rect 24163 14840 24182 14874
rect 24216 14840 24235 14874
rect 24163 14799 24235 14840
rect 23273 14780 24235 14799
rect 23273 14746 23370 14780
rect 23404 14746 23460 14780
rect 23494 14746 23550 14780
rect 23584 14746 23640 14780
rect 23674 14746 23730 14780
rect 23764 14746 23820 14780
rect 23854 14746 23910 14780
rect 23944 14746 24000 14780
rect 24034 14746 24090 14780
rect 24124 14746 24235 14780
rect 23273 14727 24235 14746
rect 12945 11152 13907 11171
rect 12945 11118 13076 11152
rect 13110 11118 13166 11152
rect 13200 11118 13256 11152
rect 13290 11118 13346 11152
rect 13380 11118 13436 11152
rect 13470 11118 13526 11152
rect 13560 11118 13616 11152
rect 13650 11118 13706 11152
rect 13740 11118 13796 11152
rect 13830 11118 13907 11152
rect 12945 11099 13907 11118
rect 12945 11095 13017 11099
rect 12945 11061 12964 11095
rect 12998 11061 13017 11095
rect 12945 11005 13017 11061
rect 13835 11076 13907 11099
rect 13835 11042 13854 11076
rect 13888 11042 13907 11076
rect 12945 10971 12964 11005
rect 12998 10971 13017 11005
rect 12945 10915 13017 10971
rect 12945 10881 12964 10915
rect 12998 10881 13017 10915
rect 12945 10825 13017 10881
rect 12945 10791 12964 10825
rect 12998 10791 13017 10825
rect 12945 10735 13017 10791
rect 12945 10701 12964 10735
rect 12998 10701 13017 10735
rect 12945 10645 13017 10701
rect 12945 10611 12964 10645
rect 12998 10611 13017 10645
rect 12945 10555 13017 10611
rect 12945 10521 12964 10555
rect 12998 10521 13017 10555
rect 12945 10465 13017 10521
rect 12945 10431 12964 10465
rect 12998 10431 13017 10465
rect 12945 10375 13017 10431
rect 12945 10341 12964 10375
rect 12998 10341 13017 10375
rect 13835 10986 13907 11042
rect 13835 10952 13854 10986
rect 13888 10952 13907 10986
rect 13835 10896 13907 10952
rect 13835 10862 13854 10896
rect 13888 10862 13907 10896
rect 13835 10806 13907 10862
rect 13835 10772 13854 10806
rect 13888 10772 13907 10806
rect 13835 10716 13907 10772
rect 13835 10682 13854 10716
rect 13888 10682 13907 10716
rect 13835 10626 13907 10682
rect 13835 10592 13854 10626
rect 13888 10592 13907 10626
rect 13835 10536 13907 10592
rect 13835 10502 13854 10536
rect 13888 10502 13907 10536
rect 13835 10446 13907 10502
rect 13835 10412 13854 10446
rect 13888 10412 13907 10446
rect 13835 10356 13907 10412
rect 12945 10281 13017 10341
rect 13835 10322 13854 10356
rect 13888 10322 13907 10356
rect 13835 10281 13907 10322
rect 12945 10262 13907 10281
rect 12945 10228 13042 10262
rect 13076 10228 13132 10262
rect 13166 10228 13222 10262
rect 13256 10228 13312 10262
rect 13346 10228 13402 10262
rect 13436 10228 13492 10262
rect 13526 10228 13582 10262
rect 13616 10228 13672 10262
rect 13706 10228 13762 10262
rect 13796 10228 13907 10262
rect 12945 10209 13907 10228
rect 12945 9662 13907 9681
rect 12945 9628 13076 9662
rect 13110 9628 13166 9662
rect 13200 9628 13256 9662
rect 13290 9628 13346 9662
rect 13380 9628 13436 9662
rect 13470 9628 13526 9662
rect 13560 9628 13616 9662
rect 13650 9628 13706 9662
rect 13740 9628 13796 9662
rect 13830 9628 13907 9662
rect 12945 9609 13907 9628
rect 12945 9605 13017 9609
rect 12945 9571 12964 9605
rect 12998 9571 13017 9605
rect 12945 9515 13017 9571
rect 13835 9586 13907 9609
rect 13835 9552 13854 9586
rect 13888 9552 13907 9586
rect 12945 9481 12964 9515
rect 12998 9481 13017 9515
rect 12945 9425 13017 9481
rect 12945 9391 12964 9425
rect 12998 9391 13017 9425
rect 12945 9335 13017 9391
rect 12945 9301 12964 9335
rect 12998 9301 13017 9335
rect 12945 9245 13017 9301
rect 12945 9211 12964 9245
rect 12998 9211 13017 9245
rect 12945 9155 13017 9211
rect 12945 9121 12964 9155
rect 12998 9121 13017 9155
rect 12945 9065 13017 9121
rect 12945 9031 12964 9065
rect 12998 9031 13017 9065
rect 12945 8975 13017 9031
rect 12945 8941 12964 8975
rect 12998 8941 13017 8975
rect 12945 8885 13017 8941
rect 12945 8851 12964 8885
rect 12998 8851 13017 8885
rect 13835 9496 13907 9552
rect 13835 9462 13854 9496
rect 13888 9462 13907 9496
rect 13835 9406 13907 9462
rect 13835 9372 13854 9406
rect 13888 9372 13907 9406
rect 13835 9316 13907 9372
rect 13835 9282 13854 9316
rect 13888 9282 13907 9316
rect 13835 9226 13907 9282
rect 13835 9192 13854 9226
rect 13888 9192 13907 9226
rect 13835 9136 13907 9192
rect 13835 9102 13854 9136
rect 13888 9102 13907 9136
rect 13835 9046 13907 9102
rect 13835 9012 13854 9046
rect 13888 9012 13907 9046
rect 13835 8956 13907 9012
rect 13835 8922 13854 8956
rect 13888 8922 13907 8956
rect 13835 8866 13907 8922
rect 12945 8791 13017 8851
rect 13835 8832 13854 8866
rect 13888 8832 13907 8866
rect 13835 8791 13907 8832
rect 12945 8772 13907 8791
rect 12945 8738 13042 8772
rect 13076 8738 13132 8772
rect 13166 8738 13222 8772
rect 13256 8738 13312 8772
rect 13346 8738 13402 8772
rect 13436 8738 13492 8772
rect 13526 8738 13582 8772
rect 13616 8738 13672 8772
rect 13706 8738 13762 8772
rect 13796 8738 13907 8772
rect 12945 8719 13907 8738
rect 12935 8252 13897 8271
rect 12935 8218 13066 8252
rect 13100 8218 13156 8252
rect 13190 8218 13246 8252
rect 13280 8218 13336 8252
rect 13370 8218 13426 8252
rect 13460 8218 13516 8252
rect 13550 8218 13606 8252
rect 13640 8218 13696 8252
rect 13730 8218 13786 8252
rect 13820 8218 13897 8252
rect 12935 8199 13897 8218
rect 12935 8195 13007 8199
rect 12935 8161 12954 8195
rect 12988 8161 13007 8195
rect 12935 8105 13007 8161
rect 13825 8176 13897 8199
rect 13825 8142 13844 8176
rect 13878 8142 13897 8176
rect 12935 8071 12954 8105
rect 12988 8071 13007 8105
rect 12935 8015 13007 8071
rect 12935 7981 12954 8015
rect 12988 7981 13007 8015
rect 12935 7925 13007 7981
rect 12935 7891 12954 7925
rect 12988 7891 13007 7925
rect 12935 7835 13007 7891
rect 12935 7801 12954 7835
rect 12988 7801 13007 7835
rect 12935 7745 13007 7801
rect 12935 7711 12954 7745
rect 12988 7711 13007 7745
rect 12935 7655 13007 7711
rect 12935 7621 12954 7655
rect 12988 7621 13007 7655
rect 12935 7565 13007 7621
rect 12935 7531 12954 7565
rect 12988 7531 13007 7565
rect 12935 7475 13007 7531
rect 12935 7441 12954 7475
rect 12988 7441 13007 7475
rect 13825 8086 13897 8142
rect 13825 8052 13844 8086
rect 13878 8052 13897 8086
rect 13825 7996 13897 8052
rect 13825 7962 13844 7996
rect 13878 7962 13897 7996
rect 13825 7906 13897 7962
rect 13825 7872 13844 7906
rect 13878 7872 13897 7906
rect 13825 7816 13897 7872
rect 13825 7782 13844 7816
rect 13878 7782 13897 7816
rect 13825 7726 13897 7782
rect 13825 7692 13844 7726
rect 13878 7692 13897 7726
rect 13825 7636 13897 7692
rect 13825 7602 13844 7636
rect 13878 7602 13897 7636
rect 13825 7546 13897 7602
rect 13825 7512 13844 7546
rect 13878 7512 13897 7546
rect 13825 7456 13897 7512
rect 12935 7381 13007 7441
rect 13825 7422 13844 7456
rect 13878 7422 13897 7456
rect 13825 7381 13897 7422
rect 12935 7362 13897 7381
rect 12935 7328 13032 7362
rect 13066 7328 13122 7362
rect 13156 7328 13212 7362
rect 13246 7328 13302 7362
rect 13336 7328 13392 7362
rect 13426 7328 13482 7362
rect 13516 7328 13572 7362
rect 13606 7328 13662 7362
rect 13696 7328 13752 7362
rect 13786 7328 13897 7362
rect 12935 7309 13897 7328
rect 12935 6902 13897 6921
rect 12935 6868 13066 6902
rect 13100 6868 13156 6902
rect 13190 6868 13246 6902
rect 13280 6868 13336 6902
rect 13370 6868 13426 6902
rect 13460 6868 13516 6902
rect 13550 6868 13606 6902
rect 13640 6868 13696 6902
rect 13730 6868 13786 6902
rect 13820 6868 13897 6902
rect 12935 6849 13897 6868
rect 12935 6845 13007 6849
rect 12935 6811 12954 6845
rect 12988 6811 13007 6845
rect 12935 6755 13007 6811
rect 13825 6826 13897 6849
rect 13825 6792 13844 6826
rect 13878 6792 13897 6826
rect 12935 6721 12954 6755
rect 12988 6721 13007 6755
rect 12935 6665 13007 6721
rect 12935 6631 12954 6665
rect 12988 6631 13007 6665
rect 12935 6575 13007 6631
rect 12935 6541 12954 6575
rect 12988 6541 13007 6575
rect 12935 6485 13007 6541
rect 12935 6451 12954 6485
rect 12988 6451 13007 6485
rect 12935 6395 13007 6451
rect 12935 6361 12954 6395
rect 12988 6361 13007 6395
rect 12935 6305 13007 6361
rect 12935 6271 12954 6305
rect 12988 6271 13007 6305
rect 12935 6215 13007 6271
rect 12935 6181 12954 6215
rect 12988 6181 13007 6215
rect 12935 6125 13007 6181
rect 12935 6091 12954 6125
rect 12988 6091 13007 6125
rect 13825 6736 13897 6792
rect 13825 6702 13844 6736
rect 13878 6702 13897 6736
rect 13825 6646 13897 6702
rect 13825 6612 13844 6646
rect 13878 6612 13897 6646
rect 13825 6556 13897 6612
rect 13825 6522 13844 6556
rect 13878 6522 13897 6556
rect 13825 6466 13897 6522
rect 13825 6432 13844 6466
rect 13878 6432 13897 6466
rect 13825 6376 13897 6432
rect 13825 6342 13844 6376
rect 13878 6342 13897 6376
rect 13825 6286 13897 6342
rect 13825 6252 13844 6286
rect 13878 6252 13897 6286
rect 13825 6196 13897 6252
rect 13825 6162 13844 6196
rect 13878 6162 13897 6196
rect 13825 6106 13897 6162
rect 12935 6031 13007 6091
rect 13825 6072 13844 6106
rect 13878 6072 13897 6106
rect 13825 6031 13897 6072
rect 12935 6012 13897 6031
rect 12935 5978 13032 6012
rect 13066 5978 13122 6012
rect 13156 5978 13212 6012
rect 13246 5978 13302 6012
rect 13336 5978 13392 6012
rect 13426 5978 13482 6012
rect 13516 5978 13572 6012
rect 13606 5978 13662 6012
rect 13696 5978 13752 6012
rect 13786 5978 13897 6012
rect 12935 5959 13897 5978
rect 14585 6932 15547 6951
rect 14585 6898 14716 6932
rect 14750 6898 14806 6932
rect 14840 6898 14896 6932
rect 14930 6898 14986 6932
rect 15020 6898 15076 6932
rect 15110 6898 15166 6932
rect 15200 6898 15256 6932
rect 15290 6898 15346 6932
rect 15380 6898 15436 6932
rect 15470 6898 15547 6932
rect 14585 6879 15547 6898
rect 14585 6875 14657 6879
rect 14585 6841 14604 6875
rect 14638 6841 14657 6875
rect 14585 6785 14657 6841
rect 15475 6856 15547 6879
rect 15475 6822 15494 6856
rect 15528 6822 15547 6856
rect 14585 6751 14604 6785
rect 14638 6751 14657 6785
rect 14585 6695 14657 6751
rect 14585 6661 14604 6695
rect 14638 6661 14657 6695
rect 14585 6605 14657 6661
rect 14585 6571 14604 6605
rect 14638 6571 14657 6605
rect 14585 6515 14657 6571
rect 14585 6481 14604 6515
rect 14638 6481 14657 6515
rect 14585 6425 14657 6481
rect 14585 6391 14604 6425
rect 14638 6391 14657 6425
rect 14585 6335 14657 6391
rect 14585 6301 14604 6335
rect 14638 6301 14657 6335
rect 14585 6245 14657 6301
rect 14585 6211 14604 6245
rect 14638 6211 14657 6245
rect 14585 6155 14657 6211
rect 14585 6121 14604 6155
rect 14638 6121 14657 6155
rect 15475 6766 15547 6822
rect 15475 6732 15494 6766
rect 15528 6732 15547 6766
rect 15475 6676 15547 6732
rect 15475 6642 15494 6676
rect 15528 6642 15547 6676
rect 15475 6586 15547 6642
rect 15475 6552 15494 6586
rect 15528 6552 15547 6586
rect 15475 6496 15547 6552
rect 15475 6462 15494 6496
rect 15528 6462 15547 6496
rect 15475 6406 15547 6462
rect 15475 6372 15494 6406
rect 15528 6372 15547 6406
rect 15475 6316 15547 6372
rect 15475 6282 15494 6316
rect 15528 6282 15547 6316
rect 15475 6226 15547 6282
rect 15475 6192 15494 6226
rect 15528 6192 15547 6226
rect 15475 6136 15547 6192
rect 14585 6061 14657 6121
rect 15475 6102 15494 6136
rect 15528 6102 15547 6136
rect 15475 6061 15547 6102
rect 14585 6042 15547 6061
rect 14585 6008 14682 6042
rect 14716 6008 14772 6042
rect 14806 6008 14862 6042
rect 14896 6008 14952 6042
rect 14986 6008 15042 6042
rect 15076 6008 15132 6042
rect 15166 6008 15222 6042
rect 15256 6008 15312 6042
rect 15346 6008 15402 6042
rect 15436 6008 15547 6042
rect 14585 5989 15547 6008
rect 12935 5552 13897 5571
rect 12935 5518 13066 5552
rect 13100 5518 13156 5552
rect 13190 5518 13246 5552
rect 13280 5518 13336 5552
rect 13370 5518 13426 5552
rect 13460 5518 13516 5552
rect 13550 5518 13606 5552
rect 13640 5518 13696 5552
rect 13730 5518 13786 5552
rect 13820 5518 13897 5552
rect 12935 5499 13897 5518
rect 12935 5495 13007 5499
rect 12935 5461 12954 5495
rect 12988 5461 13007 5495
rect 12935 5405 13007 5461
rect 13825 5476 13897 5499
rect 13825 5442 13844 5476
rect 13878 5442 13897 5476
rect 12935 5371 12954 5405
rect 12988 5371 13007 5405
rect 12935 5315 13007 5371
rect 12935 5281 12954 5315
rect 12988 5281 13007 5315
rect 12935 5225 13007 5281
rect 12935 5191 12954 5225
rect 12988 5191 13007 5225
rect 12935 5135 13007 5191
rect 12935 5101 12954 5135
rect 12988 5101 13007 5135
rect 12935 5045 13007 5101
rect 12935 5011 12954 5045
rect 12988 5011 13007 5045
rect 12935 4955 13007 5011
rect 12935 4921 12954 4955
rect 12988 4921 13007 4955
rect 12935 4865 13007 4921
rect 12935 4831 12954 4865
rect 12988 4831 13007 4865
rect 12935 4775 13007 4831
rect 12935 4741 12954 4775
rect 12988 4741 13007 4775
rect 13825 5386 13897 5442
rect 13825 5352 13844 5386
rect 13878 5352 13897 5386
rect 13825 5296 13897 5352
rect 13825 5262 13844 5296
rect 13878 5262 13897 5296
rect 13825 5206 13897 5262
rect 13825 5172 13844 5206
rect 13878 5172 13897 5206
rect 13825 5116 13897 5172
rect 13825 5082 13844 5116
rect 13878 5082 13897 5116
rect 13825 5026 13897 5082
rect 13825 4992 13844 5026
rect 13878 4992 13897 5026
rect 13825 4936 13897 4992
rect 13825 4902 13844 4936
rect 13878 4902 13897 4936
rect 13825 4846 13897 4902
rect 13825 4812 13844 4846
rect 13878 4812 13897 4846
rect 13825 4756 13897 4812
rect 12935 4681 13007 4741
rect 13825 4722 13844 4756
rect 13878 4722 13897 4756
rect 13825 4681 13897 4722
rect 12935 4662 13897 4681
rect 12935 4628 13032 4662
rect 13066 4628 13122 4662
rect 13156 4628 13212 4662
rect 13246 4628 13302 4662
rect 13336 4628 13392 4662
rect 13426 4628 13482 4662
rect 13516 4628 13572 4662
rect 13606 4628 13662 4662
rect 13696 4628 13752 4662
rect 13786 4628 13897 4662
rect 12935 4609 13897 4628
rect 14585 5572 15547 5591
rect 14585 5538 14716 5572
rect 14750 5538 14806 5572
rect 14840 5538 14896 5572
rect 14930 5538 14986 5572
rect 15020 5538 15076 5572
rect 15110 5538 15166 5572
rect 15200 5538 15256 5572
rect 15290 5538 15346 5572
rect 15380 5538 15436 5572
rect 15470 5538 15547 5572
rect 14585 5519 15547 5538
rect 14585 5515 14657 5519
rect 14585 5481 14604 5515
rect 14638 5481 14657 5515
rect 14585 5425 14657 5481
rect 15475 5496 15547 5519
rect 15475 5462 15494 5496
rect 15528 5462 15547 5496
rect 14585 5391 14604 5425
rect 14638 5391 14657 5425
rect 14585 5335 14657 5391
rect 14585 5301 14604 5335
rect 14638 5301 14657 5335
rect 14585 5245 14657 5301
rect 14585 5211 14604 5245
rect 14638 5211 14657 5245
rect 14585 5155 14657 5211
rect 14585 5121 14604 5155
rect 14638 5121 14657 5155
rect 14585 5065 14657 5121
rect 14585 5031 14604 5065
rect 14638 5031 14657 5065
rect 14585 4975 14657 5031
rect 14585 4941 14604 4975
rect 14638 4941 14657 4975
rect 14585 4885 14657 4941
rect 14585 4851 14604 4885
rect 14638 4851 14657 4885
rect 14585 4795 14657 4851
rect 14585 4761 14604 4795
rect 14638 4761 14657 4795
rect 15475 5406 15547 5462
rect 15475 5372 15494 5406
rect 15528 5372 15547 5406
rect 15475 5316 15547 5372
rect 15475 5282 15494 5316
rect 15528 5282 15547 5316
rect 15475 5226 15547 5282
rect 15475 5192 15494 5226
rect 15528 5192 15547 5226
rect 15475 5136 15547 5192
rect 15475 5102 15494 5136
rect 15528 5102 15547 5136
rect 15475 5046 15547 5102
rect 15475 5012 15494 5046
rect 15528 5012 15547 5046
rect 15475 4956 15547 5012
rect 15475 4922 15494 4956
rect 15528 4922 15547 4956
rect 15475 4866 15547 4922
rect 15475 4832 15494 4866
rect 15528 4832 15547 4866
rect 15475 4776 15547 4832
rect 14585 4701 14657 4761
rect 15475 4742 15494 4776
rect 15528 4742 15547 4776
rect 15475 4701 15547 4742
rect 14585 4682 15547 4701
rect 14585 4648 14682 4682
rect 14716 4648 14772 4682
rect 14806 4648 14862 4682
rect 14896 4648 14952 4682
rect 14986 4648 15042 4682
rect 15076 4648 15132 4682
rect 15166 4648 15222 4682
rect 15256 4648 15312 4682
rect 15346 4648 15402 4682
rect 15436 4648 15547 4682
rect 14585 4629 15547 4648
<< mvpsubdiff >>
rect 23004 17346 24388 17358
rect 23004 17312 23135 17346
rect 23169 17312 23203 17346
rect 23237 17312 23271 17346
rect 23305 17312 23339 17346
rect 23373 17312 23407 17346
rect 23441 17312 23475 17346
rect 23509 17312 23543 17346
rect 23577 17312 23611 17346
rect 23645 17312 23679 17346
rect 23713 17312 23747 17346
rect 23781 17312 23815 17346
rect 23849 17312 23883 17346
rect 23917 17312 23951 17346
rect 23985 17312 24019 17346
rect 24053 17312 24087 17346
rect 24121 17312 24155 17346
rect 24189 17312 24223 17346
rect 24257 17312 24388 17346
rect 23004 17300 24388 17312
rect 23004 17231 23062 17300
rect 23004 17197 23016 17231
rect 23050 17197 23062 17231
rect 24330 17231 24388 17300
rect 23004 17163 23062 17197
rect 23004 17129 23016 17163
rect 23050 17129 23062 17163
rect 24330 17197 24342 17231
rect 24376 17197 24388 17231
rect 24330 17163 24388 17197
rect 23004 17095 23062 17129
rect 23004 17061 23016 17095
rect 23050 17061 23062 17095
rect 23004 17027 23062 17061
rect 23004 16993 23016 17027
rect 23050 16993 23062 17027
rect 23004 16959 23062 16993
rect 23004 16925 23016 16959
rect 23050 16925 23062 16959
rect 23004 16891 23062 16925
rect 23004 16857 23016 16891
rect 23050 16857 23062 16891
rect 23004 16823 23062 16857
rect 23004 16789 23016 16823
rect 23050 16789 23062 16823
rect 23004 16755 23062 16789
rect 23004 16721 23016 16755
rect 23050 16721 23062 16755
rect 23004 16687 23062 16721
rect 23004 16653 23016 16687
rect 23050 16653 23062 16687
rect 23004 16619 23062 16653
rect 23004 16585 23016 16619
rect 23050 16585 23062 16619
rect 23004 16551 23062 16585
rect 23004 16517 23016 16551
rect 23050 16517 23062 16551
rect 23004 16483 23062 16517
rect 23004 16449 23016 16483
rect 23050 16449 23062 16483
rect 23004 16415 23062 16449
rect 23004 16381 23016 16415
rect 23050 16381 23062 16415
rect 23004 16347 23062 16381
rect 23004 16313 23016 16347
rect 23050 16313 23062 16347
rect 23004 16279 23062 16313
rect 23004 16245 23016 16279
rect 23050 16245 23062 16279
rect 23004 16211 23062 16245
rect 23004 16177 23016 16211
rect 23050 16177 23062 16211
rect 23004 16143 23062 16177
rect 23004 16109 23016 16143
rect 23050 16109 23062 16143
rect 24330 17129 24342 17163
rect 24376 17129 24388 17163
rect 24330 17095 24388 17129
rect 24330 17061 24342 17095
rect 24376 17061 24388 17095
rect 24330 17027 24388 17061
rect 24330 16993 24342 17027
rect 24376 16993 24388 17027
rect 24330 16959 24388 16993
rect 24330 16925 24342 16959
rect 24376 16925 24388 16959
rect 24330 16891 24388 16925
rect 24330 16857 24342 16891
rect 24376 16857 24388 16891
rect 24330 16823 24388 16857
rect 24330 16789 24342 16823
rect 24376 16789 24388 16823
rect 24330 16755 24388 16789
rect 24330 16721 24342 16755
rect 24376 16721 24388 16755
rect 24330 16687 24388 16721
rect 24330 16653 24342 16687
rect 24376 16653 24388 16687
rect 24330 16619 24388 16653
rect 24330 16585 24342 16619
rect 24376 16585 24388 16619
rect 24330 16551 24388 16585
rect 24330 16517 24342 16551
rect 24376 16517 24388 16551
rect 24330 16483 24388 16517
rect 24330 16449 24342 16483
rect 24376 16449 24388 16483
rect 24330 16415 24388 16449
rect 24330 16381 24342 16415
rect 24376 16381 24388 16415
rect 24330 16347 24388 16381
rect 24330 16313 24342 16347
rect 24376 16313 24388 16347
rect 24330 16279 24388 16313
rect 24330 16245 24342 16279
rect 24376 16245 24388 16279
rect 24330 16211 24388 16245
rect 24330 16177 24342 16211
rect 24376 16177 24388 16211
rect 24330 16143 24388 16177
rect 23004 16075 23062 16109
rect 23004 16041 23016 16075
rect 23050 16041 23062 16075
rect 24330 16109 24342 16143
rect 24376 16109 24388 16143
rect 24330 16075 24388 16109
rect 23004 15972 23062 16041
rect 24330 16041 24342 16075
rect 24376 16041 24388 16075
rect 24330 15972 24388 16041
rect 23004 15960 24388 15972
rect 23004 15926 23135 15960
rect 23169 15926 23203 15960
rect 23237 15926 23271 15960
rect 23305 15926 23339 15960
rect 23373 15926 23407 15960
rect 23441 15926 23475 15960
rect 23509 15926 23543 15960
rect 23577 15926 23611 15960
rect 23645 15926 23679 15960
rect 23713 15926 23747 15960
rect 23781 15926 23815 15960
rect 23849 15926 23883 15960
rect 23917 15926 23951 15960
rect 23985 15926 24019 15960
rect 24053 15926 24087 15960
rect 24121 15926 24155 15960
rect 24189 15926 24223 15960
rect 24257 15926 24388 15960
rect 23004 15914 24388 15926
rect -9119 11565 -3275 11608
rect -9119 11531 -8832 11565
rect -8798 11531 -8764 11565
rect -8730 11531 -8696 11565
rect -8662 11531 -8628 11565
rect -8594 11531 -8560 11565
rect -8526 11531 -8492 11565
rect -8458 11531 -8424 11565
rect -8390 11531 -8356 11565
rect -8322 11531 -8288 11565
rect -8254 11531 -8220 11565
rect -8186 11531 -8152 11565
rect -8118 11531 -8084 11565
rect -8050 11531 -8016 11565
rect -7982 11531 -7948 11565
rect -7914 11531 -7880 11565
rect -7846 11531 -7812 11565
rect -7778 11531 -7744 11565
rect -7710 11531 -7676 11565
rect -7642 11531 -7608 11565
rect -7574 11531 -7540 11565
rect -7506 11531 -7472 11565
rect -7438 11531 -7404 11565
rect -7370 11531 -7336 11565
rect -7302 11531 -7268 11565
rect -7234 11531 -7200 11565
rect -7166 11531 -7132 11565
rect -7098 11531 -7064 11565
rect -7030 11531 -6996 11565
rect -6962 11531 -6928 11565
rect -6894 11531 -6860 11565
rect -6826 11531 -6792 11565
rect -6758 11531 -6724 11565
rect -6690 11531 -6656 11565
rect -6622 11531 -6588 11565
rect -6554 11531 -6520 11565
rect -6486 11531 -6452 11565
rect -6418 11531 -6384 11565
rect -6350 11531 -6316 11565
rect -6282 11531 -6248 11565
rect -6214 11531 -6180 11565
rect -6146 11531 -6112 11565
rect -6078 11531 -6044 11565
rect -6010 11531 -5976 11565
rect -5942 11531 -5908 11565
rect -5874 11531 -5840 11565
rect -5806 11531 -5772 11565
rect -5738 11531 -5704 11565
rect -5670 11531 -5636 11565
rect -5602 11531 -5568 11565
rect -5534 11531 -5500 11565
rect -5466 11531 -5432 11565
rect -5398 11531 -5364 11565
rect -5330 11531 -5296 11565
rect -5262 11531 -5228 11565
rect -5194 11531 -5160 11565
rect -5126 11531 -5092 11565
rect -5058 11531 -5024 11565
rect -4990 11531 -4956 11565
rect -4922 11531 -4888 11565
rect -4854 11531 -4820 11565
rect -4786 11531 -4752 11565
rect -4718 11531 -4684 11565
rect -4650 11531 -4616 11565
rect -4582 11531 -4548 11565
rect -4514 11531 -4480 11565
rect -4446 11531 -4412 11565
rect -4378 11531 -4344 11565
rect -4310 11531 -4276 11565
rect -4242 11531 -4208 11565
rect -4174 11531 -4140 11565
rect -4106 11531 -4072 11565
rect -4038 11531 -4004 11565
rect -3970 11531 -3936 11565
rect -3902 11531 -3868 11565
rect -3834 11531 -3800 11565
rect -3766 11531 -3732 11565
rect -3698 11531 -3664 11565
rect -3630 11531 -3596 11565
rect -3562 11531 -3275 11565
rect -9119 11490 -3275 11531
rect -9119 11375 -9005 11490
rect -9119 11341 -9081 11375
rect -9047 11341 -9005 11375
rect -9119 11307 -9005 11341
rect -9119 11273 -9081 11307
rect -9047 11273 -9005 11307
rect -9119 11239 -9005 11273
rect -3402 11335 -3275 11490
rect -3402 11301 -3355 11335
rect -3321 11301 -3275 11335
rect -3402 11267 -3275 11301
rect -9119 11205 -9081 11239
rect -9047 11205 -9005 11239
rect -9119 11171 -9005 11205
rect -9119 11137 -9081 11171
rect -9047 11137 -9005 11171
rect -3402 11233 -3355 11267
rect -3321 11233 -3275 11267
rect -3402 11199 -3275 11233
rect -3402 11165 -3355 11199
rect -3321 11165 -3275 11199
rect -9119 11103 -9005 11137
rect -9119 11069 -9081 11103
rect -9047 11069 -9005 11103
rect -9119 11035 -9005 11069
rect -9119 11001 -9081 11035
rect -9047 11001 -9005 11035
rect -9119 10967 -9005 11001
rect -9119 10933 -9081 10967
rect -9047 10933 -9005 10967
rect -9119 10899 -9005 10933
rect -9119 10865 -9081 10899
rect -9047 10865 -9005 10899
rect -9119 10831 -9005 10865
rect -9119 10797 -9081 10831
rect -9047 10797 -9005 10831
rect -9119 10763 -9005 10797
rect -9119 10729 -9081 10763
rect -9047 10729 -9005 10763
rect -9119 10695 -9005 10729
rect -9119 10661 -9081 10695
rect -9047 10661 -9005 10695
rect -9119 10627 -9005 10661
rect -9119 10593 -9081 10627
rect -9047 10593 -9005 10627
rect -9119 10559 -9005 10593
rect -9119 10525 -9081 10559
rect -9047 10525 -9005 10559
rect -9119 10491 -9005 10525
rect -9119 10457 -9081 10491
rect -9047 10457 -9005 10491
rect -9119 10423 -9005 10457
rect -9119 10389 -9081 10423
rect -9047 10389 -9005 10423
rect -9119 10355 -9005 10389
rect -9119 10321 -9081 10355
rect -9047 10321 -9005 10355
rect -9119 10287 -9005 10321
rect -9119 10253 -9081 10287
rect -9047 10253 -9005 10287
rect -9119 10219 -9005 10253
rect -9119 10185 -9081 10219
rect -9047 10185 -9005 10219
rect -9119 10151 -9005 10185
rect -3402 11131 -3275 11165
rect -3402 11097 -3355 11131
rect -3321 11097 -3275 11131
rect -3402 11063 -3275 11097
rect -3402 11029 -3355 11063
rect -3321 11029 -3275 11063
rect -3402 10995 -3275 11029
rect -3402 10961 -3355 10995
rect -3321 10961 -3275 10995
rect -3402 10927 -3275 10961
rect -3402 10893 -3355 10927
rect -3321 10893 -3275 10927
rect -3402 10859 -3275 10893
rect -3402 10825 -3355 10859
rect -3321 10825 -3275 10859
rect -3402 10791 -3275 10825
rect -3402 10757 -3355 10791
rect -3321 10757 -3275 10791
rect -3402 10723 -3275 10757
rect -3402 10689 -3355 10723
rect -3321 10689 -3275 10723
rect -3402 10655 -3275 10689
rect -3402 10621 -3355 10655
rect -3321 10621 -3275 10655
rect -3402 10587 -3275 10621
rect -3402 10553 -3355 10587
rect -3321 10553 -3275 10587
rect -3402 10519 -3275 10553
rect -3402 10485 -3355 10519
rect -3321 10485 -3275 10519
rect -3402 10451 -3275 10485
rect -3402 10417 -3355 10451
rect -3321 10417 -3275 10451
rect -3402 10383 -3275 10417
rect -3402 10349 -3355 10383
rect -3321 10349 -3275 10383
rect -3402 10315 -3275 10349
rect -3402 10281 -3355 10315
rect -3321 10281 -3275 10315
rect -3402 10247 -3275 10281
rect -3402 10213 -3355 10247
rect -3321 10213 -3275 10247
rect -3402 10179 -3275 10213
rect -9119 10117 -9081 10151
rect -9047 10117 -9005 10151
rect -9119 10083 -9005 10117
rect -9119 10049 -9081 10083
rect -9047 10049 -9005 10083
rect -3402 10145 -3355 10179
rect -3321 10145 -3275 10179
rect -3402 10111 -3275 10145
rect -3402 10077 -3355 10111
rect -3321 10077 -3275 10111
rect -9119 10015 -9005 10049
rect -9119 9981 -9081 10015
rect -9047 9981 -9005 10015
rect -9119 9947 -9005 9981
rect -9119 9913 -9081 9947
rect -9047 9913 -9005 9947
rect -9119 9879 -9005 9913
rect -3402 10043 -3275 10077
rect -3402 10009 -3355 10043
rect -3321 10009 -3275 10043
rect -3402 9975 -3275 10009
rect -3402 9941 -3355 9975
rect -3321 9941 -3275 9975
rect -3402 9907 -3275 9941
rect -9119 9845 -9081 9879
rect -9047 9845 -9005 9879
rect -9119 9811 -9005 9845
rect -9119 9777 -9081 9811
rect -9047 9777 -9005 9811
rect -3402 9873 -3355 9907
rect -3321 9873 -3275 9907
rect -3402 9839 -3275 9873
rect -3402 9805 -3355 9839
rect -3321 9805 -3275 9839
rect -9119 9743 -9005 9777
rect -9119 9709 -9081 9743
rect -9047 9709 -9005 9743
rect -9119 9675 -9005 9709
rect -9119 9641 -9081 9675
rect -9047 9641 -9005 9675
rect -9119 9607 -9005 9641
rect -9119 9573 -9081 9607
rect -9047 9573 -9005 9607
rect -9119 9539 -9005 9573
rect -9119 9505 -9081 9539
rect -9047 9505 -9005 9539
rect -9119 9471 -9005 9505
rect -9119 9437 -9081 9471
rect -9047 9437 -9005 9471
rect -9119 9403 -9005 9437
rect -9119 9369 -9081 9403
rect -9047 9369 -9005 9403
rect -9119 9335 -9005 9369
rect -9119 9301 -9081 9335
rect -9047 9301 -9005 9335
rect -9119 9267 -9005 9301
rect -9119 9233 -9081 9267
rect -9047 9233 -9005 9267
rect -9119 9199 -9005 9233
rect -9119 9165 -9081 9199
rect -9047 9165 -9005 9199
rect -9119 9131 -9005 9165
rect -9119 9097 -9081 9131
rect -9047 9097 -9005 9131
rect -9119 9063 -9005 9097
rect -9119 9029 -9081 9063
rect -9047 9029 -9005 9063
rect -9119 8995 -9005 9029
rect -9119 8961 -9081 8995
rect -9047 8961 -9005 8995
rect -9119 8927 -9005 8961
rect -9119 8893 -9081 8927
rect -9047 8893 -9005 8927
rect -9119 8859 -9005 8893
rect -9119 8825 -9081 8859
rect -9047 8825 -9005 8859
rect -9119 8791 -9005 8825
rect -3402 9771 -3275 9805
rect -3402 9737 -3355 9771
rect -3321 9737 -3275 9771
rect -3402 9703 -3275 9737
rect -3402 9669 -3355 9703
rect -3321 9669 -3275 9703
rect -3402 9635 -3275 9669
rect -3402 9601 -3355 9635
rect -3321 9601 -3275 9635
rect -3402 9567 -3275 9601
rect -3402 9533 -3355 9567
rect -3321 9533 -3275 9567
rect -3402 9499 -3275 9533
rect -3402 9465 -3355 9499
rect -3321 9465 -3275 9499
rect -3402 9431 -3275 9465
rect -3402 9397 -3355 9431
rect -3321 9397 -3275 9431
rect -3402 9363 -3275 9397
rect -3402 9329 -3355 9363
rect -3321 9329 -3275 9363
rect -3402 9295 -3275 9329
rect -3402 9261 -3355 9295
rect -3321 9261 -3275 9295
rect -3402 9227 -3275 9261
rect -3402 9193 -3355 9227
rect -3321 9193 -3275 9227
rect -3402 9159 -3275 9193
rect -3402 9125 -3355 9159
rect -3321 9125 -3275 9159
rect -3402 9091 -3275 9125
rect -3402 9057 -3355 9091
rect -3321 9057 -3275 9091
rect -3402 9023 -3275 9057
rect -3402 8989 -3355 9023
rect -3321 8989 -3275 9023
rect -3402 8955 -3275 8989
rect -3402 8921 -3355 8955
rect -3321 8921 -3275 8955
rect -3402 8887 -3275 8921
rect -3402 8853 -3355 8887
rect -3321 8853 -3275 8887
rect -3402 8819 -3275 8853
rect -9119 8757 -9081 8791
rect -9047 8757 -9005 8791
rect -9119 8723 -9005 8757
rect -9119 8689 -9081 8723
rect -9047 8689 -9005 8723
rect -3402 8785 -3355 8819
rect -3321 8785 -3275 8819
rect -3402 8751 -3275 8785
rect -3402 8717 -3355 8751
rect -3321 8717 -3275 8751
rect -9119 8655 -9005 8689
rect -9119 8621 -9081 8655
rect -9047 8621 -9005 8655
rect -9119 8440 -9005 8621
rect -3402 8683 -3275 8717
rect -3402 8649 -3355 8683
rect -3321 8649 -3275 8683
rect -3402 8615 -3275 8649
rect -3402 8581 -3355 8615
rect -3321 8581 -3275 8615
rect -3402 8440 -3275 8581
rect -9119 8399 -3275 8440
rect -9119 8365 -8813 8399
rect -8779 8365 -8745 8399
rect -8711 8365 -8677 8399
rect -8643 8365 -8609 8399
rect -8575 8365 -8541 8399
rect -8507 8365 -8473 8399
rect -8439 8365 -8405 8399
rect -8371 8365 -8337 8399
rect -8303 8365 -8269 8399
rect -8235 8365 -8201 8399
rect -8167 8365 -8133 8399
rect -8099 8365 -8065 8399
rect -8031 8365 -7997 8399
rect -7963 8365 -7929 8399
rect -7895 8365 -7861 8399
rect -7827 8365 -7793 8399
rect -7759 8365 -7725 8399
rect -7691 8365 -7657 8399
rect -7623 8365 -7589 8399
rect -7555 8365 -7521 8399
rect -7487 8365 -7453 8399
rect -7419 8365 -7385 8399
rect -7351 8365 -7317 8399
rect -7283 8365 -7249 8399
rect -7215 8365 -7181 8399
rect -7147 8365 -7113 8399
rect -7079 8365 -7045 8399
rect -7011 8365 -6977 8399
rect -6943 8365 -6909 8399
rect -6875 8365 -6841 8399
rect -6807 8365 -6773 8399
rect -6739 8365 -6705 8399
rect -6671 8365 -6637 8399
rect -6603 8365 -6569 8399
rect -6535 8365 -6501 8399
rect -6467 8365 -6433 8399
rect -6399 8365 -6365 8399
rect -6331 8365 -6297 8399
rect -6263 8365 -6229 8399
rect -6195 8365 -6161 8399
rect -6127 8365 -6093 8399
rect -6059 8365 -6025 8399
rect -5991 8365 -5957 8399
rect -5923 8365 -5889 8399
rect -5855 8365 -5821 8399
rect -5787 8365 -5753 8399
rect -5719 8365 -5685 8399
rect -5651 8365 -5617 8399
rect -5583 8365 -5549 8399
rect -5515 8365 -5481 8399
rect -5447 8365 -5413 8399
rect -5379 8365 -5345 8399
rect -5311 8365 -5277 8399
rect -5243 8365 -5209 8399
rect -5175 8365 -5141 8399
rect -5107 8365 -5073 8399
rect -5039 8365 -5005 8399
rect -4971 8365 -4937 8399
rect -4903 8365 -4869 8399
rect -4835 8365 -4801 8399
rect -4767 8365 -4733 8399
rect -4699 8365 -4665 8399
rect -4631 8365 -4597 8399
rect -4563 8365 -4529 8399
rect -4495 8365 -4461 8399
rect -4427 8365 -4393 8399
rect -4359 8365 -4325 8399
rect -4291 8365 -4257 8399
rect -4223 8365 -4189 8399
rect -4155 8365 -4121 8399
rect -4087 8365 -4053 8399
rect -4019 8365 -3985 8399
rect -3951 8365 -3917 8399
rect -3883 8365 -3849 8399
rect -3815 8365 -3781 8399
rect -3747 8365 -3713 8399
rect -3679 8365 -3645 8399
rect -3611 8365 -3577 8399
rect -3543 8365 -3275 8399
rect -9119 8326 -3275 8365
rect -7992 7859 -3398 7882
rect -7992 7825 -7749 7859
rect -7715 7825 -7681 7859
rect -7647 7825 -7613 7859
rect -7579 7825 -7545 7859
rect -7511 7825 -7477 7859
rect -7443 7825 -7409 7859
rect -7375 7825 -7341 7859
rect -7307 7825 -7273 7859
rect -7239 7825 -7205 7859
rect -7171 7825 -7137 7859
rect -7103 7825 -7069 7859
rect -7035 7825 -7001 7859
rect -6967 7825 -6933 7859
rect -6899 7825 -6865 7859
rect -6831 7825 -6797 7859
rect -6763 7825 -6729 7859
rect -6695 7825 -6661 7859
rect -6627 7825 -6593 7859
rect -6559 7825 -6525 7859
rect -6491 7825 -6457 7859
rect -6423 7825 -6389 7859
rect -6355 7825 -6321 7859
rect -6287 7825 -6253 7859
rect -6219 7825 -6185 7859
rect -6151 7825 -6117 7859
rect -6083 7825 -6049 7859
rect -6015 7825 -5981 7859
rect -5947 7825 -5913 7859
rect -5879 7825 -5845 7859
rect -5811 7825 -5777 7859
rect -5743 7825 -5709 7859
rect -5675 7825 -5641 7859
rect -5607 7825 -5573 7859
rect -5539 7825 -5505 7859
rect -5471 7825 -5437 7859
rect -5403 7825 -5369 7859
rect -5335 7825 -5301 7859
rect -5267 7825 -5233 7859
rect -5199 7825 -5165 7859
rect -5131 7825 -5097 7859
rect -5063 7825 -5029 7859
rect -4995 7825 -4961 7859
rect -4927 7825 -4893 7859
rect -4859 7825 -4825 7859
rect -4791 7825 -4757 7859
rect -4723 7825 -4689 7859
rect -4655 7825 -4621 7859
rect -4587 7825 -4553 7859
rect -4519 7825 -4485 7859
rect -4451 7825 -4417 7859
rect -4383 7825 -4349 7859
rect -4315 7825 -4281 7859
rect -4247 7825 -4213 7859
rect -4179 7825 -4145 7859
rect -4111 7825 -4077 7859
rect -4043 7825 -4009 7859
rect -3975 7825 -3941 7859
rect -3907 7825 -3873 7859
rect -3839 7825 -3805 7859
rect -3771 7825 -3737 7859
rect -3703 7825 -3669 7859
rect -3635 7825 -3601 7859
rect -3567 7825 -3398 7859
rect -7992 7806 -3398 7825
rect -7992 7682 -7910 7806
rect -7992 7648 -7968 7682
rect -7934 7648 -7910 7682
rect -7992 7614 -7910 7648
rect -3480 7694 -3398 7806
rect -3480 7660 -3456 7694
rect -3422 7660 -3398 7694
rect -3480 7626 -3398 7660
rect -7992 7580 -7968 7614
rect -7934 7580 -7910 7614
rect -7992 7546 -7910 7580
rect -7992 7512 -7968 7546
rect -7934 7512 -7910 7546
rect -3480 7592 -3456 7626
rect -3422 7592 -3398 7626
rect -3480 7558 -3398 7592
rect -7992 7478 -7910 7512
rect -7992 7444 -7968 7478
rect -7934 7444 -7910 7478
rect -7992 7410 -7910 7444
rect -7992 7376 -7968 7410
rect -7934 7376 -7910 7410
rect -7992 7342 -7910 7376
rect -7992 7308 -7968 7342
rect -7934 7308 -7910 7342
rect -7992 7274 -7910 7308
rect -7992 7240 -7968 7274
rect -7934 7240 -7910 7274
rect -7992 7206 -7910 7240
rect -7992 7172 -7968 7206
rect -7934 7172 -7910 7206
rect -7992 7138 -7910 7172
rect -7992 7104 -7968 7138
rect -7934 7104 -7910 7138
rect -7992 7070 -7910 7104
rect -7992 7036 -7968 7070
rect -7934 7036 -7910 7070
rect -7992 7002 -7910 7036
rect -7992 6968 -7968 7002
rect -7934 6968 -7910 7002
rect -7992 6934 -7910 6968
rect -7992 6900 -7968 6934
rect -7934 6900 -7910 6934
rect -7992 6866 -7910 6900
rect -7992 6832 -7968 6866
rect -7934 6832 -7910 6866
rect -7992 6798 -7910 6832
rect -7992 6764 -7968 6798
rect -7934 6764 -7910 6798
rect -7992 6730 -7910 6764
rect -7992 6696 -7968 6730
rect -7934 6696 -7910 6730
rect -7992 6662 -7910 6696
rect -7992 6628 -7968 6662
rect -7934 6628 -7910 6662
rect -7992 6594 -7910 6628
rect -7992 6560 -7968 6594
rect -7934 6560 -7910 6594
rect -7992 6526 -7910 6560
rect -7992 6492 -7968 6526
rect -7934 6492 -7910 6526
rect -7992 6458 -7910 6492
rect -7992 6424 -7968 6458
rect -7934 6424 -7910 6458
rect -7992 6390 -7910 6424
rect -7992 6356 -7968 6390
rect -7934 6356 -7910 6390
rect -7992 6322 -7910 6356
rect -7992 6288 -7968 6322
rect -7934 6288 -7910 6322
rect -7992 6254 -7910 6288
rect -7992 6220 -7968 6254
rect -7934 6220 -7910 6254
rect -7992 6186 -7910 6220
rect -7992 6152 -7968 6186
rect -7934 6152 -7910 6186
rect -7992 6118 -7910 6152
rect -7992 6084 -7968 6118
rect -7934 6084 -7910 6118
rect -7992 6050 -7910 6084
rect -7992 6016 -7968 6050
rect -7934 6016 -7910 6050
rect -7992 5982 -7910 6016
rect -7992 5948 -7968 5982
rect -7934 5948 -7910 5982
rect -7992 5914 -7910 5948
rect -7992 5880 -7968 5914
rect -7934 5880 -7910 5914
rect -7992 5846 -7910 5880
rect -7992 5812 -7968 5846
rect -7934 5812 -7910 5846
rect -7992 5778 -7910 5812
rect -7992 5744 -7968 5778
rect -7934 5744 -7910 5778
rect -7992 5710 -7910 5744
rect -7992 5676 -7968 5710
rect -7934 5676 -7910 5710
rect -7992 5642 -7910 5676
rect -7992 5608 -7968 5642
rect -7934 5608 -7910 5642
rect -7992 5574 -7910 5608
rect -7992 5540 -7968 5574
rect -7934 5540 -7910 5574
rect -7992 5506 -7910 5540
rect -3480 7524 -3456 7558
rect -3422 7524 -3398 7558
rect -3480 7490 -3398 7524
rect -3480 7456 -3456 7490
rect -3422 7456 -3398 7490
rect -3480 7422 -3398 7456
rect -3480 7388 -3456 7422
rect -3422 7388 -3398 7422
rect -3480 7354 -3398 7388
rect -3480 7320 -3456 7354
rect -3422 7320 -3398 7354
rect -3480 7286 -3398 7320
rect -3480 7252 -3456 7286
rect -3422 7252 -3398 7286
rect -3480 7218 -3398 7252
rect -3480 7184 -3456 7218
rect -3422 7184 -3398 7218
rect -3480 7150 -3398 7184
rect -3480 7116 -3456 7150
rect -3422 7116 -3398 7150
rect 17288 7758 18672 7770
rect 17288 7724 17419 7758
rect 17453 7724 17487 7758
rect 17521 7724 17555 7758
rect 17589 7724 17623 7758
rect 17657 7724 17691 7758
rect 17725 7724 17759 7758
rect 17793 7724 17827 7758
rect 17861 7724 17895 7758
rect 17929 7724 17963 7758
rect 17997 7724 18031 7758
rect 18065 7724 18099 7758
rect 18133 7724 18167 7758
rect 18201 7724 18235 7758
rect 18269 7724 18303 7758
rect 18337 7724 18371 7758
rect 18405 7724 18439 7758
rect 18473 7724 18507 7758
rect 18541 7724 18672 7758
rect 17288 7712 18672 7724
rect 17288 7629 17346 7712
rect 17288 7595 17300 7629
rect 17334 7595 17346 7629
rect 17288 7561 17346 7595
rect 17288 7527 17300 7561
rect 17334 7527 17346 7561
rect 18614 7629 18672 7712
rect 18614 7595 18626 7629
rect 18660 7595 18672 7629
rect 18614 7561 18672 7595
rect 17288 7493 17346 7527
rect 17288 7459 17300 7493
rect 17334 7459 17346 7493
rect 17288 7425 17346 7459
rect 17288 7391 17300 7425
rect 17334 7391 17346 7425
rect 17288 7357 17346 7391
rect 17288 7323 17300 7357
rect 17334 7323 17346 7357
rect 17288 7289 17346 7323
rect 17288 7255 17300 7289
rect 17334 7255 17346 7289
rect -3480 7082 -3398 7116
rect -3480 7048 -3456 7082
rect -3422 7048 -3398 7082
rect -3480 7014 -3398 7048
rect -3480 6980 -3456 7014
rect -3422 6980 -3398 7014
rect -3480 6946 -3398 6980
rect -3480 6912 -3456 6946
rect -3422 6912 -3398 6946
rect -3480 6878 -3398 6912
rect -3480 6844 -3456 6878
rect -3422 6844 -3398 6878
rect -3480 6810 -3398 6844
rect -3480 6776 -3456 6810
rect -3422 6776 -3398 6810
rect -3480 6742 -3398 6776
rect -3480 6708 -3456 6742
rect -3422 6708 -3398 6742
rect -3480 6674 -3398 6708
rect -3480 6640 -3456 6674
rect -3422 6640 -3398 6674
rect -3480 6606 -3398 6640
rect -3480 6572 -3456 6606
rect -3422 6572 -3398 6606
rect -3480 6538 -3398 6572
rect -3480 6504 -3456 6538
rect -3422 6504 -3398 6538
rect -3480 6470 -3398 6504
rect -3480 6436 -3456 6470
rect -3422 6436 -3398 6470
rect -3480 6402 -3398 6436
rect -3480 6368 -3456 6402
rect -3422 6368 -3398 6402
rect -3480 6334 -3398 6368
rect -3480 6300 -3456 6334
rect -3422 6300 -3398 6334
rect -3480 6266 -3398 6300
rect -3480 6232 -3456 6266
rect -3422 6232 -3398 6266
rect -3480 6198 -3398 6232
rect -3480 6164 -3456 6198
rect -3422 6164 -3398 6198
rect -3480 6130 -3398 6164
rect -3480 6096 -3456 6130
rect -3422 6096 -3398 6130
rect -3480 6062 -3398 6096
rect -3480 6028 -3456 6062
rect -3422 6028 -3398 6062
rect -3480 5994 -3398 6028
rect -3480 5960 -3456 5994
rect -3422 5960 -3398 5994
rect -3480 5926 -3398 5960
rect -3480 5892 -3456 5926
rect -3422 5892 -3398 5926
rect -3480 5858 -3398 5892
rect -3480 5824 -3456 5858
rect -3422 5824 -3398 5858
rect -3480 5790 -3398 5824
rect -3480 5756 -3456 5790
rect -3422 5756 -3398 5790
rect -3480 5722 -3398 5756
rect -3480 5688 -3456 5722
rect -3422 5688 -3398 5722
rect -3480 5654 -3398 5688
rect -3480 5620 -3456 5654
rect -3422 5620 -3398 5654
rect -3480 5586 -3398 5620
rect -3480 5552 -3456 5586
rect -3422 5552 -3398 5586
rect -7992 5472 -7968 5506
rect -7934 5472 -7910 5506
rect -7992 5438 -7910 5472
rect -3480 5518 -3398 5552
rect -3480 5484 -3456 5518
rect -3422 5484 -3398 5518
rect -3480 5450 -3398 5484
rect -7992 5404 -7968 5438
rect -7934 5404 -7910 5438
rect -7992 5300 -7910 5404
rect -3480 5416 -3456 5450
rect -3422 5416 -3398 5450
rect -3480 5300 -3398 5416
rect -7992 5279 -3398 5300
rect -7992 5245 -7773 5279
rect -7739 5245 -7705 5279
rect -7671 5245 -7637 5279
rect -7603 5245 -7569 5279
rect -7535 5245 -7501 5279
rect -7467 5245 -7433 5279
rect -7399 5245 -7365 5279
rect -7331 5245 -7297 5279
rect -7263 5245 -7229 5279
rect -7195 5245 -7161 5279
rect -7127 5245 -7093 5279
rect -7059 5245 -7025 5279
rect -6991 5245 -6957 5279
rect -6923 5245 -6889 5279
rect -6855 5245 -6821 5279
rect -6787 5245 -6753 5279
rect -6719 5245 -6685 5279
rect -6651 5245 -6617 5279
rect -6583 5245 -6549 5279
rect -6515 5245 -6481 5279
rect -6447 5245 -6413 5279
rect -6379 5245 -6345 5279
rect -6311 5245 -6277 5279
rect -6243 5245 -6209 5279
rect -6175 5245 -6141 5279
rect -6107 5245 -6073 5279
rect -6039 5245 -6005 5279
rect -5971 5245 -5937 5279
rect -5903 5245 -5869 5279
rect -5835 5245 -5801 5279
rect -5767 5245 -5733 5279
rect -5699 5245 -5665 5279
rect -5631 5245 -5597 5279
rect -5563 5245 -5529 5279
rect -5495 5245 -5461 5279
rect -5427 5245 -5393 5279
rect -5359 5245 -5325 5279
rect -5291 5245 -5257 5279
rect -5223 5245 -5189 5279
rect -5155 5245 -5121 5279
rect -5087 5245 -5053 5279
rect -5019 5245 -4985 5279
rect -4951 5245 -4917 5279
rect -4883 5245 -4849 5279
rect -4815 5245 -4781 5279
rect -4747 5245 -4713 5279
rect -4679 5245 -4645 5279
rect -4611 5245 -4577 5279
rect -4543 5245 -4509 5279
rect -4475 5245 -4441 5279
rect -4407 5245 -4373 5279
rect -4339 5245 -4305 5279
rect -4271 5245 -4237 5279
rect -4203 5245 -4169 5279
rect -4135 5245 -4101 5279
rect -4067 5245 -4033 5279
rect -3999 5245 -3965 5279
rect -3931 5245 -3897 5279
rect -3863 5245 -3829 5279
rect -3795 5245 -3761 5279
rect -3727 5245 -3693 5279
rect -3659 5245 -3625 5279
rect -3591 5245 -3398 5279
rect -7992 5226 -3398 5245
rect 17288 7221 17346 7255
rect 17288 7187 17300 7221
rect 17334 7187 17346 7221
rect 17288 7153 17346 7187
rect 17288 7119 17300 7153
rect 17334 7119 17346 7153
rect 17288 7085 17346 7119
rect 17288 7051 17300 7085
rect 17334 7051 17346 7085
rect 17288 7017 17346 7051
rect 17288 6983 17300 7017
rect 17334 6983 17346 7017
rect 17288 6949 17346 6983
rect 17288 6915 17300 6949
rect 17334 6915 17346 6949
rect 17288 6881 17346 6915
rect 17288 6847 17300 6881
rect 17334 6847 17346 6881
rect 17288 6813 17346 6847
rect 17288 6779 17300 6813
rect 17334 6779 17346 6813
rect 17288 6745 17346 6779
rect 17288 6711 17300 6745
rect 17334 6711 17346 6745
rect 17288 6677 17346 6711
rect 17288 6643 17300 6677
rect 17334 6643 17346 6677
rect 17288 6609 17346 6643
rect 17288 6575 17300 6609
rect 17334 6575 17346 6609
rect 17288 6541 17346 6575
rect 17288 6507 17300 6541
rect 17334 6507 17346 6541
rect 17288 6473 17346 6507
rect 17288 6439 17300 6473
rect 17334 6439 17346 6473
rect 17288 6405 17346 6439
rect 17288 6371 17300 6405
rect 17334 6371 17346 6405
rect 17288 6337 17346 6371
rect 17288 6303 17300 6337
rect 17334 6303 17346 6337
rect 17288 6269 17346 6303
rect 17288 6235 17300 6269
rect 17334 6235 17346 6269
rect 17288 6201 17346 6235
rect 17288 6167 17300 6201
rect 17334 6167 17346 6201
rect 17288 6133 17346 6167
rect 17288 6099 17300 6133
rect 17334 6099 17346 6133
rect 17288 6065 17346 6099
rect 17288 6031 17300 6065
rect 17334 6031 17346 6065
rect 17288 5997 17346 6031
rect 17288 5963 17300 5997
rect 17334 5963 17346 5997
rect 17288 5929 17346 5963
rect 17288 5895 17300 5929
rect 17334 5895 17346 5929
rect 17288 5861 17346 5895
rect 17288 5827 17300 5861
rect 17334 5827 17346 5861
rect 17288 5793 17346 5827
rect 17288 5759 17300 5793
rect 17334 5759 17346 5793
rect 17288 5725 17346 5759
rect 17288 5691 17300 5725
rect 17334 5691 17346 5725
rect 17288 5657 17346 5691
rect 17288 5623 17300 5657
rect 17334 5623 17346 5657
rect 17288 5589 17346 5623
rect 17288 5555 17300 5589
rect 17334 5555 17346 5589
rect 17288 5521 17346 5555
rect 17288 5487 17300 5521
rect 17334 5487 17346 5521
rect 17288 5453 17346 5487
rect 17288 5419 17300 5453
rect 17334 5419 17346 5453
rect 17288 5385 17346 5419
rect 17288 5351 17300 5385
rect 17334 5351 17346 5385
rect 17288 5317 17346 5351
rect 17288 5283 17300 5317
rect 17334 5283 17346 5317
rect 17288 5249 17346 5283
rect 17288 5215 17300 5249
rect 17334 5215 17346 5249
rect 17288 5181 17346 5215
rect 17288 5147 17300 5181
rect 17334 5147 17346 5181
rect 17288 5113 17346 5147
rect 17288 5079 17300 5113
rect 17334 5079 17346 5113
rect 17288 5045 17346 5079
rect 17288 5011 17300 5045
rect 17334 5011 17346 5045
rect 17288 4977 17346 5011
rect 17288 4943 17300 4977
rect 17334 4943 17346 4977
rect 17288 4909 17346 4943
rect 17288 4875 17300 4909
rect 17334 4875 17346 4909
rect 17288 4841 17346 4875
rect 17288 4807 17300 4841
rect 17334 4807 17346 4841
rect 17288 4773 17346 4807
rect 17288 4739 17300 4773
rect 17334 4739 17346 4773
rect 17288 4705 17346 4739
rect 17288 4671 17300 4705
rect 17334 4671 17346 4705
rect 17288 4637 17346 4671
rect 17288 4603 17300 4637
rect 17334 4603 17346 4637
rect 17288 4569 17346 4603
rect 17288 4535 17300 4569
rect 17334 4535 17346 4569
rect 18614 7527 18626 7561
rect 18660 7527 18672 7561
rect 18614 7493 18672 7527
rect 18614 7459 18626 7493
rect 18660 7459 18672 7493
rect 18614 7425 18672 7459
rect 18614 7391 18626 7425
rect 18660 7391 18672 7425
rect 18614 7357 18672 7391
rect 18614 7323 18626 7357
rect 18660 7323 18672 7357
rect 18614 7289 18672 7323
rect 18614 7255 18626 7289
rect 18660 7255 18672 7289
rect 18614 7221 18672 7255
rect 18614 7187 18626 7221
rect 18660 7187 18672 7221
rect 18614 7153 18672 7187
rect 18614 7119 18626 7153
rect 18660 7119 18672 7153
rect 18614 7085 18672 7119
rect 18614 7051 18626 7085
rect 18660 7051 18672 7085
rect 18614 7017 18672 7051
rect 18614 6983 18626 7017
rect 18660 6983 18672 7017
rect 18614 6949 18672 6983
rect 18614 6915 18626 6949
rect 18660 6915 18672 6949
rect 18614 6881 18672 6915
rect 18614 6847 18626 6881
rect 18660 6847 18672 6881
rect 18614 6813 18672 6847
rect 18614 6779 18626 6813
rect 18660 6779 18672 6813
rect 18614 6745 18672 6779
rect 18614 6711 18626 6745
rect 18660 6711 18672 6745
rect 18614 6677 18672 6711
rect 18614 6643 18626 6677
rect 18660 6643 18672 6677
rect 18614 6609 18672 6643
rect 18614 6575 18626 6609
rect 18660 6575 18672 6609
rect 18614 6541 18672 6575
rect 18614 6507 18626 6541
rect 18660 6507 18672 6541
rect 18614 6473 18672 6507
rect 18614 6439 18626 6473
rect 18660 6439 18672 6473
rect 18614 6405 18672 6439
rect 18614 6371 18626 6405
rect 18660 6371 18672 6405
rect 18614 6337 18672 6371
rect 18614 6303 18626 6337
rect 18660 6303 18672 6337
rect 18614 6269 18672 6303
rect 18614 6235 18626 6269
rect 18660 6235 18672 6269
rect 18614 6201 18672 6235
rect 18614 6167 18626 6201
rect 18660 6167 18672 6201
rect 18614 6133 18672 6167
rect 18614 6099 18626 6133
rect 18660 6099 18672 6133
rect 18614 6065 18672 6099
rect 18614 6031 18626 6065
rect 18660 6031 18672 6065
rect 18614 5997 18672 6031
rect 18614 5963 18626 5997
rect 18660 5963 18672 5997
rect 18614 5929 18672 5963
rect 18614 5895 18626 5929
rect 18660 5895 18672 5929
rect 18614 5861 18672 5895
rect 18614 5827 18626 5861
rect 18660 5827 18672 5861
rect 18614 5793 18672 5827
rect 18614 5759 18626 5793
rect 18660 5759 18672 5793
rect 18614 5725 18672 5759
rect 18614 5691 18626 5725
rect 18660 5691 18672 5725
rect 18614 5657 18672 5691
rect 18614 5623 18626 5657
rect 18660 5623 18672 5657
rect 18614 5589 18672 5623
rect 18614 5555 18626 5589
rect 18660 5555 18672 5589
rect 18614 5521 18672 5555
rect 18614 5487 18626 5521
rect 18660 5487 18672 5521
rect 18614 5453 18672 5487
rect 18614 5419 18626 5453
rect 18660 5419 18672 5453
rect 18614 5385 18672 5419
rect 18614 5351 18626 5385
rect 18660 5351 18672 5385
rect 18614 5317 18672 5351
rect 18614 5283 18626 5317
rect 18660 5283 18672 5317
rect 18614 5249 18672 5283
rect 18614 5215 18626 5249
rect 18660 5215 18672 5249
rect 18614 5181 18672 5215
rect 18614 5147 18626 5181
rect 18660 5147 18672 5181
rect 18614 5113 18672 5147
rect 18614 5079 18626 5113
rect 18660 5079 18672 5113
rect 18614 5045 18672 5079
rect 18614 5011 18626 5045
rect 18660 5011 18672 5045
rect 18614 4977 18672 5011
rect 18614 4943 18626 4977
rect 18660 4943 18672 4977
rect 18614 4909 18672 4943
rect 18614 4875 18626 4909
rect 18660 4875 18672 4909
rect 18614 4841 18672 4875
rect 18614 4807 18626 4841
rect 18660 4807 18672 4841
rect 18614 4773 18672 4807
rect 18614 4739 18626 4773
rect 18660 4739 18672 4773
rect 18614 4705 18672 4739
rect 18614 4671 18626 4705
rect 18660 4671 18672 4705
rect 18614 4637 18672 4671
rect 18614 4603 18626 4637
rect 18660 4603 18672 4637
rect 18614 4569 18672 4603
rect 17288 4501 17346 4535
rect 17288 4467 17300 4501
rect 17334 4467 17346 4501
rect 17288 4384 17346 4467
rect 18614 4535 18626 4569
rect 18660 4535 18672 4569
rect 18614 4501 18672 4535
rect 18614 4467 18626 4501
rect 18660 4467 18672 4501
rect 18614 4384 18672 4467
rect 17288 4372 18672 4384
rect 17288 4338 17419 4372
rect 17453 4338 17487 4372
rect 17521 4338 17555 4372
rect 17589 4338 17623 4372
rect 17657 4338 17691 4372
rect 17725 4338 17759 4372
rect 17793 4338 17827 4372
rect 17861 4338 17895 4372
rect 17929 4338 17963 4372
rect 17997 4338 18031 4372
rect 18065 4338 18099 4372
rect 18133 4338 18167 4372
rect 18201 4338 18235 4372
rect 18269 4338 18303 4372
rect 18337 4338 18371 4372
rect 18405 4338 18439 4372
rect 18473 4338 18507 4372
rect 18541 4338 18672 4372
rect 17288 4326 18672 4338
rect 18738 7758 20122 7770
rect 18738 7724 18869 7758
rect 18903 7724 18937 7758
rect 18971 7724 19005 7758
rect 19039 7724 19073 7758
rect 19107 7724 19141 7758
rect 19175 7724 19209 7758
rect 19243 7724 19277 7758
rect 19311 7724 19345 7758
rect 19379 7724 19413 7758
rect 19447 7724 19481 7758
rect 19515 7724 19549 7758
rect 19583 7724 19617 7758
rect 19651 7724 19685 7758
rect 19719 7724 19753 7758
rect 19787 7724 19821 7758
rect 19855 7724 19889 7758
rect 19923 7724 19957 7758
rect 19991 7724 20122 7758
rect 18738 7712 20122 7724
rect 18738 7629 18796 7712
rect 18738 7595 18750 7629
rect 18784 7595 18796 7629
rect 18738 7561 18796 7595
rect 18738 7527 18750 7561
rect 18784 7527 18796 7561
rect 20064 7629 20122 7712
rect 20064 7595 20076 7629
rect 20110 7595 20122 7629
rect 20064 7561 20122 7595
rect 18738 7493 18796 7527
rect 18738 7459 18750 7493
rect 18784 7459 18796 7493
rect 18738 7425 18796 7459
rect 18738 7391 18750 7425
rect 18784 7391 18796 7425
rect 18738 7357 18796 7391
rect 18738 7323 18750 7357
rect 18784 7323 18796 7357
rect 18738 7289 18796 7323
rect 18738 7255 18750 7289
rect 18784 7255 18796 7289
rect 18738 7221 18796 7255
rect 18738 7187 18750 7221
rect 18784 7187 18796 7221
rect 18738 7153 18796 7187
rect 18738 7119 18750 7153
rect 18784 7119 18796 7153
rect 18738 7085 18796 7119
rect 18738 7051 18750 7085
rect 18784 7051 18796 7085
rect 18738 7017 18796 7051
rect 18738 6983 18750 7017
rect 18784 6983 18796 7017
rect 18738 6949 18796 6983
rect 18738 6915 18750 6949
rect 18784 6915 18796 6949
rect 18738 6881 18796 6915
rect 18738 6847 18750 6881
rect 18784 6847 18796 6881
rect 18738 6813 18796 6847
rect 18738 6779 18750 6813
rect 18784 6779 18796 6813
rect 18738 6745 18796 6779
rect 18738 6711 18750 6745
rect 18784 6711 18796 6745
rect 18738 6677 18796 6711
rect 18738 6643 18750 6677
rect 18784 6643 18796 6677
rect 18738 6609 18796 6643
rect 18738 6575 18750 6609
rect 18784 6575 18796 6609
rect 18738 6541 18796 6575
rect 18738 6507 18750 6541
rect 18784 6507 18796 6541
rect 18738 6473 18796 6507
rect 18738 6439 18750 6473
rect 18784 6439 18796 6473
rect 18738 6405 18796 6439
rect 18738 6371 18750 6405
rect 18784 6371 18796 6405
rect 18738 6337 18796 6371
rect 18738 6303 18750 6337
rect 18784 6303 18796 6337
rect 18738 6269 18796 6303
rect 18738 6235 18750 6269
rect 18784 6235 18796 6269
rect 18738 6201 18796 6235
rect 18738 6167 18750 6201
rect 18784 6167 18796 6201
rect 18738 6133 18796 6167
rect 18738 6099 18750 6133
rect 18784 6099 18796 6133
rect 18738 6065 18796 6099
rect 18738 6031 18750 6065
rect 18784 6031 18796 6065
rect 18738 5997 18796 6031
rect 18738 5963 18750 5997
rect 18784 5963 18796 5997
rect 18738 5929 18796 5963
rect 18738 5895 18750 5929
rect 18784 5895 18796 5929
rect 18738 5861 18796 5895
rect 18738 5827 18750 5861
rect 18784 5827 18796 5861
rect 18738 5793 18796 5827
rect 18738 5759 18750 5793
rect 18784 5759 18796 5793
rect 18738 5725 18796 5759
rect 18738 5691 18750 5725
rect 18784 5691 18796 5725
rect 18738 5657 18796 5691
rect 18738 5623 18750 5657
rect 18784 5623 18796 5657
rect 18738 5589 18796 5623
rect 18738 5555 18750 5589
rect 18784 5555 18796 5589
rect 18738 5521 18796 5555
rect 18738 5487 18750 5521
rect 18784 5487 18796 5521
rect 18738 5453 18796 5487
rect 18738 5419 18750 5453
rect 18784 5419 18796 5453
rect 18738 5385 18796 5419
rect 18738 5351 18750 5385
rect 18784 5351 18796 5385
rect 18738 5317 18796 5351
rect 18738 5283 18750 5317
rect 18784 5283 18796 5317
rect 18738 5249 18796 5283
rect 18738 5215 18750 5249
rect 18784 5215 18796 5249
rect 18738 5181 18796 5215
rect 18738 5147 18750 5181
rect 18784 5147 18796 5181
rect 18738 5113 18796 5147
rect 18738 5079 18750 5113
rect 18784 5079 18796 5113
rect 18738 5045 18796 5079
rect 18738 5011 18750 5045
rect 18784 5011 18796 5045
rect 18738 4977 18796 5011
rect 18738 4943 18750 4977
rect 18784 4943 18796 4977
rect 18738 4909 18796 4943
rect 18738 4875 18750 4909
rect 18784 4875 18796 4909
rect 18738 4841 18796 4875
rect 18738 4807 18750 4841
rect 18784 4807 18796 4841
rect 18738 4773 18796 4807
rect 18738 4739 18750 4773
rect 18784 4739 18796 4773
rect 18738 4705 18796 4739
rect 18738 4671 18750 4705
rect 18784 4671 18796 4705
rect 18738 4637 18796 4671
rect 18738 4603 18750 4637
rect 18784 4603 18796 4637
rect 18738 4569 18796 4603
rect 18738 4535 18750 4569
rect 18784 4535 18796 4569
rect 20064 7527 20076 7561
rect 20110 7527 20122 7561
rect 20064 7493 20122 7527
rect 20064 7459 20076 7493
rect 20110 7459 20122 7493
rect 20064 7425 20122 7459
rect 20064 7391 20076 7425
rect 20110 7391 20122 7425
rect 20064 7357 20122 7391
rect 20064 7323 20076 7357
rect 20110 7323 20122 7357
rect 20064 7289 20122 7323
rect 20064 7255 20076 7289
rect 20110 7255 20122 7289
rect 20064 7221 20122 7255
rect 20064 7187 20076 7221
rect 20110 7187 20122 7221
rect 20064 7153 20122 7187
rect 20064 7119 20076 7153
rect 20110 7119 20122 7153
rect 20064 7085 20122 7119
rect 20064 7051 20076 7085
rect 20110 7051 20122 7085
rect 20064 7017 20122 7051
rect 20064 6983 20076 7017
rect 20110 6983 20122 7017
rect 20064 6949 20122 6983
rect 20064 6915 20076 6949
rect 20110 6915 20122 6949
rect 20064 6881 20122 6915
rect 20064 6847 20076 6881
rect 20110 6847 20122 6881
rect 20064 6813 20122 6847
rect 20064 6779 20076 6813
rect 20110 6779 20122 6813
rect 20064 6745 20122 6779
rect 20064 6711 20076 6745
rect 20110 6711 20122 6745
rect 20064 6677 20122 6711
rect 20064 6643 20076 6677
rect 20110 6643 20122 6677
rect 20064 6609 20122 6643
rect 20064 6575 20076 6609
rect 20110 6575 20122 6609
rect 20064 6541 20122 6575
rect 20064 6507 20076 6541
rect 20110 6507 20122 6541
rect 20064 6473 20122 6507
rect 20064 6439 20076 6473
rect 20110 6439 20122 6473
rect 20064 6405 20122 6439
rect 20064 6371 20076 6405
rect 20110 6371 20122 6405
rect 20064 6337 20122 6371
rect 20064 6303 20076 6337
rect 20110 6303 20122 6337
rect 20064 6269 20122 6303
rect 20064 6235 20076 6269
rect 20110 6235 20122 6269
rect 20064 6201 20122 6235
rect 20064 6167 20076 6201
rect 20110 6167 20122 6201
rect 20064 6133 20122 6167
rect 20064 6099 20076 6133
rect 20110 6099 20122 6133
rect 20064 6065 20122 6099
rect 20064 6031 20076 6065
rect 20110 6031 20122 6065
rect 20064 5997 20122 6031
rect 20064 5963 20076 5997
rect 20110 5963 20122 5997
rect 20064 5929 20122 5963
rect 20064 5895 20076 5929
rect 20110 5895 20122 5929
rect 20064 5861 20122 5895
rect 20064 5827 20076 5861
rect 20110 5827 20122 5861
rect 20064 5793 20122 5827
rect 20064 5759 20076 5793
rect 20110 5759 20122 5793
rect 20064 5725 20122 5759
rect 20064 5691 20076 5725
rect 20110 5691 20122 5725
rect 20064 5657 20122 5691
rect 20064 5623 20076 5657
rect 20110 5623 20122 5657
rect 20064 5589 20122 5623
rect 20064 5555 20076 5589
rect 20110 5555 20122 5589
rect 20064 5521 20122 5555
rect 20064 5487 20076 5521
rect 20110 5487 20122 5521
rect 20064 5453 20122 5487
rect 20064 5419 20076 5453
rect 20110 5419 20122 5453
rect 20064 5385 20122 5419
rect 20064 5351 20076 5385
rect 20110 5351 20122 5385
rect 20064 5317 20122 5351
rect 20064 5283 20076 5317
rect 20110 5283 20122 5317
rect 20064 5249 20122 5283
rect 20064 5215 20076 5249
rect 20110 5215 20122 5249
rect 20064 5181 20122 5215
rect 20064 5147 20076 5181
rect 20110 5147 20122 5181
rect 20064 5113 20122 5147
rect 20064 5079 20076 5113
rect 20110 5079 20122 5113
rect 20064 5045 20122 5079
rect 20064 5011 20076 5045
rect 20110 5011 20122 5045
rect 20064 4977 20122 5011
rect 20064 4943 20076 4977
rect 20110 4943 20122 4977
rect 20064 4909 20122 4943
rect 20064 4875 20076 4909
rect 20110 4875 20122 4909
rect 20064 4841 20122 4875
rect 20064 4807 20076 4841
rect 20110 4807 20122 4841
rect 20064 4773 20122 4807
rect 20064 4739 20076 4773
rect 20110 4739 20122 4773
rect 20064 4705 20122 4739
rect 20064 4671 20076 4705
rect 20110 4671 20122 4705
rect 20064 4637 20122 4671
rect 20064 4603 20076 4637
rect 20110 4603 20122 4637
rect 20064 4569 20122 4603
rect 22908 11950 24352 11962
rect 22908 11916 23035 11950
rect 23069 11916 23103 11950
rect 23137 11916 23171 11950
rect 23205 11916 23239 11950
rect 23273 11916 23307 11950
rect 23341 11916 23375 11950
rect 23409 11916 23443 11950
rect 23477 11916 23511 11950
rect 23545 11916 23579 11950
rect 23613 11916 23647 11950
rect 23681 11916 23715 11950
rect 23749 11916 23783 11950
rect 23817 11916 23851 11950
rect 23885 11916 23919 11950
rect 23953 11916 23987 11950
rect 24021 11916 24055 11950
rect 24089 11916 24123 11950
rect 24157 11916 24191 11950
rect 24225 11916 24352 11950
rect 22908 11904 24352 11916
rect 22908 11831 22966 11904
rect 22908 11797 22920 11831
rect 22954 11797 22966 11831
rect 24294 11831 24352 11904
rect 22908 11763 22966 11797
rect 24294 11797 24306 11831
rect 24340 11797 24352 11831
rect 22908 11729 22920 11763
rect 22954 11729 22966 11763
rect 22908 11695 22966 11729
rect 22908 11661 22920 11695
rect 22954 11661 22966 11695
rect 22908 11627 22966 11661
rect 22908 11593 22920 11627
rect 22954 11593 22966 11627
rect 22908 11559 22966 11593
rect 22908 11525 22920 11559
rect 22954 11525 22966 11559
rect 22908 11491 22966 11525
rect 22908 11457 22920 11491
rect 22954 11457 22966 11491
rect 22908 11423 22966 11457
rect 22908 11389 22920 11423
rect 22954 11389 22966 11423
rect 22908 11355 22966 11389
rect 22908 11321 22920 11355
rect 22954 11321 22966 11355
rect 22908 11287 22966 11321
rect 22908 11253 22920 11287
rect 22954 11253 22966 11287
rect 22908 11219 22966 11253
rect 22908 11185 22920 11219
rect 22954 11185 22966 11219
rect 22908 11151 22966 11185
rect 22908 11117 22920 11151
rect 22954 11117 22966 11151
rect 22908 11083 22966 11117
rect 22908 11049 22920 11083
rect 22954 11049 22966 11083
rect 22908 11015 22966 11049
rect 22908 10981 22920 11015
rect 22954 10981 22966 11015
rect 22908 10947 22966 10981
rect 22908 10913 22920 10947
rect 22954 10913 22966 10947
rect 22908 10879 22966 10913
rect 22908 10845 22920 10879
rect 22954 10845 22966 10879
rect 22908 10811 22966 10845
rect 22908 10777 22920 10811
rect 22954 10777 22966 10811
rect 22908 10743 22966 10777
rect 24294 11763 24352 11797
rect 24294 11729 24306 11763
rect 24340 11729 24352 11763
rect 24294 11695 24352 11729
rect 24294 11661 24306 11695
rect 24340 11661 24352 11695
rect 24294 11627 24352 11661
rect 24294 11593 24306 11627
rect 24340 11593 24352 11627
rect 24294 11559 24352 11593
rect 24294 11525 24306 11559
rect 24340 11525 24352 11559
rect 24294 11491 24352 11525
rect 24294 11457 24306 11491
rect 24340 11457 24352 11491
rect 24294 11423 24352 11457
rect 24294 11389 24306 11423
rect 24340 11389 24352 11423
rect 24294 11355 24352 11389
rect 24294 11321 24306 11355
rect 24340 11321 24352 11355
rect 24294 11287 24352 11321
rect 24294 11253 24306 11287
rect 24340 11253 24352 11287
rect 24294 11219 24352 11253
rect 24294 11185 24306 11219
rect 24340 11185 24352 11219
rect 24294 11151 24352 11185
rect 24294 11117 24306 11151
rect 24340 11117 24352 11151
rect 24294 11083 24352 11117
rect 24294 11049 24306 11083
rect 24340 11049 24352 11083
rect 24294 11015 24352 11049
rect 24294 10981 24306 11015
rect 24340 10981 24352 11015
rect 24294 10947 24352 10981
rect 24294 10913 24306 10947
rect 24340 10913 24352 10947
rect 24294 10879 24352 10913
rect 24294 10845 24306 10879
rect 24340 10845 24352 10879
rect 24294 10811 24352 10845
rect 24294 10777 24306 10811
rect 24340 10777 24352 10811
rect 22908 10709 22920 10743
rect 22954 10709 22966 10743
rect 24294 10743 24352 10777
rect 22908 10636 22966 10709
rect 24294 10709 24306 10743
rect 24340 10709 24352 10743
rect 24294 10636 24352 10709
rect 22908 10624 24352 10636
rect 22908 10590 23035 10624
rect 23069 10590 23103 10624
rect 23137 10590 23171 10624
rect 23205 10590 23239 10624
rect 23273 10590 23307 10624
rect 23341 10590 23375 10624
rect 23409 10590 23443 10624
rect 23477 10590 23511 10624
rect 23545 10590 23579 10624
rect 23613 10590 23647 10624
rect 23681 10590 23715 10624
rect 23749 10590 23783 10624
rect 23817 10590 23851 10624
rect 23885 10590 23919 10624
rect 23953 10590 23987 10624
rect 24021 10590 24055 10624
rect 24089 10590 24123 10624
rect 24157 10590 24191 10624
rect 24225 10590 24352 10624
rect 22908 10578 24352 10590
rect 23388 8014 24832 8026
rect 23388 7980 23515 8014
rect 23549 7980 23583 8014
rect 23617 7980 23651 8014
rect 23685 7980 23719 8014
rect 23753 7980 23787 8014
rect 23821 7980 23855 8014
rect 23889 7980 23923 8014
rect 23957 7980 23991 8014
rect 24025 7980 24059 8014
rect 24093 7980 24127 8014
rect 24161 7980 24195 8014
rect 24229 7980 24263 8014
rect 24297 7980 24331 8014
rect 24365 7980 24399 8014
rect 24433 7980 24467 8014
rect 24501 7980 24535 8014
rect 24569 7980 24603 8014
rect 24637 7980 24671 8014
rect 24705 7980 24832 8014
rect 23388 7968 24832 7980
rect 23388 7906 23446 7968
rect 23388 7872 23400 7906
rect 23434 7872 23446 7906
rect 24774 7906 24832 7968
rect 23388 7838 23446 7872
rect 23388 7804 23400 7838
rect 23434 7804 23446 7838
rect 24774 7872 24786 7906
rect 24820 7872 24832 7906
rect 24774 7838 24832 7872
rect 23388 7770 23446 7804
rect 23388 7736 23400 7770
rect 23434 7736 23446 7770
rect 23388 7702 23446 7736
rect 23388 7668 23400 7702
rect 23434 7668 23446 7702
rect 23388 7634 23446 7668
rect 23388 7600 23400 7634
rect 23434 7600 23446 7634
rect 23388 7566 23446 7600
rect 23388 7532 23400 7566
rect 23434 7532 23446 7566
rect 23388 7498 23446 7532
rect 23388 7464 23400 7498
rect 23434 7464 23446 7498
rect 23388 7430 23446 7464
rect 23388 7396 23400 7430
rect 23434 7396 23446 7430
rect 23388 7362 23446 7396
rect 23388 7328 23400 7362
rect 23434 7328 23446 7362
rect 23388 7294 23446 7328
rect 23388 7260 23400 7294
rect 23434 7260 23446 7294
rect 23388 7226 23446 7260
rect 23388 7192 23400 7226
rect 23434 7192 23446 7226
rect 23388 7158 23446 7192
rect 23388 7124 23400 7158
rect 23434 7124 23446 7158
rect 23388 7090 23446 7124
rect 23388 7056 23400 7090
rect 23434 7056 23446 7090
rect 23388 7022 23446 7056
rect 23388 6988 23400 7022
rect 23434 6988 23446 7022
rect 23388 6954 23446 6988
rect 23388 6920 23400 6954
rect 23434 6920 23446 6954
rect 23388 6886 23446 6920
rect 23388 6852 23400 6886
rect 23434 6852 23446 6886
rect 23388 6818 23446 6852
rect 24774 7804 24786 7838
rect 24820 7804 24832 7838
rect 24774 7770 24832 7804
rect 24774 7736 24786 7770
rect 24820 7736 24832 7770
rect 24774 7702 24832 7736
rect 24774 7668 24786 7702
rect 24820 7668 24832 7702
rect 24774 7634 24832 7668
rect 24774 7600 24786 7634
rect 24820 7600 24832 7634
rect 24774 7566 24832 7600
rect 24774 7532 24786 7566
rect 24820 7532 24832 7566
rect 24774 7498 24832 7532
rect 24774 7464 24786 7498
rect 24820 7464 24832 7498
rect 24774 7430 24832 7464
rect 24774 7396 24786 7430
rect 24820 7396 24832 7430
rect 24774 7362 24832 7396
rect 24774 7328 24786 7362
rect 24820 7328 24832 7362
rect 24774 7294 24832 7328
rect 24774 7260 24786 7294
rect 24820 7260 24832 7294
rect 24774 7226 24832 7260
rect 24774 7192 24786 7226
rect 24820 7192 24832 7226
rect 24774 7158 24832 7192
rect 24774 7124 24786 7158
rect 24820 7124 24832 7158
rect 24774 7090 24832 7124
rect 24774 7056 24786 7090
rect 24820 7056 24832 7090
rect 24774 7022 24832 7056
rect 24774 6988 24786 7022
rect 24820 6988 24832 7022
rect 24774 6954 24832 6988
rect 24774 6920 24786 6954
rect 24820 6920 24832 6954
rect 24774 6886 24832 6920
rect 24774 6852 24786 6886
rect 24820 6852 24832 6886
rect 23388 6784 23400 6818
rect 23434 6784 23446 6818
rect 23388 6750 23446 6784
rect 24774 6818 24832 6852
rect 24774 6784 24786 6818
rect 24820 6784 24832 6818
rect 23388 6716 23400 6750
rect 23434 6716 23446 6750
rect 23388 6682 23446 6716
rect 23388 6648 23400 6682
rect 23434 6648 23446 6682
rect 23388 6614 23446 6648
rect 23388 6580 23400 6614
rect 23434 6580 23446 6614
rect 23388 6546 23446 6580
rect 23388 6512 23400 6546
rect 23434 6512 23446 6546
rect 23388 6478 23446 6512
rect 23388 6444 23400 6478
rect 23434 6444 23446 6478
rect 23388 6410 23446 6444
rect 23388 6376 23400 6410
rect 23434 6376 23446 6410
rect 23388 6342 23446 6376
rect 23388 6308 23400 6342
rect 23434 6308 23446 6342
rect 23388 6274 23446 6308
rect 23388 6240 23400 6274
rect 23434 6240 23446 6274
rect 23388 6206 23446 6240
rect 23388 6172 23400 6206
rect 23434 6172 23446 6206
rect 23388 6138 23446 6172
rect 23388 6104 23400 6138
rect 23434 6104 23446 6138
rect 23388 6070 23446 6104
rect 23388 6036 23400 6070
rect 23434 6036 23446 6070
rect 23388 6002 23446 6036
rect 23388 5968 23400 6002
rect 23434 5968 23446 6002
rect 23388 5934 23446 5968
rect 23388 5900 23400 5934
rect 23434 5900 23446 5934
rect 23388 5866 23446 5900
rect 23388 5832 23400 5866
rect 23434 5832 23446 5866
rect 23388 5798 23446 5832
rect 23388 5764 23400 5798
rect 23434 5764 23446 5798
rect 24774 6750 24832 6784
rect 24774 6716 24786 6750
rect 24820 6716 24832 6750
rect 24774 6682 24832 6716
rect 24774 6648 24786 6682
rect 24820 6648 24832 6682
rect 24774 6614 24832 6648
rect 24774 6580 24786 6614
rect 24820 6580 24832 6614
rect 24774 6546 24832 6580
rect 24774 6512 24786 6546
rect 24820 6512 24832 6546
rect 24774 6478 24832 6512
rect 24774 6444 24786 6478
rect 24820 6444 24832 6478
rect 24774 6410 24832 6444
rect 24774 6376 24786 6410
rect 24820 6376 24832 6410
rect 24774 6342 24832 6376
rect 24774 6308 24786 6342
rect 24820 6308 24832 6342
rect 24774 6274 24832 6308
rect 24774 6240 24786 6274
rect 24820 6240 24832 6274
rect 24774 6206 24832 6240
rect 24774 6172 24786 6206
rect 24820 6172 24832 6206
rect 24774 6138 24832 6172
rect 24774 6104 24786 6138
rect 24820 6104 24832 6138
rect 24774 6070 24832 6104
rect 24774 6036 24786 6070
rect 24820 6036 24832 6070
rect 24774 6002 24832 6036
rect 24774 5968 24786 6002
rect 24820 5968 24832 6002
rect 24774 5934 24832 5968
rect 24774 5900 24786 5934
rect 24820 5900 24832 5934
rect 24774 5866 24832 5900
rect 24774 5832 24786 5866
rect 24820 5832 24832 5866
rect 24774 5798 24832 5832
rect 23388 5730 23446 5764
rect 23388 5696 23400 5730
rect 23434 5696 23446 5730
rect 24774 5764 24786 5798
rect 24820 5764 24832 5798
rect 24774 5730 24832 5764
rect 23388 5662 23446 5696
rect 23388 5628 23400 5662
rect 23434 5628 23446 5662
rect 23388 5594 23446 5628
rect 23388 5560 23400 5594
rect 23434 5560 23446 5594
rect 23388 5526 23446 5560
rect 23388 5492 23400 5526
rect 23434 5492 23446 5526
rect 23388 5458 23446 5492
rect 23388 5424 23400 5458
rect 23434 5424 23446 5458
rect 23388 5390 23446 5424
rect 23388 5356 23400 5390
rect 23434 5356 23446 5390
rect 23388 5322 23446 5356
rect 23388 5288 23400 5322
rect 23434 5288 23446 5322
rect 23388 5254 23446 5288
rect 23388 5220 23400 5254
rect 23434 5220 23446 5254
rect 23388 5186 23446 5220
rect 23388 5152 23400 5186
rect 23434 5152 23446 5186
rect 23388 5118 23446 5152
rect 23388 5084 23400 5118
rect 23434 5084 23446 5118
rect 23388 5050 23446 5084
rect 23388 5016 23400 5050
rect 23434 5016 23446 5050
rect 23388 4982 23446 5016
rect 23388 4948 23400 4982
rect 23434 4948 23446 4982
rect 23388 4914 23446 4948
rect 23388 4880 23400 4914
rect 23434 4880 23446 4914
rect 23388 4846 23446 4880
rect 23388 4812 23400 4846
rect 23434 4812 23446 4846
rect 23388 4778 23446 4812
rect 23388 4744 23400 4778
rect 23434 4744 23446 4778
rect 23388 4710 23446 4744
rect 24774 5696 24786 5730
rect 24820 5696 24832 5730
rect 24774 5662 24832 5696
rect 24774 5628 24786 5662
rect 24820 5628 24832 5662
rect 24774 5594 24832 5628
rect 24774 5560 24786 5594
rect 24820 5560 24832 5594
rect 24774 5526 24832 5560
rect 24774 5492 24786 5526
rect 24820 5492 24832 5526
rect 24774 5458 24832 5492
rect 24774 5424 24786 5458
rect 24820 5424 24832 5458
rect 24774 5390 24832 5424
rect 24774 5356 24786 5390
rect 24820 5356 24832 5390
rect 24774 5322 24832 5356
rect 24774 5288 24786 5322
rect 24820 5288 24832 5322
rect 24774 5254 24832 5288
rect 24774 5220 24786 5254
rect 24820 5220 24832 5254
rect 24774 5186 24832 5220
rect 24774 5152 24786 5186
rect 24820 5152 24832 5186
rect 24774 5118 24832 5152
rect 24774 5084 24786 5118
rect 24820 5084 24832 5118
rect 24774 5050 24832 5084
rect 24774 5016 24786 5050
rect 24820 5016 24832 5050
rect 24774 4982 24832 5016
rect 24774 4948 24786 4982
rect 24820 4948 24832 4982
rect 24774 4914 24832 4948
rect 24774 4880 24786 4914
rect 24820 4880 24832 4914
rect 24774 4846 24832 4880
rect 24774 4812 24786 4846
rect 24820 4812 24832 4846
rect 24774 4778 24832 4812
rect 24774 4744 24786 4778
rect 24820 4744 24832 4778
rect 23388 4676 23400 4710
rect 23434 4676 23446 4710
rect 23388 4642 23446 4676
rect 24774 4710 24832 4744
rect 24774 4676 24786 4710
rect 24820 4676 24832 4710
rect 23388 4608 23400 4642
rect 23434 4608 23446 4642
rect 18738 4501 18796 4535
rect 18738 4467 18750 4501
rect 18784 4467 18796 4501
rect 18738 4384 18796 4467
rect 20064 4535 20076 4569
rect 20110 4535 20122 4569
rect 20064 4501 20122 4535
rect 20064 4467 20076 4501
rect 20110 4467 20122 4501
rect 20064 4384 20122 4467
rect 18738 4372 20122 4384
rect 18738 4338 18869 4372
rect 18903 4338 18937 4372
rect 18971 4338 19005 4372
rect 19039 4338 19073 4372
rect 19107 4338 19141 4372
rect 19175 4338 19209 4372
rect 19243 4338 19277 4372
rect 19311 4338 19345 4372
rect 19379 4338 19413 4372
rect 19447 4338 19481 4372
rect 19515 4338 19549 4372
rect 19583 4338 19617 4372
rect 19651 4338 19685 4372
rect 19719 4338 19753 4372
rect 19787 4338 19821 4372
rect 19855 4338 19889 4372
rect 19923 4338 19957 4372
rect 19991 4338 20122 4372
rect 18738 4326 20122 4338
rect 23388 4574 23446 4608
rect 23388 4540 23400 4574
rect 23434 4540 23446 4574
rect 23388 4506 23446 4540
rect 23388 4472 23400 4506
rect 23434 4472 23446 4506
rect 23388 4438 23446 4472
rect 23388 4404 23400 4438
rect 23434 4404 23446 4438
rect 23388 4370 23446 4404
rect 23388 4336 23400 4370
rect 23434 4336 23446 4370
rect 23388 4302 23446 4336
rect 23388 4268 23400 4302
rect 23434 4268 23446 4302
rect 23388 4234 23446 4268
rect 23388 4200 23400 4234
rect 23434 4200 23446 4234
rect 23388 4166 23446 4200
rect 23388 4132 23400 4166
rect 23434 4132 23446 4166
rect 23388 4098 23446 4132
rect 23388 4064 23400 4098
rect 23434 4064 23446 4098
rect 23388 4030 23446 4064
rect 23388 3996 23400 4030
rect 23434 3996 23446 4030
rect 23388 3962 23446 3996
rect 23388 3928 23400 3962
rect 23434 3928 23446 3962
rect 23388 3894 23446 3928
rect 23388 3860 23400 3894
rect 23434 3860 23446 3894
rect 23388 3826 23446 3860
rect 23388 3792 23400 3826
rect 23434 3792 23446 3826
rect 23388 3758 23446 3792
rect 23388 3724 23400 3758
rect 23434 3724 23446 3758
rect 23388 3690 23446 3724
rect 23388 3656 23400 3690
rect 23434 3656 23446 3690
rect 24774 4642 24832 4676
rect 24774 4608 24786 4642
rect 24820 4608 24832 4642
rect 24774 4574 24832 4608
rect 24774 4540 24786 4574
rect 24820 4540 24832 4574
rect 24774 4506 24832 4540
rect 24774 4472 24786 4506
rect 24820 4472 24832 4506
rect 24774 4438 24832 4472
rect 24774 4404 24786 4438
rect 24820 4404 24832 4438
rect 24774 4370 24832 4404
rect 24774 4336 24786 4370
rect 24820 4336 24832 4370
rect 24774 4302 24832 4336
rect 24774 4268 24786 4302
rect 24820 4268 24832 4302
rect 24774 4234 24832 4268
rect 24774 4200 24786 4234
rect 24820 4200 24832 4234
rect 24774 4166 24832 4200
rect 24774 4132 24786 4166
rect 24820 4132 24832 4166
rect 24774 4098 24832 4132
rect 24774 4064 24786 4098
rect 24820 4064 24832 4098
rect 24774 4030 24832 4064
rect 24774 3996 24786 4030
rect 24820 3996 24832 4030
rect 24774 3962 24832 3996
rect 24774 3928 24786 3962
rect 24820 3928 24832 3962
rect 24774 3894 24832 3928
rect 24774 3860 24786 3894
rect 24820 3860 24832 3894
rect 24774 3826 24832 3860
rect 24774 3792 24786 3826
rect 24820 3792 24832 3826
rect 24774 3758 24832 3792
rect 24774 3724 24786 3758
rect 24820 3724 24832 3758
rect 24774 3690 24832 3724
rect 23388 3622 23446 3656
rect 23388 3588 23400 3622
rect 23434 3588 23446 3622
rect 24774 3656 24786 3690
rect 24820 3656 24832 3690
rect 24774 3622 24832 3656
rect 23388 3526 23446 3588
rect 24774 3588 24786 3622
rect 24820 3588 24832 3622
rect 24774 3526 24832 3588
rect 23388 3514 24832 3526
rect 23388 3480 23515 3514
rect 23549 3480 23583 3514
rect 23617 3480 23651 3514
rect 23685 3480 23719 3514
rect 23753 3480 23787 3514
rect 23821 3480 23855 3514
rect 23889 3480 23923 3514
rect 23957 3480 23991 3514
rect 24025 3480 24059 3514
rect 24093 3480 24127 3514
rect 24161 3480 24195 3514
rect 24229 3480 24263 3514
rect 24297 3480 24331 3514
rect 24365 3480 24399 3514
rect 24433 3480 24467 3514
rect 24501 3480 24535 3514
rect 24569 3480 24603 3514
rect 24637 3480 24671 3514
rect 24705 3480 24832 3514
rect 23388 3468 24832 3480
rect 24888 8014 26332 8026
rect 24888 7980 25015 8014
rect 25049 7980 25083 8014
rect 25117 7980 25151 8014
rect 25185 7980 25219 8014
rect 25253 7980 25287 8014
rect 25321 7980 25355 8014
rect 25389 7980 25423 8014
rect 25457 7980 25491 8014
rect 25525 7980 25559 8014
rect 25593 7980 25627 8014
rect 25661 7980 25695 8014
rect 25729 7980 25763 8014
rect 25797 7980 25831 8014
rect 25865 7980 25899 8014
rect 25933 7980 25967 8014
rect 26001 7980 26035 8014
rect 26069 7980 26103 8014
rect 26137 7980 26171 8014
rect 26205 7980 26332 8014
rect 24888 7968 26332 7980
rect 24888 7906 24946 7968
rect 24888 7872 24900 7906
rect 24934 7872 24946 7906
rect 26274 7906 26332 7968
rect 24888 7838 24946 7872
rect 24888 7804 24900 7838
rect 24934 7804 24946 7838
rect 26274 7872 26286 7906
rect 26320 7872 26332 7906
rect 26274 7838 26332 7872
rect 24888 7770 24946 7804
rect 24888 7736 24900 7770
rect 24934 7736 24946 7770
rect 24888 7702 24946 7736
rect 24888 7668 24900 7702
rect 24934 7668 24946 7702
rect 24888 7634 24946 7668
rect 24888 7600 24900 7634
rect 24934 7600 24946 7634
rect 24888 7566 24946 7600
rect 24888 7532 24900 7566
rect 24934 7532 24946 7566
rect 24888 7498 24946 7532
rect 24888 7464 24900 7498
rect 24934 7464 24946 7498
rect 24888 7430 24946 7464
rect 24888 7396 24900 7430
rect 24934 7396 24946 7430
rect 24888 7362 24946 7396
rect 24888 7328 24900 7362
rect 24934 7328 24946 7362
rect 24888 7294 24946 7328
rect 24888 7260 24900 7294
rect 24934 7260 24946 7294
rect 24888 7226 24946 7260
rect 24888 7192 24900 7226
rect 24934 7192 24946 7226
rect 24888 7158 24946 7192
rect 24888 7124 24900 7158
rect 24934 7124 24946 7158
rect 24888 7090 24946 7124
rect 24888 7056 24900 7090
rect 24934 7056 24946 7090
rect 24888 7022 24946 7056
rect 24888 6988 24900 7022
rect 24934 6988 24946 7022
rect 24888 6954 24946 6988
rect 24888 6920 24900 6954
rect 24934 6920 24946 6954
rect 24888 6886 24946 6920
rect 24888 6852 24900 6886
rect 24934 6852 24946 6886
rect 24888 6818 24946 6852
rect 26274 7804 26286 7838
rect 26320 7804 26332 7838
rect 26274 7770 26332 7804
rect 26274 7736 26286 7770
rect 26320 7736 26332 7770
rect 26274 7702 26332 7736
rect 26274 7668 26286 7702
rect 26320 7668 26332 7702
rect 26274 7634 26332 7668
rect 26274 7600 26286 7634
rect 26320 7600 26332 7634
rect 26274 7566 26332 7600
rect 26274 7532 26286 7566
rect 26320 7532 26332 7566
rect 26274 7498 26332 7532
rect 26274 7464 26286 7498
rect 26320 7464 26332 7498
rect 26274 7430 26332 7464
rect 26274 7396 26286 7430
rect 26320 7396 26332 7430
rect 26274 7362 26332 7396
rect 26274 7328 26286 7362
rect 26320 7328 26332 7362
rect 26274 7294 26332 7328
rect 26274 7260 26286 7294
rect 26320 7260 26332 7294
rect 26274 7226 26332 7260
rect 26274 7192 26286 7226
rect 26320 7192 26332 7226
rect 26274 7158 26332 7192
rect 26274 7124 26286 7158
rect 26320 7124 26332 7158
rect 26274 7090 26332 7124
rect 26274 7056 26286 7090
rect 26320 7056 26332 7090
rect 26274 7022 26332 7056
rect 26274 6988 26286 7022
rect 26320 6988 26332 7022
rect 26274 6954 26332 6988
rect 26274 6920 26286 6954
rect 26320 6920 26332 6954
rect 26274 6886 26332 6920
rect 26274 6852 26286 6886
rect 26320 6852 26332 6886
rect 24888 6784 24900 6818
rect 24934 6784 24946 6818
rect 24888 6750 24946 6784
rect 26274 6818 26332 6852
rect 26274 6784 26286 6818
rect 26320 6784 26332 6818
rect 24888 6716 24900 6750
rect 24934 6716 24946 6750
rect 24888 6682 24946 6716
rect 24888 6648 24900 6682
rect 24934 6648 24946 6682
rect 24888 6614 24946 6648
rect 24888 6580 24900 6614
rect 24934 6580 24946 6614
rect 24888 6546 24946 6580
rect 24888 6512 24900 6546
rect 24934 6512 24946 6546
rect 24888 6478 24946 6512
rect 24888 6444 24900 6478
rect 24934 6444 24946 6478
rect 24888 6410 24946 6444
rect 24888 6376 24900 6410
rect 24934 6376 24946 6410
rect 24888 6342 24946 6376
rect 24888 6308 24900 6342
rect 24934 6308 24946 6342
rect 24888 6274 24946 6308
rect 24888 6240 24900 6274
rect 24934 6240 24946 6274
rect 24888 6206 24946 6240
rect 24888 6172 24900 6206
rect 24934 6172 24946 6206
rect 24888 6138 24946 6172
rect 24888 6104 24900 6138
rect 24934 6104 24946 6138
rect 24888 6070 24946 6104
rect 24888 6036 24900 6070
rect 24934 6036 24946 6070
rect 24888 6002 24946 6036
rect 24888 5968 24900 6002
rect 24934 5968 24946 6002
rect 24888 5934 24946 5968
rect 24888 5900 24900 5934
rect 24934 5900 24946 5934
rect 24888 5866 24946 5900
rect 24888 5832 24900 5866
rect 24934 5832 24946 5866
rect 24888 5798 24946 5832
rect 24888 5764 24900 5798
rect 24934 5764 24946 5798
rect 26274 6750 26332 6784
rect 26274 6716 26286 6750
rect 26320 6716 26332 6750
rect 26274 6682 26332 6716
rect 26274 6648 26286 6682
rect 26320 6648 26332 6682
rect 26274 6614 26332 6648
rect 26274 6580 26286 6614
rect 26320 6580 26332 6614
rect 26274 6546 26332 6580
rect 26274 6512 26286 6546
rect 26320 6512 26332 6546
rect 26274 6478 26332 6512
rect 26274 6444 26286 6478
rect 26320 6444 26332 6478
rect 26274 6410 26332 6444
rect 26274 6376 26286 6410
rect 26320 6376 26332 6410
rect 26274 6342 26332 6376
rect 26274 6308 26286 6342
rect 26320 6308 26332 6342
rect 26274 6274 26332 6308
rect 26274 6240 26286 6274
rect 26320 6240 26332 6274
rect 26274 6206 26332 6240
rect 26274 6172 26286 6206
rect 26320 6172 26332 6206
rect 26274 6138 26332 6172
rect 26274 6104 26286 6138
rect 26320 6104 26332 6138
rect 26274 6070 26332 6104
rect 26274 6036 26286 6070
rect 26320 6036 26332 6070
rect 26274 6002 26332 6036
rect 26274 5968 26286 6002
rect 26320 5968 26332 6002
rect 26274 5934 26332 5968
rect 26274 5900 26286 5934
rect 26320 5900 26332 5934
rect 26274 5866 26332 5900
rect 26274 5832 26286 5866
rect 26320 5832 26332 5866
rect 26274 5798 26332 5832
rect 24888 5730 24946 5764
rect 24888 5696 24900 5730
rect 24934 5696 24946 5730
rect 26274 5764 26286 5798
rect 26320 5764 26332 5798
rect 26274 5730 26332 5764
rect 24888 5662 24946 5696
rect 24888 5628 24900 5662
rect 24934 5628 24946 5662
rect 24888 5594 24946 5628
rect 24888 5560 24900 5594
rect 24934 5560 24946 5594
rect 24888 5526 24946 5560
rect 24888 5492 24900 5526
rect 24934 5492 24946 5526
rect 24888 5458 24946 5492
rect 24888 5424 24900 5458
rect 24934 5424 24946 5458
rect 24888 5390 24946 5424
rect 24888 5356 24900 5390
rect 24934 5356 24946 5390
rect 24888 5322 24946 5356
rect 24888 5288 24900 5322
rect 24934 5288 24946 5322
rect 24888 5254 24946 5288
rect 24888 5220 24900 5254
rect 24934 5220 24946 5254
rect 24888 5186 24946 5220
rect 24888 5152 24900 5186
rect 24934 5152 24946 5186
rect 24888 5118 24946 5152
rect 24888 5084 24900 5118
rect 24934 5084 24946 5118
rect 24888 5050 24946 5084
rect 24888 5016 24900 5050
rect 24934 5016 24946 5050
rect 24888 4982 24946 5016
rect 24888 4948 24900 4982
rect 24934 4948 24946 4982
rect 24888 4914 24946 4948
rect 24888 4880 24900 4914
rect 24934 4880 24946 4914
rect 24888 4846 24946 4880
rect 24888 4812 24900 4846
rect 24934 4812 24946 4846
rect 24888 4778 24946 4812
rect 24888 4744 24900 4778
rect 24934 4744 24946 4778
rect 24888 4710 24946 4744
rect 26274 5696 26286 5730
rect 26320 5696 26332 5730
rect 26274 5662 26332 5696
rect 26274 5628 26286 5662
rect 26320 5628 26332 5662
rect 26274 5594 26332 5628
rect 26274 5560 26286 5594
rect 26320 5560 26332 5594
rect 26274 5526 26332 5560
rect 26274 5492 26286 5526
rect 26320 5492 26332 5526
rect 26274 5458 26332 5492
rect 26274 5424 26286 5458
rect 26320 5424 26332 5458
rect 26274 5390 26332 5424
rect 26274 5356 26286 5390
rect 26320 5356 26332 5390
rect 26274 5322 26332 5356
rect 26274 5288 26286 5322
rect 26320 5288 26332 5322
rect 26274 5254 26332 5288
rect 26274 5220 26286 5254
rect 26320 5220 26332 5254
rect 26274 5186 26332 5220
rect 26274 5152 26286 5186
rect 26320 5152 26332 5186
rect 26274 5118 26332 5152
rect 26274 5084 26286 5118
rect 26320 5084 26332 5118
rect 26274 5050 26332 5084
rect 26274 5016 26286 5050
rect 26320 5016 26332 5050
rect 26274 4982 26332 5016
rect 26274 4948 26286 4982
rect 26320 4948 26332 4982
rect 26274 4914 26332 4948
rect 26274 4880 26286 4914
rect 26320 4880 26332 4914
rect 26274 4846 26332 4880
rect 26274 4812 26286 4846
rect 26320 4812 26332 4846
rect 26274 4778 26332 4812
rect 26274 4744 26286 4778
rect 26320 4744 26332 4778
rect 24888 4676 24900 4710
rect 24934 4676 24946 4710
rect 24888 4642 24946 4676
rect 26274 4710 26332 4744
rect 26274 4676 26286 4710
rect 26320 4676 26332 4710
rect 24888 4608 24900 4642
rect 24934 4608 24946 4642
rect 24888 4574 24946 4608
rect 24888 4540 24900 4574
rect 24934 4540 24946 4574
rect 24888 4506 24946 4540
rect 24888 4472 24900 4506
rect 24934 4472 24946 4506
rect 24888 4438 24946 4472
rect 24888 4404 24900 4438
rect 24934 4404 24946 4438
rect 24888 4370 24946 4404
rect 24888 4336 24900 4370
rect 24934 4336 24946 4370
rect 24888 4302 24946 4336
rect 24888 4268 24900 4302
rect 24934 4268 24946 4302
rect 24888 4234 24946 4268
rect 24888 4200 24900 4234
rect 24934 4200 24946 4234
rect 24888 4166 24946 4200
rect 24888 4132 24900 4166
rect 24934 4132 24946 4166
rect 24888 4098 24946 4132
rect 24888 4064 24900 4098
rect 24934 4064 24946 4098
rect 24888 4030 24946 4064
rect 24888 3996 24900 4030
rect 24934 3996 24946 4030
rect 24888 3962 24946 3996
rect 24888 3928 24900 3962
rect 24934 3928 24946 3962
rect 24888 3894 24946 3928
rect 24888 3860 24900 3894
rect 24934 3860 24946 3894
rect 24888 3826 24946 3860
rect 24888 3792 24900 3826
rect 24934 3792 24946 3826
rect 24888 3758 24946 3792
rect 24888 3724 24900 3758
rect 24934 3724 24946 3758
rect 24888 3690 24946 3724
rect 24888 3656 24900 3690
rect 24934 3656 24946 3690
rect 26274 4642 26332 4676
rect 26274 4608 26286 4642
rect 26320 4608 26332 4642
rect 26274 4574 26332 4608
rect 26274 4540 26286 4574
rect 26320 4540 26332 4574
rect 26274 4506 26332 4540
rect 26274 4472 26286 4506
rect 26320 4472 26332 4506
rect 26274 4438 26332 4472
rect 26274 4404 26286 4438
rect 26320 4404 26332 4438
rect 26274 4370 26332 4404
rect 26274 4336 26286 4370
rect 26320 4336 26332 4370
rect 26274 4302 26332 4336
rect 26274 4268 26286 4302
rect 26320 4268 26332 4302
rect 26274 4234 26332 4268
rect 26274 4200 26286 4234
rect 26320 4200 26332 4234
rect 26274 4166 26332 4200
rect 26274 4132 26286 4166
rect 26320 4132 26332 4166
rect 26274 4098 26332 4132
rect 26274 4064 26286 4098
rect 26320 4064 26332 4098
rect 26274 4030 26332 4064
rect 26274 3996 26286 4030
rect 26320 3996 26332 4030
rect 26274 3962 26332 3996
rect 26274 3928 26286 3962
rect 26320 3928 26332 3962
rect 26274 3894 26332 3928
rect 26274 3860 26286 3894
rect 26320 3860 26332 3894
rect 26274 3826 26332 3860
rect 26274 3792 26286 3826
rect 26320 3792 26332 3826
rect 26274 3758 26332 3792
rect 26274 3724 26286 3758
rect 26320 3724 26332 3758
rect 26274 3690 26332 3724
rect 24888 3622 24946 3656
rect 24888 3588 24900 3622
rect 24934 3588 24946 3622
rect 26274 3656 26286 3690
rect 26320 3656 26332 3690
rect 26274 3622 26332 3656
rect 24888 3526 24946 3588
rect 26274 3588 26286 3622
rect 26320 3588 26332 3622
rect 26274 3526 26332 3588
rect 24888 3514 26332 3526
rect 24888 3480 25015 3514
rect 25049 3480 25083 3514
rect 25117 3480 25151 3514
rect 25185 3480 25219 3514
rect 25253 3480 25287 3514
rect 25321 3480 25355 3514
rect 25389 3480 25423 3514
rect 25457 3480 25491 3514
rect 25525 3480 25559 3514
rect 25593 3480 25627 3514
rect 25661 3480 25695 3514
rect 25729 3480 25763 3514
rect 25797 3480 25831 3514
rect 25865 3480 25899 3514
rect 25933 3480 25967 3514
rect 26001 3480 26035 3514
rect 26069 3480 26103 3514
rect 26137 3480 26171 3514
rect 26205 3480 26332 3514
rect 24888 3468 26332 3480
rect 36473 12315 42317 12358
rect 36473 12281 36760 12315
rect 36794 12281 36828 12315
rect 36862 12281 36896 12315
rect 36930 12281 36964 12315
rect 36998 12281 37032 12315
rect 37066 12281 37100 12315
rect 37134 12281 37168 12315
rect 37202 12281 37236 12315
rect 37270 12281 37304 12315
rect 37338 12281 37372 12315
rect 37406 12281 37440 12315
rect 37474 12281 37508 12315
rect 37542 12281 37576 12315
rect 37610 12281 37644 12315
rect 37678 12281 37712 12315
rect 37746 12281 37780 12315
rect 37814 12281 37848 12315
rect 37882 12281 37916 12315
rect 37950 12281 37984 12315
rect 38018 12281 38052 12315
rect 38086 12281 38120 12315
rect 38154 12281 38188 12315
rect 38222 12281 38256 12315
rect 38290 12281 38324 12315
rect 38358 12281 38392 12315
rect 38426 12281 38460 12315
rect 38494 12281 38528 12315
rect 38562 12281 38596 12315
rect 38630 12281 38664 12315
rect 38698 12281 38732 12315
rect 38766 12281 38800 12315
rect 38834 12281 38868 12315
rect 38902 12281 38936 12315
rect 38970 12281 39004 12315
rect 39038 12281 39072 12315
rect 39106 12281 39140 12315
rect 39174 12281 39208 12315
rect 39242 12281 39276 12315
rect 39310 12281 39344 12315
rect 39378 12281 39412 12315
rect 39446 12281 39480 12315
rect 39514 12281 39548 12315
rect 39582 12281 39616 12315
rect 39650 12281 39684 12315
rect 39718 12281 39752 12315
rect 39786 12281 39820 12315
rect 39854 12281 39888 12315
rect 39922 12281 39956 12315
rect 39990 12281 40024 12315
rect 40058 12281 40092 12315
rect 40126 12281 40160 12315
rect 40194 12281 40228 12315
rect 40262 12281 40296 12315
rect 40330 12281 40364 12315
rect 40398 12281 40432 12315
rect 40466 12281 40500 12315
rect 40534 12281 40568 12315
rect 40602 12281 40636 12315
rect 40670 12281 40704 12315
rect 40738 12281 40772 12315
rect 40806 12281 40840 12315
rect 40874 12281 40908 12315
rect 40942 12281 40976 12315
rect 41010 12281 41044 12315
rect 41078 12281 41112 12315
rect 41146 12281 41180 12315
rect 41214 12281 41248 12315
rect 41282 12281 41316 12315
rect 41350 12281 41384 12315
rect 41418 12281 41452 12315
rect 41486 12281 41520 12315
rect 41554 12281 41588 12315
rect 41622 12281 41656 12315
rect 41690 12281 41724 12315
rect 41758 12281 41792 12315
rect 41826 12281 41860 12315
rect 41894 12281 41928 12315
rect 41962 12281 41996 12315
rect 42030 12281 42317 12315
rect 36473 12240 42317 12281
rect 36473 12125 36587 12240
rect 36473 12091 36511 12125
rect 36545 12091 36587 12125
rect 36473 12057 36587 12091
rect 36473 12023 36511 12057
rect 36545 12023 36587 12057
rect 36473 11989 36587 12023
rect 42190 12085 42317 12240
rect 42190 12051 42237 12085
rect 42271 12051 42317 12085
rect 42190 12017 42317 12051
rect 36473 11955 36511 11989
rect 36545 11955 36587 11989
rect 36473 11921 36587 11955
rect 36473 11887 36511 11921
rect 36545 11887 36587 11921
rect 42190 11983 42237 12017
rect 42271 11983 42317 12017
rect 42190 11949 42317 11983
rect 42190 11915 42237 11949
rect 42271 11915 42317 11949
rect 36473 11853 36587 11887
rect 36473 11819 36511 11853
rect 36545 11819 36587 11853
rect 36473 11785 36587 11819
rect 36473 11751 36511 11785
rect 36545 11751 36587 11785
rect 36473 11717 36587 11751
rect 36473 11683 36511 11717
rect 36545 11683 36587 11717
rect 36473 11649 36587 11683
rect 36473 11615 36511 11649
rect 36545 11615 36587 11649
rect 36473 11581 36587 11615
rect 36473 11547 36511 11581
rect 36545 11547 36587 11581
rect 36473 11513 36587 11547
rect 36473 11479 36511 11513
rect 36545 11479 36587 11513
rect 36473 11445 36587 11479
rect 36473 11411 36511 11445
rect 36545 11411 36587 11445
rect 36473 11377 36587 11411
rect 36473 11343 36511 11377
rect 36545 11343 36587 11377
rect 36473 11309 36587 11343
rect 36473 11275 36511 11309
rect 36545 11275 36587 11309
rect 36473 11241 36587 11275
rect 36473 11207 36511 11241
rect 36545 11207 36587 11241
rect 36473 11173 36587 11207
rect 36473 11139 36511 11173
rect 36545 11139 36587 11173
rect 36473 11105 36587 11139
rect 36473 11071 36511 11105
rect 36545 11071 36587 11105
rect 36473 11037 36587 11071
rect 36473 11003 36511 11037
rect 36545 11003 36587 11037
rect 36473 10969 36587 11003
rect 36473 10935 36511 10969
rect 36545 10935 36587 10969
rect 36473 10901 36587 10935
rect 42190 11881 42317 11915
rect 42190 11847 42237 11881
rect 42271 11847 42317 11881
rect 42190 11813 42317 11847
rect 42190 11779 42237 11813
rect 42271 11779 42317 11813
rect 42190 11745 42317 11779
rect 42190 11711 42237 11745
rect 42271 11711 42317 11745
rect 42190 11677 42317 11711
rect 42190 11643 42237 11677
rect 42271 11643 42317 11677
rect 42190 11609 42317 11643
rect 42190 11575 42237 11609
rect 42271 11575 42317 11609
rect 42190 11541 42317 11575
rect 42190 11507 42237 11541
rect 42271 11507 42317 11541
rect 42190 11473 42317 11507
rect 42190 11439 42237 11473
rect 42271 11439 42317 11473
rect 42190 11405 42317 11439
rect 42190 11371 42237 11405
rect 42271 11371 42317 11405
rect 42190 11337 42317 11371
rect 42190 11303 42237 11337
rect 42271 11303 42317 11337
rect 42190 11269 42317 11303
rect 42190 11235 42237 11269
rect 42271 11235 42317 11269
rect 42190 11201 42317 11235
rect 42190 11167 42237 11201
rect 42271 11167 42317 11201
rect 42190 11133 42317 11167
rect 42190 11099 42237 11133
rect 42271 11099 42317 11133
rect 42190 11065 42317 11099
rect 42190 11031 42237 11065
rect 42271 11031 42317 11065
rect 42190 10997 42317 11031
rect 42190 10963 42237 10997
rect 42271 10963 42317 10997
rect 42190 10929 42317 10963
rect 36473 10867 36511 10901
rect 36545 10867 36587 10901
rect 36473 10833 36587 10867
rect 36473 10799 36511 10833
rect 36545 10799 36587 10833
rect 42190 10895 42237 10929
rect 42271 10895 42317 10929
rect 42190 10861 42317 10895
rect 42190 10827 42237 10861
rect 42271 10827 42317 10861
rect 36473 10765 36587 10799
rect 36473 10731 36511 10765
rect 36545 10731 36587 10765
rect 36473 10697 36587 10731
rect 36473 10663 36511 10697
rect 36545 10663 36587 10697
rect 36473 10629 36587 10663
rect 42190 10793 42317 10827
rect 42190 10759 42237 10793
rect 42271 10759 42317 10793
rect 42190 10725 42317 10759
rect 42190 10691 42237 10725
rect 42271 10691 42317 10725
rect 42190 10657 42317 10691
rect 36473 10595 36511 10629
rect 36545 10595 36587 10629
rect 36473 10561 36587 10595
rect 36473 10527 36511 10561
rect 36545 10527 36587 10561
rect 42190 10623 42237 10657
rect 42271 10623 42317 10657
rect 42190 10589 42317 10623
rect 42190 10555 42237 10589
rect 42271 10555 42317 10589
rect 36473 10493 36587 10527
rect 36473 10459 36511 10493
rect 36545 10459 36587 10493
rect 36473 10425 36587 10459
rect 36473 10391 36511 10425
rect 36545 10391 36587 10425
rect 36473 10357 36587 10391
rect 36473 10323 36511 10357
rect 36545 10323 36587 10357
rect 36473 10289 36587 10323
rect 36473 10255 36511 10289
rect 36545 10255 36587 10289
rect 36473 10221 36587 10255
rect 36473 10187 36511 10221
rect 36545 10187 36587 10221
rect 36473 10153 36587 10187
rect 36473 10119 36511 10153
rect 36545 10119 36587 10153
rect 36473 10085 36587 10119
rect 36473 10051 36511 10085
rect 36545 10051 36587 10085
rect 36473 10017 36587 10051
rect 36473 9983 36511 10017
rect 36545 9983 36587 10017
rect 36473 9949 36587 9983
rect 36473 9915 36511 9949
rect 36545 9915 36587 9949
rect 36473 9881 36587 9915
rect 36473 9847 36511 9881
rect 36545 9847 36587 9881
rect 36473 9813 36587 9847
rect 36473 9779 36511 9813
rect 36545 9779 36587 9813
rect 36473 9745 36587 9779
rect 36473 9711 36511 9745
rect 36545 9711 36587 9745
rect 36473 9677 36587 9711
rect 36473 9643 36511 9677
rect 36545 9643 36587 9677
rect 36473 9609 36587 9643
rect 36473 9575 36511 9609
rect 36545 9575 36587 9609
rect 36473 9541 36587 9575
rect 42190 10521 42317 10555
rect 42190 10487 42237 10521
rect 42271 10487 42317 10521
rect 42190 10453 42317 10487
rect 42190 10419 42237 10453
rect 42271 10419 42317 10453
rect 42190 10385 42317 10419
rect 42190 10351 42237 10385
rect 42271 10351 42317 10385
rect 42190 10317 42317 10351
rect 42190 10283 42237 10317
rect 42271 10283 42317 10317
rect 42190 10249 42317 10283
rect 42190 10215 42237 10249
rect 42271 10215 42317 10249
rect 42190 10181 42317 10215
rect 42190 10147 42237 10181
rect 42271 10147 42317 10181
rect 42190 10113 42317 10147
rect 42190 10079 42237 10113
rect 42271 10079 42317 10113
rect 42190 10045 42317 10079
rect 42190 10011 42237 10045
rect 42271 10011 42317 10045
rect 42190 9977 42317 10011
rect 42190 9943 42237 9977
rect 42271 9943 42317 9977
rect 42190 9909 42317 9943
rect 42190 9875 42237 9909
rect 42271 9875 42317 9909
rect 42190 9841 42317 9875
rect 42190 9807 42237 9841
rect 42271 9807 42317 9841
rect 42190 9773 42317 9807
rect 42190 9739 42237 9773
rect 42271 9739 42317 9773
rect 42190 9705 42317 9739
rect 42190 9671 42237 9705
rect 42271 9671 42317 9705
rect 42190 9637 42317 9671
rect 42190 9603 42237 9637
rect 42271 9603 42317 9637
rect 42190 9569 42317 9603
rect 36473 9507 36511 9541
rect 36545 9507 36587 9541
rect 36473 9473 36587 9507
rect 36473 9439 36511 9473
rect 36545 9439 36587 9473
rect 42190 9535 42237 9569
rect 42271 9535 42317 9569
rect 42190 9501 42317 9535
rect 42190 9467 42237 9501
rect 42271 9467 42317 9501
rect 36473 9405 36587 9439
rect 36473 9371 36511 9405
rect 36545 9371 36587 9405
rect 36473 9190 36587 9371
rect 42190 9433 42317 9467
rect 42190 9399 42237 9433
rect 42271 9399 42317 9433
rect 42190 9365 42317 9399
rect 42190 9331 42237 9365
rect 42271 9331 42317 9365
rect 42190 9190 42317 9331
rect 36473 9149 42317 9190
rect 36473 9115 36779 9149
rect 36813 9115 36847 9149
rect 36881 9115 36915 9149
rect 36949 9115 36983 9149
rect 37017 9115 37051 9149
rect 37085 9115 37119 9149
rect 37153 9115 37187 9149
rect 37221 9115 37255 9149
rect 37289 9115 37323 9149
rect 37357 9115 37391 9149
rect 37425 9115 37459 9149
rect 37493 9115 37527 9149
rect 37561 9115 37595 9149
rect 37629 9115 37663 9149
rect 37697 9115 37731 9149
rect 37765 9115 37799 9149
rect 37833 9115 37867 9149
rect 37901 9115 37935 9149
rect 37969 9115 38003 9149
rect 38037 9115 38071 9149
rect 38105 9115 38139 9149
rect 38173 9115 38207 9149
rect 38241 9115 38275 9149
rect 38309 9115 38343 9149
rect 38377 9115 38411 9149
rect 38445 9115 38479 9149
rect 38513 9115 38547 9149
rect 38581 9115 38615 9149
rect 38649 9115 38683 9149
rect 38717 9115 38751 9149
rect 38785 9115 38819 9149
rect 38853 9115 38887 9149
rect 38921 9115 38955 9149
rect 38989 9115 39023 9149
rect 39057 9115 39091 9149
rect 39125 9115 39159 9149
rect 39193 9115 39227 9149
rect 39261 9115 39295 9149
rect 39329 9115 39363 9149
rect 39397 9115 39431 9149
rect 39465 9115 39499 9149
rect 39533 9115 39567 9149
rect 39601 9115 39635 9149
rect 39669 9115 39703 9149
rect 39737 9115 39771 9149
rect 39805 9115 39839 9149
rect 39873 9115 39907 9149
rect 39941 9115 39975 9149
rect 40009 9115 40043 9149
rect 40077 9115 40111 9149
rect 40145 9115 40179 9149
rect 40213 9115 40247 9149
rect 40281 9115 40315 9149
rect 40349 9115 40383 9149
rect 40417 9115 40451 9149
rect 40485 9115 40519 9149
rect 40553 9115 40587 9149
rect 40621 9115 40655 9149
rect 40689 9115 40723 9149
rect 40757 9115 40791 9149
rect 40825 9115 40859 9149
rect 40893 9115 40927 9149
rect 40961 9115 40995 9149
rect 41029 9115 41063 9149
rect 41097 9115 41131 9149
rect 41165 9115 41199 9149
rect 41233 9115 41267 9149
rect 41301 9115 41335 9149
rect 41369 9115 41403 9149
rect 41437 9115 41471 9149
rect 41505 9115 41539 9149
rect 41573 9115 41607 9149
rect 41641 9115 41675 9149
rect 41709 9115 41743 9149
rect 41777 9115 41811 9149
rect 41845 9115 41879 9149
rect 41913 9115 41947 9149
rect 41981 9115 42015 9149
rect 42049 9115 42317 9149
rect 36473 9076 42317 9115
rect 37600 8609 42194 8632
rect 37600 8575 37843 8609
rect 37877 8575 37911 8609
rect 37945 8575 37979 8609
rect 38013 8575 38047 8609
rect 38081 8575 38115 8609
rect 38149 8575 38183 8609
rect 38217 8575 38251 8609
rect 38285 8575 38319 8609
rect 38353 8575 38387 8609
rect 38421 8575 38455 8609
rect 38489 8575 38523 8609
rect 38557 8575 38591 8609
rect 38625 8575 38659 8609
rect 38693 8575 38727 8609
rect 38761 8575 38795 8609
rect 38829 8575 38863 8609
rect 38897 8575 38931 8609
rect 38965 8575 38999 8609
rect 39033 8575 39067 8609
rect 39101 8575 39135 8609
rect 39169 8575 39203 8609
rect 39237 8575 39271 8609
rect 39305 8575 39339 8609
rect 39373 8575 39407 8609
rect 39441 8575 39475 8609
rect 39509 8575 39543 8609
rect 39577 8575 39611 8609
rect 39645 8575 39679 8609
rect 39713 8575 39747 8609
rect 39781 8575 39815 8609
rect 39849 8575 39883 8609
rect 39917 8575 39951 8609
rect 39985 8575 40019 8609
rect 40053 8575 40087 8609
rect 40121 8575 40155 8609
rect 40189 8575 40223 8609
rect 40257 8575 40291 8609
rect 40325 8575 40359 8609
rect 40393 8575 40427 8609
rect 40461 8575 40495 8609
rect 40529 8575 40563 8609
rect 40597 8575 40631 8609
rect 40665 8575 40699 8609
rect 40733 8575 40767 8609
rect 40801 8575 40835 8609
rect 40869 8575 40903 8609
rect 40937 8575 40971 8609
rect 41005 8575 41039 8609
rect 41073 8575 41107 8609
rect 41141 8575 41175 8609
rect 41209 8575 41243 8609
rect 41277 8575 41311 8609
rect 41345 8575 41379 8609
rect 41413 8575 41447 8609
rect 41481 8575 41515 8609
rect 41549 8575 41583 8609
rect 41617 8575 41651 8609
rect 41685 8575 41719 8609
rect 41753 8575 41787 8609
rect 41821 8575 41855 8609
rect 41889 8575 41923 8609
rect 41957 8575 41991 8609
rect 42025 8575 42194 8609
rect 37600 8556 42194 8575
rect 37600 8432 37682 8556
rect 37600 8398 37624 8432
rect 37658 8398 37682 8432
rect 37600 8364 37682 8398
rect 42112 8444 42194 8556
rect 42112 8410 42136 8444
rect 42170 8410 42194 8444
rect 42112 8376 42194 8410
rect 37600 8330 37624 8364
rect 37658 8330 37682 8364
rect 37600 8296 37682 8330
rect 37600 8262 37624 8296
rect 37658 8262 37682 8296
rect 42112 8342 42136 8376
rect 42170 8342 42194 8376
rect 42112 8308 42194 8342
rect 37600 8228 37682 8262
rect 37600 8194 37624 8228
rect 37658 8194 37682 8228
rect 37600 8160 37682 8194
rect 37600 8126 37624 8160
rect 37658 8126 37682 8160
rect 37600 8092 37682 8126
rect 37600 8058 37624 8092
rect 37658 8058 37682 8092
rect 37600 8024 37682 8058
rect 37600 7990 37624 8024
rect 37658 7990 37682 8024
rect 37600 7956 37682 7990
rect 37600 7922 37624 7956
rect 37658 7922 37682 7956
rect 37600 7888 37682 7922
rect 37600 7854 37624 7888
rect 37658 7854 37682 7888
rect 37600 7820 37682 7854
rect 37600 7786 37624 7820
rect 37658 7786 37682 7820
rect 37600 7752 37682 7786
rect 37600 7718 37624 7752
rect 37658 7718 37682 7752
rect 37600 7684 37682 7718
rect 37600 7650 37624 7684
rect 37658 7650 37682 7684
rect 37600 7616 37682 7650
rect 37600 7582 37624 7616
rect 37658 7582 37682 7616
rect 37600 7548 37682 7582
rect 37600 7514 37624 7548
rect 37658 7514 37682 7548
rect 37600 7480 37682 7514
rect 37600 7446 37624 7480
rect 37658 7446 37682 7480
rect 37600 7412 37682 7446
rect 37600 7378 37624 7412
rect 37658 7378 37682 7412
rect 37600 7344 37682 7378
rect 37600 7310 37624 7344
rect 37658 7310 37682 7344
rect 37600 7276 37682 7310
rect 37600 7242 37624 7276
rect 37658 7242 37682 7276
rect 37600 7208 37682 7242
rect 37600 7174 37624 7208
rect 37658 7174 37682 7208
rect 37600 7140 37682 7174
rect 37600 7106 37624 7140
rect 37658 7106 37682 7140
rect 37600 7072 37682 7106
rect 37600 7038 37624 7072
rect 37658 7038 37682 7072
rect 37600 7004 37682 7038
rect 37600 6970 37624 7004
rect 37658 6970 37682 7004
rect 37600 6936 37682 6970
rect 37600 6902 37624 6936
rect 37658 6902 37682 6936
rect 37600 6868 37682 6902
rect 37600 6834 37624 6868
rect 37658 6834 37682 6868
rect 37600 6800 37682 6834
rect 37600 6766 37624 6800
rect 37658 6766 37682 6800
rect 37600 6732 37682 6766
rect 37600 6698 37624 6732
rect 37658 6698 37682 6732
rect 37600 6664 37682 6698
rect 37600 6630 37624 6664
rect 37658 6630 37682 6664
rect 37600 6596 37682 6630
rect 37600 6562 37624 6596
rect 37658 6562 37682 6596
rect 37600 6528 37682 6562
rect 37600 6494 37624 6528
rect 37658 6494 37682 6528
rect 37600 6460 37682 6494
rect 37600 6426 37624 6460
rect 37658 6426 37682 6460
rect 37600 6392 37682 6426
rect 37600 6358 37624 6392
rect 37658 6358 37682 6392
rect 37600 6324 37682 6358
rect 37600 6290 37624 6324
rect 37658 6290 37682 6324
rect 37600 6256 37682 6290
rect 42112 8274 42136 8308
rect 42170 8274 42194 8308
rect 42112 8240 42194 8274
rect 42112 8206 42136 8240
rect 42170 8206 42194 8240
rect 42112 8172 42194 8206
rect 42112 8138 42136 8172
rect 42170 8138 42194 8172
rect 42112 8104 42194 8138
rect 42112 8070 42136 8104
rect 42170 8070 42194 8104
rect 42112 8036 42194 8070
rect 42112 8002 42136 8036
rect 42170 8002 42194 8036
rect 42112 7968 42194 8002
rect 42112 7934 42136 7968
rect 42170 7934 42194 7968
rect 42112 7900 42194 7934
rect 42112 7866 42136 7900
rect 42170 7866 42194 7900
rect 42112 7832 42194 7866
rect 42112 7798 42136 7832
rect 42170 7798 42194 7832
rect 42112 7764 42194 7798
rect 42112 7730 42136 7764
rect 42170 7730 42194 7764
rect 42112 7696 42194 7730
rect 42112 7662 42136 7696
rect 42170 7662 42194 7696
rect 42112 7628 42194 7662
rect 42112 7594 42136 7628
rect 42170 7594 42194 7628
rect 42112 7560 42194 7594
rect 42112 7526 42136 7560
rect 42170 7526 42194 7560
rect 42112 7492 42194 7526
rect 42112 7458 42136 7492
rect 42170 7458 42194 7492
rect 42112 7424 42194 7458
rect 42112 7390 42136 7424
rect 42170 7390 42194 7424
rect 42112 7356 42194 7390
rect 42112 7322 42136 7356
rect 42170 7322 42194 7356
rect 42112 7288 42194 7322
rect 42112 7254 42136 7288
rect 42170 7254 42194 7288
rect 42112 7220 42194 7254
rect 42112 7186 42136 7220
rect 42170 7186 42194 7220
rect 42112 7152 42194 7186
rect 42112 7118 42136 7152
rect 42170 7118 42194 7152
rect 42112 7084 42194 7118
rect 42112 7050 42136 7084
rect 42170 7050 42194 7084
rect 42112 7016 42194 7050
rect 42112 6982 42136 7016
rect 42170 6982 42194 7016
rect 42112 6948 42194 6982
rect 42112 6914 42136 6948
rect 42170 6914 42194 6948
rect 42112 6880 42194 6914
rect 42112 6846 42136 6880
rect 42170 6846 42194 6880
rect 42112 6812 42194 6846
rect 42112 6778 42136 6812
rect 42170 6778 42194 6812
rect 42112 6744 42194 6778
rect 42112 6710 42136 6744
rect 42170 6710 42194 6744
rect 42112 6676 42194 6710
rect 42112 6642 42136 6676
rect 42170 6642 42194 6676
rect 42112 6608 42194 6642
rect 42112 6574 42136 6608
rect 42170 6574 42194 6608
rect 42112 6540 42194 6574
rect 42112 6506 42136 6540
rect 42170 6506 42194 6540
rect 42112 6472 42194 6506
rect 42112 6438 42136 6472
rect 42170 6438 42194 6472
rect 42112 6404 42194 6438
rect 42112 6370 42136 6404
rect 42170 6370 42194 6404
rect 42112 6336 42194 6370
rect 42112 6302 42136 6336
rect 42170 6302 42194 6336
rect 37600 6222 37624 6256
rect 37658 6222 37682 6256
rect 37600 6188 37682 6222
rect 42112 6268 42194 6302
rect 42112 6234 42136 6268
rect 42170 6234 42194 6268
rect 42112 6200 42194 6234
rect 37600 6154 37624 6188
rect 37658 6154 37682 6188
rect 37600 6050 37682 6154
rect 42112 6166 42136 6200
rect 42170 6166 42194 6200
rect 42112 6050 42194 6166
rect 37600 6029 42194 6050
rect 37600 5995 37819 6029
rect 37853 5995 37887 6029
rect 37921 5995 37955 6029
rect 37989 5995 38023 6029
rect 38057 5995 38091 6029
rect 38125 5995 38159 6029
rect 38193 5995 38227 6029
rect 38261 5995 38295 6029
rect 38329 5995 38363 6029
rect 38397 5995 38431 6029
rect 38465 5995 38499 6029
rect 38533 5995 38567 6029
rect 38601 5995 38635 6029
rect 38669 5995 38703 6029
rect 38737 5995 38771 6029
rect 38805 5995 38839 6029
rect 38873 5995 38907 6029
rect 38941 5995 38975 6029
rect 39009 5995 39043 6029
rect 39077 5995 39111 6029
rect 39145 5995 39179 6029
rect 39213 5995 39247 6029
rect 39281 5995 39315 6029
rect 39349 5995 39383 6029
rect 39417 5995 39451 6029
rect 39485 5995 39519 6029
rect 39553 5995 39587 6029
rect 39621 5995 39655 6029
rect 39689 5995 39723 6029
rect 39757 5995 39791 6029
rect 39825 5995 39859 6029
rect 39893 5995 39927 6029
rect 39961 5995 39995 6029
rect 40029 5995 40063 6029
rect 40097 5995 40131 6029
rect 40165 5995 40199 6029
rect 40233 5995 40267 6029
rect 40301 5995 40335 6029
rect 40369 5995 40403 6029
rect 40437 5995 40471 6029
rect 40505 5995 40539 6029
rect 40573 5995 40607 6029
rect 40641 5995 40675 6029
rect 40709 5995 40743 6029
rect 40777 5995 40811 6029
rect 40845 5995 40879 6029
rect 40913 5995 40947 6029
rect 40981 5995 41015 6029
rect 41049 5995 41083 6029
rect 41117 5995 41151 6029
rect 41185 5995 41219 6029
rect 41253 5995 41287 6029
rect 41321 5995 41355 6029
rect 41389 5995 41423 6029
rect 41457 5995 41491 6029
rect 41525 5995 41559 6029
rect 41593 5995 41627 6029
rect 41661 5995 41695 6029
rect 41729 5995 41763 6029
rect 41797 5995 41831 6029
rect 41865 5995 41899 6029
rect 41933 5995 41967 6029
rect 42001 5995 42194 6029
rect 37600 5976 42194 5995
<< mvnsubdiff >>
rect 42466 19062 45372 19074
rect 42466 19028 42576 19062
rect 42610 19028 42644 19062
rect 42678 19028 42712 19062
rect 42746 19028 42780 19062
rect 42814 19028 42848 19062
rect 42882 19028 42916 19062
rect 42950 19028 42984 19062
rect 43018 19028 43052 19062
rect 43086 19028 43120 19062
rect 43154 19028 43188 19062
rect 43222 19028 43256 19062
rect 43290 19028 43324 19062
rect 43358 19028 43392 19062
rect 43426 19028 43460 19062
rect 43494 19028 43528 19062
rect 43562 19028 43596 19062
rect 43630 19028 43664 19062
rect 43698 19028 43732 19062
rect 43766 19028 43800 19062
rect 43834 19028 43868 19062
rect 43902 19028 43936 19062
rect 43970 19028 44004 19062
rect 44038 19028 44072 19062
rect 44106 19028 44140 19062
rect 44174 19028 44208 19062
rect 44242 19028 44276 19062
rect 44310 19028 44344 19062
rect 44378 19028 44412 19062
rect 44446 19028 44480 19062
rect 44514 19028 44548 19062
rect 44582 19028 44616 19062
rect 44650 19028 44684 19062
rect 44718 19028 44752 19062
rect 44786 19028 44820 19062
rect 44854 19028 44888 19062
rect 44922 19028 44956 19062
rect 44990 19028 45024 19062
rect 45058 19028 45092 19062
rect 45126 19028 45160 19062
rect 45194 19028 45228 19062
rect 45262 19028 45372 19062
rect 42466 19016 45372 19028
rect 23030 18966 24414 18978
rect 23030 18932 23161 18966
rect 23195 18932 23229 18966
rect 23263 18932 23297 18966
rect 23331 18932 23365 18966
rect 23399 18932 23433 18966
rect 23467 18932 23501 18966
rect 23535 18932 23569 18966
rect 23603 18932 23637 18966
rect 23671 18932 23705 18966
rect 23739 18932 23773 18966
rect 23807 18932 23841 18966
rect 23875 18932 23909 18966
rect 23943 18932 23977 18966
rect 24011 18932 24045 18966
rect 24079 18932 24113 18966
rect 24147 18932 24181 18966
rect 24215 18932 24249 18966
rect 24283 18932 24414 18966
rect 23030 18920 24414 18932
rect 23030 18842 23088 18920
rect 23030 18808 23042 18842
rect 23076 18808 23088 18842
rect 23030 18774 23088 18808
rect 23030 18740 23042 18774
rect 23076 18740 23088 18774
rect 24356 18842 24414 18920
rect 24356 18808 24368 18842
rect 24402 18808 24414 18842
rect 24356 18774 24414 18808
rect 23030 18706 23088 18740
rect 23030 18672 23042 18706
rect 23076 18672 23088 18706
rect 23030 18638 23088 18672
rect 23030 18604 23042 18638
rect 23076 18604 23088 18638
rect 23030 18570 23088 18604
rect 23030 18536 23042 18570
rect 23076 18536 23088 18570
rect 23030 18502 23088 18536
rect 23030 18468 23042 18502
rect 23076 18468 23088 18502
rect 23030 18434 23088 18468
rect 23030 18400 23042 18434
rect 23076 18400 23088 18434
rect 23030 18366 23088 18400
rect 23030 18332 23042 18366
rect 23076 18332 23088 18366
rect -3126 18312 -220 18324
rect -3126 18278 -3016 18312
rect -2982 18278 -2948 18312
rect -2914 18278 -2880 18312
rect -2846 18278 -2812 18312
rect -2778 18278 -2744 18312
rect -2710 18278 -2676 18312
rect -2642 18278 -2608 18312
rect -2574 18278 -2540 18312
rect -2506 18278 -2472 18312
rect -2438 18278 -2404 18312
rect -2370 18278 -2336 18312
rect -2302 18278 -2268 18312
rect -2234 18278 -2200 18312
rect -2166 18278 -2132 18312
rect -2098 18278 -2064 18312
rect -2030 18278 -1996 18312
rect -1962 18278 -1928 18312
rect -1894 18278 -1860 18312
rect -1826 18278 -1792 18312
rect -1758 18278 -1724 18312
rect -1690 18278 -1656 18312
rect -1622 18278 -1588 18312
rect -1554 18278 -1520 18312
rect -1486 18278 -1452 18312
rect -1418 18278 -1384 18312
rect -1350 18278 -1316 18312
rect -1282 18278 -1248 18312
rect -1214 18278 -1180 18312
rect -1146 18278 -1112 18312
rect -1078 18278 -1044 18312
rect -1010 18278 -976 18312
rect -942 18278 -908 18312
rect -874 18278 -840 18312
rect -806 18278 -772 18312
rect -738 18278 -704 18312
rect -670 18278 -636 18312
rect -602 18278 -568 18312
rect -534 18278 -500 18312
rect -466 18278 -432 18312
rect -398 18278 -364 18312
rect -330 18278 -220 18312
rect -3126 18266 -220 18278
rect -3126 18198 -3068 18266
rect -3126 18164 -3114 18198
rect -3080 18164 -3068 18198
rect -278 18198 -220 18266
rect -3126 18130 -3068 18164
rect -3126 18096 -3114 18130
rect -3080 18096 -3068 18130
rect -3126 18062 -3068 18096
rect -278 18164 -266 18198
rect -232 18164 -220 18198
rect -278 18130 -220 18164
rect -278 18096 -266 18130
rect -232 18096 -220 18130
rect -3126 18028 -3114 18062
rect -3080 18028 -3068 18062
rect -3126 17994 -3068 18028
rect -3126 17960 -3114 17994
rect -3080 17960 -3068 17994
rect -3126 17926 -3068 17960
rect -3126 17892 -3114 17926
rect -3080 17892 -3068 17926
rect -3126 17858 -3068 17892
rect -3126 17824 -3114 17858
rect -3080 17824 -3068 17858
rect -3126 17790 -3068 17824
rect -3126 17756 -3114 17790
rect -3080 17756 -3068 17790
rect -3126 17722 -3068 17756
rect -3126 17688 -3114 17722
rect -3080 17688 -3068 17722
rect -3126 17654 -3068 17688
rect -3126 17620 -3114 17654
rect -3080 17620 -3068 17654
rect -3126 17586 -3068 17620
rect -6816 17536 -5446 17564
rect -6816 17502 -6702 17536
rect -6668 17502 -6634 17536
rect -6600 17502 -6566 17536
rect -6532 17502 -6498 17536
rect -6464 17502 -6430 17536
rect -6396 17502 -6362 17536
rect -6328 17502 -6294 17536
rect -6260 17502 -6226 17536
rect -6192 17502 -6158 17536
rect -6124 17502 -6090 17536
rect -6056 17502 -6022 17536
rect -5988 17502 -5954 17536
rect -5920 17502 -5886 17536
rect -5852 17502 -5818 17536
rect -5784 17502 -5750 17536
rect -5716 17502 -5682 17536
rect -5648 17502 -5614 17536
rect -5580 17502 -5446 17536
rect -6816 17484 -5446 17502
rect -6816 17441 -6736 17484
rect -6816 17407 -6798 17441
rect -6764 17407 -6736 17441
rect -6816 17373 -6736 17407
rect -6816 17339 -6798 17373
rect -6764 17339 -6736 17373
rect -6816 17305 -6736 17339
rect -5526 17461 -5446 17484
rect -5526 17427 -5508 17461
rect -5474 17427 -5446 17461
rect -5526 17393 -5446 17427
rect -5526 17359 -5508 17393
rect -5474 17359 -5446 17393
rect -5526 17325 -5446 17359
rect -6816 17271 -6798 17305
rect -6764 17271 -6736 17305
rect -6816 17237 -6736 17271
rect -6816 17203 -6798 17237
rect -6764 17203 -6736 17237
rect -5526 17291 -5508 17325
rect -5474 17291 -5446 17325
rect -5526 17257 -5446 17291
rect -6816 17169 -6736 17203
rect -6816 17135 -6798 17169
rect -6764 17135 -6736 17169
rect -6816 17101 -6736 17135
rect -6816 17067 -6798 17101
rect -6764 17067 -6736 17101
rect -6816 17033 -6736 17067
rect -6816 16999 -6798 17033
rect -6764 16999 -6736 17033
rect -6816 16965 -6736 16999
rect -6816 16931 -6798 16965
rect -6764 16931 -6736 16965
rect -6816 16897 -6736 16931
rect -6816 16863 -6798 16897
rect -6764 16863 -6736 16897
rect -6816 16829 -6736 16863
rect -6816 16795 -6798 16829
rect -6764 16795 -6736 16829
rect -6816 16761 -6736 16795
rect -6816 16727 -6798 16761
rect -6764 16727 -6736 16761
rect -6816 16693 -6736 16727
rect -6816 16659 -6798 16693
rect -6764 16659 -6736 16693
rect -6816 16625 -6736 16659
rect -6816 16591 -6798 16625
rect -6764 16591 -6736 16625
rect -6816 16557 -6736 16591
rect -6816 16523 -6798 16557
rect -6764 16523 -6736 16557
rect -6816 16489 -6736 16523
rect -6816 16455 -6798 16489
rect -6764 16455 -6736 16489
rect -6816 16421 -6736 16455
rect -6816 16387 -6798 16421
rect -6764 16387 -6736 16421
rect -6816 16353 -6736 16387
rect -6816 16319 -6798 16353
rect -6764 16319 -6736 16353
rect -6816 16285 -6736 16319
rect -6816 16251 -6798 16285
rect -6764 16251 -6736 16285
rect -6816 16217 -6736 16251
rect -5526 17223 -5508 17257
rect -5474 17223 -5446 17257
rect -5526 17189 -5446 17223
rect -5526 17155 -5508 17189
rect -5474 17155 -5446 17189
rect -5526 17121 -5446 17155
rect -5526 17087 -5508 17121
rect -5474 17087 -5446 17121
rect -5526 17053 -5446 17087
rect -5526 17019 -5508 17053
rect -5474 17019 -5446 17053
rect -5526 16985 -5446 17019
rect -5526 16951 -5508 16985
rect -5474 16951 -5446 16985
rect -5526 16917 -5446 16951
rect -5526 16883 -5508 16917
rect -5474 16883 -5446 16917
rect -5526 16849 -5446 16883
rect -5526 16815 -5508 16849
rect -5474 16815 -5446 16849
rect -5526 16781 -5446 16815
rect -5526 16747 -5508 16781
rect -5474 16747 -5446 16781
rect -5526 16713 -5446 16747
rect -5526 16679 -5508 16713
rect -5474 16679 -5446 16713
rect -5526 16645 -5446 16679
rect -5526 16611 -5508 16645
rect -5474 16611 -5446 16645
rect -5526 16577 -5446 16611
rect -5526 16543 -5508 16577
rect -5474 16543 -5446 16577
rect -5526 16509 -5446 16543
rect -5526 16475 -5508 16509
rect -5474 16475 -5446 16509
rect -5526 16441 -5446 16475
rect -5526 16407 -5508 16441
rect -5474 16407 -5446 16441
rect -5526 16373 -5446 16407
rect -5526 16339 -5508 16373
rect -5474 16339 -5446 16373
rect -5526 16305 -5446 16339
rect -5526 16271 -5508 16305
rect -5474 16271 -5446 16305
rect -5526 16237 -5446 16271
rect -6816 16183 -6798 16217
rect -6764 16183 -6736 16217
rect -6816 16149 -6736 16183
rect -6816 16115 -6798 16149
rect -6764 16115 -6736 16149
rect -5526 16203 -5508 16237
rect -5474 16203 -5446 16237
rect -5526 16169 -5446 16203
rect -5526 16135 -5508 16169
rect -5474 16135 -5446 16169
rect -6816 16081 -6736 16115
rect -6816 16047 -6798 16081
rect -6764 16047 -6736 16081
rect -6816 16024 -6736 16047
rect -5526 16101 -5446 16135
rect -5526 16067 -5508 16101
rect -5474 16067 -5446 16101
rect -5526 16024 -5446 16067
rect -6816 15996 -5446 16024
rect -6816 15962 -6682 15996
rect -6648 15962 -6614 15996
rect -6580 15962 -6546 15996
rect -6512 15962 -6478 15996
rect -6444 15962 -6410 15996
rect -6376 15962 -6342 15996
rect -6308 15962 -6274 15996
rect -6240 15962 -6206 15996
rect -6172 15962 -6138 15996
rect -6104 15962 -6070 15996
rect -6036 15962 -6002 15996
rect -5968 15962 -5934 15996
rect -5900 15962 -5866 15996
rect -5832 15962 -5798 15996
rect -5764 15962 -5730 15996
rect -5696 15962 -5662 15996
rect -5628 15962 -5594 15996
rect -5560 15962 -5446 15996
rect -6816 15944 -5446 15962
rect -3126 17552 -3114 17586
rect -3080 17552 -3068 17586
rect -3126 17518 -3068 17552
rect -3126 17484 -3114 17518
rect -3080 17484 -3068 17518
rect -3126 17450 -3068 17484
rect -3126 17416 -3114 17450
rect -3080 17416 -3068 17450
rect -3126 17382 -3068 17416
rect -3126 17348 -3114 17382
rect -3080 17348 -3068 17382
rect -3126 17314 -3068 17348
rect -3126 17280 -3114 17314
rect -3080 17280 -3068 17314
rect -3126 17246 -3068 17280
rect -3126 17212 -3114 17246
rect -3080 17212 -3068 17246
rect -3126 17178 -3068 17212
rect -3126 17144 -3114 17178
rect -3080 17144 -3068 17178
rect -3126 17110 -3068 17144
rect -3126 17076 -3114 17110
rect -3080 17076 -3068 17110
rect -3126 17042 -3068 17076
rect -3126 17008 -3114 17042
rect -3080 17008 -3068 17042
rect -3126 16974 -3068 17008
rect -3126 16940 -3114 16974
rect -3080 16940 -3068 16974
rect -3126 16906 -3068 16940
rect -3126 16872 -3114 16906
rect -3080 16872 -3068 16906
rect -3126 16838 -3068 16872
rect -3126 16804 -3114 16838
rect -3080 16804 -3068 16838
rect -3126 16770 -3068 16804
rect -3126 16736 -3114 16770
rect -3080 16736 -3068 16770
rect -3126 16702 -3068 16736
rect -3126 16668 -3114 16702
rect -3080 16668 -3068 16702
rect -3126 16634 -3068 16668
rect -3126 16600 -3114 16634
rect -3080 16600 -3068 16634
rect -3126 16566 -3068 16600
rect -3126 16532 -3114 16566
rect -3080 16532 -3068 16566
rect -3126 16498 -3068 16532
rect -3126 16464 -3114 16498
rect -3080 16464 -3068 16498
rect -3126 16430 -3068 16464
rect -3126 16396 -3114 16430
rect -3080 16396 -3068 16430
rect -3126 16362 -3068 16396
rect -3126 16328 -3114 16362
rect -3080 16328 -3068 16362
rect -3126 16294 -3068 16328
rect -3126 16260 -3114 16294
rect -3080 16260 -3068 16294
rect -3126 16226 -3068 16260
rect -3126 16192 -3114 16226
rect -3080 16192 -3068 16226
rect -3126 16158 -3068 16192
rect -3126 16124 -3114 16158
rect -3080 16124 -3068 16158
rect -3126 16090 -3068 16124
rect -278 18062 -220 18096
rect -278 18028 -266 18062
rect -232 18028 -220 18062
rect -278 17994 -220 18028
rect -278 17960 -266 17994
rect -232 17960 -220 17994
rect -278 17926 -220 17960
rect -278 17892 -266 17926
rect -232 17892 -220 17926
rect -278 17858 -220 17892
rect -278 17824 -266 17858
rect -232 17824 -220 17858
rect -278 17790 -220 17824
rect -278 17756 -266 17790
rect -232 17756 -220 17790
rect -278 17722 -220 17756
rect -278 17688 -266 17722
rect -232 17688 -220 17722
rect -278 17654 -220 17688
rect -278 17620 -266 17654
rect -232 17620 -220 17654
rect -278 17586 -220 17620
rect -278 17552 -266 17586
rect -232 17552 -220 17586
rect -278 17518 -220 17552
rect -278 17484 -266 17518
rect -232 17484 -220 17518
rect 23030 18298 23088 18332
rect 23030 18264 23042 18298
rect 23076 18264 23088 18298
rect 23030 18230 23088 18264
rect 23030 18196 23042 18230
rect 23076 18196 23088 18230
rect 23030 18162 23088 18196
rect 23030 18128 23042 18162
rect 23076 18128 23088 18162
rect 23030 18094 23088 18128
rect 23030 18060 23042 18094
rect 23076 18060 23088 18094
rect 23030 18026 23088 18060
rect 23030 17992 23042 18026
rect 23076 17992 23088 18026
rect 23030 17958 23088 17992
rect 23030 17924 23042 17958
rect 23076 17924 23088 17958
rect 23030 17890 23088 17924
rect 23030 17856 23042 17890
rect 23076 17856 23088 17890
rect 23030 17822 23088 17856
rect 23030 17788 23042 17822
rect 23076 17788 23088 17822
rect 23030 17754 23088 17788
rect 23030 17720 23042 17754
rect 23076 17720 23088 17754
rect 24356 18740 24368 18774
rect 24402 18740 24414 18774
rect 24356 18706 24414 18740
rect 24356 18672 24368 18706
rect 24402 18672 24414 18706
rect 24356 18638 24414 18672
rect 24356 18604 24368 18638
rect 24402 18604 24414 18638
rect 24356 18570 24414 18604
rect 24356 18536 24368 18570
rect 24402 18536 24414 18570
rect 24356 18502 24414 18536
rect 24356 18468 24368 18502
rect 24402 18468 24414 18502
rect 24356 18434 24414 18468
rect 24356 18400 24368 18434
rect 24402 18400 24414 18434
rect 24356 18366 24414 18400
rect 24356 18332 24368 18366
rect 24402 18332 24414 18366
rect 24356 18298 24414 18332
rect 24356 18264 24368 18298
rect 24402 18264 24414 18298
rect 24356 18230 24414 18264
rect 24356 18196 24368 18230
rect 24402 18196 24414 18230
rect 24356 18162 24414 18196
rect 24356 18128 24368 18162
rect 24402 18128 24414 18162
rect 24356 18094 24414 18128
rect 24356 18060 24368 18094
rect 24402 18060 24414 18094
rect 24356 18026 24414 18060
rect 24356 17992 24368 18026
rect 24402 17992 24414 18026
rect 24356 17958 24414 17992
rect 24356 17924 24368 17958
rect 24402 17924 24414 17958
rect 24356 17890 24414 17924
rect 24356 17856 24368 17890
rect 24402 17856 24414 17890
rect 24356 17822 24414 17856
rect 24356 17788 24368 17822
rect 24402 17788 24414 17822
rect 24356 17754 24414 17788
rect 23030 17686 23088 17720
rect 23030 17652 23042 17686
rect 23076 17652 23088 17686
rect 23030 17574 23088 17652
rect 24356 17720 24368 17754
rect 24402 17720 24414 17754
rect 24356 17686 24414 17720
rect 24356 17652 24368 17686
rect 24402 17652 24414 17686
rect 24356 17574 24414 17652
rect 23030 17562 24414 17574
rect 23030 17528 23161 17562
rect 23195 17528 23229 17562
rect 23263 17528 23297 17562
rect 23331 17528 23365 17562
rect 23399 17528 23433 17562
rect 23467 17528 23501 17562
rect 23535 17528 23569 17562
rect 23603 17528 23637 17562
rect 23671 17528 23705 17562
rect 23739 17528 23773 17562
rect 23807 17528 23841 17562
rect 23875 17528 23909 17562
rect 23943 17528 23977 17562
rect 24011 17528 24045 17562
rect 24079 17528 24113 17562
rect 24147 17528 24181 17562
rect 24215 17528 24249 17562
rect 24283 17528 24414 17562
rect 23030 17516 24414 17528
rect 24546 18966 28046 18978
rect 24546 18932 24681 18966
rect 24715 18932 24749 18966
rect 24783 18932 24817 18966
rect 24851 18932 24885 18966
rect 24919 18932 24953 18966
rect 24987 18932 25021 18966
rect 25055 18932 25089 18966
rect 25123 18932 25157 18966
rect 25191 18932 25225 18966
rect 25259 18932 25293 18966
rect 25327 18932 25361 18966
rect 25395 18932 25429 18966
rect 25463 18932 25497 18966
rect 25531 18932 25565 18966
rect 25599 18932 25633 18966
rect 25667 18932 25701 18966
rect 25735 18932 25769 18966
rect 25803 18932 25837 18966
rect 25871 18932 25905 18966
rect 25939 18932 25973 18966
rect 26007 18932 26041 18966
rect 26075 18932 26109 18966
rect 26143 18932 26177 18966
rect 26211 18932 26245 18966
rect 26279 18932 26313 18966
rect 26347 18932 26381 18966
rect 26415 18932 26449 18966
rect 26483 18932 26517 18966
rect 26551 18932 26585 18966
rect 26619 18932 26653 18966
rect 26687 18932 26721 18966
rect 26755 18932 26789 18966
rect 26823 18932 26857 18966
rect 26891 18932 26925 18966
rect 26959 18932 26993 18966
rect 27027 18932 27061 18966
rect 27095 18932 27129 18966
rect 27163 18932 27197 18966
rect 27231 18932 27265 18966
rect 27299 18932 27333 18966
rect 27367 18932 27401 18966
rect 27435 18932 27469 18966
rect 27503 18932 27537 18966
rect 27571 18932 27605 18966
rect 27639 18932 27673 18966
rect 27707 18932 27741 18966
rect 27775 18932 27809 18966
rect 27843 18932 27877 18966
rect 27911 18932 28046 18966
rect 24546 18920 28046 18932
rect 24546 18848 24604 18920
rect 24546 18814 24558 18848
rect 24592 18814 24604 18848
rect 27988 18848 28046 18920
rect 24546 18780 24604 18814
rect 24546 18746 24558 18780
rect 24592 18746 24604 18780
rect 27988 18814 28000 18848
rect 28034 18814 28046 18848
rect 27988 18780 28046 18814
rect 24546 18712 24604 18746
rect 24546 18678 24558 18712
rect 24592 18678 24604 18712
rect 24546 18644 24604 18678
rect 24546 18610 24558 18644
rect 24592 18610 24604 18644
rect 24546 18576 24604 18610
rect 24546 18542 24558 18576
rect 24592 18542 24604 18576
rect 24546 18508 24604 18542
rect 24546 18474 24558 18508
rect 24592 18474 24604 18508
rect 24546 18440 24604 18474
rect 24546 18406 24558 18440
rect 24592 18406 24604 18440
rect 24546 18372 24604 18406
rect 24546 18338 24558 18372
rect 24592 18338 24604 18372
rect 24546 18304 24604 18338
rect 24546 18270 24558 18304
rect 24592 18270 24604 18304
rect 24546 18236 24604 18270
rect 24546 18202 24558 18236
rect 24592 18202 24604 18236
rect 24546 18168 24604 18202
rect 24546 18134 24558 18168
rect 24592 18134 24604 18168
rect 24546 18100 24604 18134
rect 24546 18066 24558 18100
rect 24592 18066 24604 18100
rect 24546 18032 24604 18066
rect 24546 17998 24558 18032
rect 24592 17998 24604 18032
rect 24546 17964 24604 17998
rect 24546 17930 24558 17964
rect 24592 17930 24604 17964
rect 24546 17896 24604 17930
rect 24546 17862 24558 17896
rect 24592 17862 24604 17896
rect 24546 17828 24604 17862
rect 24546 17794 24558 17828
rect 24592 17794 24604 17828
rect 24546 17760 24604 17794
rect 24546 17726 24558 17760
rect 24592 17726 24604 17760
rect 24546 17692 24604 17726
rect 24546 17658 24558 17692
rect 24592 17658 24604 17692
rect 24546 17624 24604 17658
rect 24546 17590 24558 17624
rect 24592 17590 24604 17624
rect 24546 17556 24604 17590
rect 24546 17522 24558 17556
rect 24592 17522 24604 17556
rect -278 17450 -220 17484
rect -278 17416 -266 17450
rect -232 17416 -220 17450
rect -278 17382 -220 17416
rect -278 17348 -266 17382
rect -232 17348 -220 17382
rect 24546 17488 24604 17522
rect 24546 17454 24558 17488
rect 24592 17454 24604 17488
rect 24546 17420 24604 17454
rect 24546 17386 24558 17420
rect 24592 17386 24604 17420
rect -278 17314 -220 17348
rect -278 17280 -266 17314
rect -232 17280 -220 17314
rect -278 17246 -220 17280
rect -278 17212 -266 17246
rect -232 17212 -220 17246
rect -278 17178 -220 17212
rect -278 17144 -266 17178
rect -232 17144 -220 17178
rect -278 17110 -220 17144
rect -278 17076 -266 17110
rect -232 17076 -220 17110
rect -278 17042 -220 17076
rect -278 17008 -266 17042
rect -232 17008 -220 17042
rect -278 16974 -220 17008
rect -278 16940 -266 16974
rect -232 16940 -220 16974
rect -278 16906 -220 16940
rect -278 16872 -266 16906
rect -232 16872 -220 16906
rect -278 16838 -220 16872
rect -278 16804 -266 16838
rect -232 16804 -220 16838
rect -278 16770 -220 16804
rect -278 16736 -266 16770
rect -232 16736 -220 16770
rect -278 16702 -220 16736
rect -278 16668 -266 16702
rect -232 16668 -220 16702
rect -278 16634 -220 16668
rect -278 16600 -266 16634
rect -232 16600 -220 16634
rect -278 16566 -220 16600
rect -278 16532 -266 16566
rect -232 16532 -220 16566
rect -278 16498 -220 16532
rect -278 16464 -266 16498
rect -232 16464 -220 16498
rect -278 16430 -220 16464
rect -278 16396 -266 16430
rect -232 16396 -220 16430
rect -278 16362 -220 16396
rect -278 16328 -266 16362
rect -232 16328 -220 16362
rect -278 16294 -220 16328
rect -278 16260 -266 16294
rect -232 16260 -220 16294
rect -278 16226 -220 16260
rect -278 16192 -266 16226
rect -232 16192 -220 16226
rect -278 16158 -220 16192
rect -278 16124 -266 16158
rect -232 16124 -220 16158
rect -3126 16056 -3114 16090
rect -3080 16056 -3068 16090
rect -3126 16022 -3068 16056
rect -3126 15988 -3114 16022
rect -3080 15988 -3068 16022
rect -278 16090 -220 16124
rect -278 16056 -266 16090
rect -232 16056 -220 16090
rect -278 16022 -220 16056
rect -3126 15920 -3068 15988
rect -278 15988 -266 16022
rect -232 15988 -220 16022
rect -278 15920 -220 15988
rect -3126 15908 -220 15920
rect 24546 17352 24604 17386
rect 24546 17318 24558 17352
rect 24592 17318 24604 17352
rect 24546 17284 24604 17318
rect 24546 17250 24558 17284
rect 24592 17250 24604 17284
rect 24546 17216 24604 17250
rect 24546 17182 24558 17216
rect 24592 17182 24604 17216
rect 24546 17148 24604 17182
rect 24546 17114 24558 17148
rect 24592 17114 24604 17148
rect 27988 18746 28000 18780
rect 28034 18746 28046 18780
rect 27988 18712 28046 18746
rect 27988 18678 28000 18712
rect 28034 18678 28046 18712
rect 27988 18644 28046 18678
rect 27988 18610 28000 18644
rect 28034 18610 28046 18644
rect 27988 18576 28046 18610
rect 27988 18542 28000 18576
rect 28034 18542 28046 18576
rect 27988 18508 28046 18542
rect 27988 18474 28000 18508
rect 28034 18474 28046 18508
rect 27988 18440 28046 18474
rect 27988 18406 28000 18440
rect 28034 18406 28046 18440
rect 27988 18372 28046 18406
rect 27988 18338 28000 18372
rect 28034 18338 28046 18372
rect 27988 18304 28046 18338
rect 42466 18948 42524 19016
rect 42466 18914 42478 18948
rect 42512 18914 42524 18948
rect 45314 18948 45372 19016
rect 42466 18880 42524 18914
rect 42466 18846 42478 18880
rect 42512 18846 42524 18880
rect 42466 18812 42524 18846
rect 45314 18914 45326 18948
rect 45360 18914 45372 18948
rect 45314 18880 45372 18914
rect 45314 18846 45326 18880
rect 45360 18846 45372 18880
rect 42466 18778 42478 18812
rect 42512 18778 42524 18812
rect 42466 18744 42524 18778
rect 42466 18710 42478 18744
rect 42512 18710 42524 18744
rect 42466 18676 42524 18710
rect 42466 18642 42478 18676
rect 42512 18642 42524 18676
rect 42466 18608 42524 18642
rect 42466 18574 42478 18608
rect 42512 18574 42524 18608
rect 42466 18540 42524 18574
rect 42466 18506 42478 18540
rect 42512 18506 42524 18540
rect 42466 18472 42524 18506
rect 42466 18438 42478 18472
rect 42512 18438 42524 18472
rect 42466 18404 42524 18438
rect 42466 18370 42478 18404
rect 42512 18370 42524 18404
rect 42466 18336 42524 18370
rect 27988 18270 28000 18304
rect 28034 18270 28046 18304
rect 27988 18236 28046 18270
rect 27988 18202 28000 18236
rect 28034 18202 28046 18236
rect 27988 18168 28046 18202
rect 27988 18134 28000 18168
rect 28034 18134 28046 18168
rect 27988 18100 28046 18134
rect 27988 18066 28000 18100
rect 28034 18066 28046 18100
rect 27988 18032 28046 18066
rect 27988 17998 28000 18032
rect 28034 17998 28046 18032
rect 27988 17964 28046 17998
rect 27988 17930 28000 17964
rect 28034 17930 28046 17964
rect 27988 17896 28046 17930
rect 27988 17862 28000 17896
rect 28034 17862 28046 17896
rect 27988 17828 28046 17862
rect 27988 17794 28000 17828
rect 28034 17794 28046 17828
rect 27988 17760 28046 17794
rect 27988 17726 28000 17760
rect 28034 17726 28046 17760
rect 27988 17692 28046 17726
rect 27988 17658 28000 17692
rect 28034 17658 28046 17692
rect 27988 17624 28046 17658
rect 27988 17590 28000 17624
rect 28034 17590 28046 17624
rect 27988 17556 28046 17590
rect 27988 17522 28000 17556
rect 28034 17522 28046 17556
rect 27988 17488 28046 17522
rect 27988 17454 28000 17488
rect 28034 17454 28046 17488
rect 27988 17420 28046 17454
rect 27988 17386 28000 17420
rect 28034 17386 28046 17420
rect 27988 17352 28046 17386
rect 27988 17318 28000 17352
rect 28034 17318 28046 17352
rect 27988 17284 28046 17318
rect 27988 17250 28000 17284
rect 28034 17250 28046 17284
rect 27988 17216 28046 17250
rect 27988 17182 28000 17216
rect 28034 17182 28046 17216
rect 27988 17148 28046 17182
rect 24546 17080 24604 17114
rect 24546 17046 24558 17080
rect 24592 17046 24604 17080
rect 27988 17114 28000 17148
rect 28034 17114 28046 17148
rect 27988 17080 28046 17114
rect 24546 16974 24604 17046
rect 27988 17046 28000 17080
rect 28034 17046 28046 17080
rect 27988 16974 28046 17046
rect 24546 16962 28046 16974
rect 24546 16928 24681 16962
rect 24715 16928 24749 16962
rect 24783 16928 24817 16962
rect 24851 16928 24885 16962
rect 24919 16928 24953 16962
rect 24987 16928 25021 16962
rect 25055 16928 25089 16962
rect 25123 16928 25157 16962
rect 25191 16928 25225 16962
rect 25259 16928 25293 16962
rect 25327 16928 25361 16962
rect 25395 16928 25429 16962
rect 25463 16928 25497 16962
rect 25531 16928 25565 16962
rect 25599 16928 25633 16962
rect 25667 16928 25701 16962
rect 25735 16928 25769 16962
rect 25803 16928 25837 16962
rect 25871 16928 25905 16962
rect 25939 16928 25973 16962
rect 26007 16928 26041 16962
rect 26075 16928 26109 16962
rect 26143 16928 26177 16962
rect 26211 16928 26245 16962
rect 26279 16928 26313 16962
rect 26347 16928 26381 16962
rect 26415 16928 26449 16962
rect 26483 16928 26517 16962
rect 26551 16928 26585 16962
rect 26619 16928 26653 16962
rect 26687 16928 26721 16962
rect 26755 16928 26789 16962
rect 26823 16928 26857 16962
rect 26891 16928 26925 16962
rect 26959 16928 26993 16962
rect 27027 16928 27061 16962
rect 27095 16928 27129 16962
rect 27163 16928 27197 16962
rect 27231 16928 27265 16962
rect 27299 16928 27333 16962
rect 27367 16928 27401 16962
rect 27435 16928 27469 16962
rect 27503 16928 27537 16962
rect 27571 16928 27605 16962
rect 27639 16928 27673 16962
rect 27707 16928 27741 16962
rect 27775 16928 27809 16962
rect 27843 16928 27877 16962
rect 27911 16928 28046 16962
rect 24546 16916 28046 16928
rect 38776 18286 40146 18314
rect 38776 18252 38890 18286
rect 38924 18252 38958 18286
rect 38992 18252 39026 18286
rect 39060 18252 39094 18286
rect 39128 18252 39162 18286
rect 39196 18252 39230 18286
rect 39264 18252 39298 18286
rect 39332 18252 39366 18286
rect 39400 18252 39434 18286
rect 39468 18252 39502 18286
rect 39536 18252 39570 18286
rect 39604 18252 39638 18286
rect 39672 18252 39706 18286
rect 39740 18252 39774 18286
rect 39808 18252 39842 18286
rect 39876 18252 39910 18286
rect 39944 18252 39978 18286
rect 40012 18252 40146 18286
rect 38776 18234 40146 18252
rect 38776 18191 38856 18234
rect 38776 18157 38794 18191
rect 38828 18157 38856 18191
rect 38776 18123 38856 18157
rect 38776 18089 38794 18123
rect 38828 18089 38856 18123
rect 38776 18055 38856 18089
rect 40066 18211 40146 18234
rect 40066 18177 40084 18211
rect 40118 18177 40146 18211
rect 40066 18143 40146 18177
rect 40066 18109 40084 18143
rect 40118 18109 40146 18143
rect 40066 18075 40146 18109
rect 38776 18021 38794 18055
rect 38828 18021 38856 18055
rect 38776 17987 38856 18021
rect 38776 17953 38794 17987
rect 38828 17953 38856 17987
rect 40066 18041 40084 18075
rect 40118 18041 40146 18075
rect 40066 18007 40146 18041
rect 38776 17919 38856 17953
rect 38776 17885 38794 17919
rect 38828 17885 38856 17919
rect 38776 17851 38856 17885
rect 38776 17817 38794 17851
rect 38828 17817 38856 17851
rect 38776 17783 38856 17817
rect 38776 17749 38794 17783
rect 38828 17749 38856 17783
rect 38776 17715 38856 17749
rect 38776 17681 38794 17715
rect 38828 17681 38856 17715
rect 38776 17647 38856 17681
rect 38776 17613 38794 17647
rect 38828 17613 38856 17647
rect 38776 17579 38856 17613
rect 38776 17545 38794 17579
rect 38828 17545 38856 17579
rect 38776 17511 38856 17545
rect 38776 17477 38794 17511
rect 38828 17477 38856 17511
rect 38776 17443 38856 17477
rect 38776 17409 38794 17443
rect 38828 17409 38856 17443
rect 38776 17375 38856 17409
rect 38776 17341 38794 17375
rect 38828 17341 38856 17375
rect 38776 17307 38856 17341
rect 38776 17273 38794 17307
rect 38828 17273 38856 17307
rect 38776 17239 38856 17273
rect 38776 17205 38794 17239
rect 38828 17205 38856 17239
rect 38776 17171 38856 17205
rect 38776 17137 38794 17171
rect 38828 17137 38856 17171
rect 38776 17103 38856 17137
rect 38776 17069 38794 17103
rect 38828 17069 38856 17103
rect 38776 17035 38856 17069
rect 38776 17001 38794 17035
rect 38828 17001 38856 17035
rect 38776 16967 38856 17001
rect 40066 17973 40084 18007
rect 40118 17973 40146 18007
rect 40066 17939 40146 17973
rect 40066 17905 40084 17939
rect 40118 17905 40146 17939
rect 40066 17871 40146 17905
rect 40066 17837 40084 17871
rect 40118 17837 40146 17871
rect 40066 17803 40146 17837
rect 40066 17769 40084 17803
rect 40118 17769 40146 17803
rect 40066 17735 40146 17769
rect 40066 17701 40084 17735
rect 40118 17701 40146 17735
rect 40066 17667 40146 17701
rect 40066 17633 40084 17667
rect 40118 17633 40146 17667
rect 40066 17599 40146 17633
rect 40066 17565 40084 17599
rect 40118 17565 40146 17599
rect 40066 17531 40146 17565
rect 40066 17497 40084 17531
rect 40118 17497 40146 17531
rect 40066 17463 40146 17497
rect 40066 17429 40084 17463
rect 40118 17429 40146 17463
rect 40066 17395 40146 17429
rect 40066 17361 40084 17395
rect 40118 17361 40146 17395
rect 40066 17327 40146 17361
rect 40066 17293 40084 17327
rect 40118 17293 40146 17327
rect 40066 17259 40146 17293
rect 40066 17225 40084 17259
rect 40118 17225 40146 17259
rect 40066 17191 40146 17225
rect 40066 17157 40084 17191
rect 40118 17157 40146 17191
rect 40066 17123 40146 17157
rect 40066 17089 40084 17123
rect 40118 17089 40146 17123
rect 40066 17055 40146 17089
rect 40066 17021 40084 17055
rect 40118 17021 40146 17055
rect 40066 16987 40146 17021
rect 38776 16933 38794 16967
rect 38828 16933 38856 16967
rect 38776 16899 38856 16933
rect 38776 16865 38794 16899
rect 38828 16865 38856 16899
rect 40066 16953 40084 16987
rect 40118 16953 40146 16987
rect 40066 16919 40146 16953
rect 40066 16885 40084 16919
rect 40118 16885 40146 16919
rect 38776 16831 38856 16865
rect 38776 16797 38794 16831
rect 38828 16797 38856 16831
rect 38776 16774 38856 16797
rect 40066 16851 40146 16885
rect 40066 16817 40084 16851
rect 40118 16817 40146 16851
rect 40066 16774 40146 16817
rect 38776 16746 40146 16774
rect 38776 16712 38910 16746
rect 38944 16712 38978 16746
rect 39012 16712 39046 16746
rect 39080 16712 39114 16746
rect 39148 16712 39182 16746
rect 39216 16712 39250 16746
rect 39284 16712 39318 16746
rect 39352 16712 39386 16746
rect 39420 16712 39454 16746
rect 39488 16712 39522 16746
rect 39556 16712 39590 16746
rect 39624 16712 39658 16746
rect 39692 16712 39726 16746
rect 39760 16712 39794 16746
rect 39828 16712 39862 16746
rect 39896 16712 39930 16746
rect 39964 16712 39998 16746
rect 40032 16712 40146 16746
rect 38776 16694 40146 16712
rect 42466 18302 42478 18336
rect 42512 18302 42524 18336
rect 42466 18268 42524 18302
rect 42466 18234 42478 18268
rect 42512 18234 42524 18268
rect 42466 18200 42524 18234
rect 42466 18166 42478 18200
rect 42512 18166 42524 18200
rect 42466 18132 42524 18166
rect 42466 18098 42478 18132
rect 42512 18098 42524 18132
rect 42466 18064 42524 18098
rect 42466 18030 42478 18064
rect 42512 18030 42524 18064
rect 42466 17996 42524 18030
rect 42466 17962 42478 17996
rect 42512 17962 42524 17996
rect 42466 17928 42524 17962
rect 42466 17894 42478 17928
rect 42512 17894 42524 17928
rect 42466 17860 42524 17894
rect 42466 17826 42478 17860
rect 42512 17826 42524 17860
rect 42466 17792 42524 17826
rect 42466 17758 42478 17792
rect 42512 17758 42524 17792
rect 42466 17724 42524 17758
rect 42466 17690 42478 17724
rect 42512 17690 42524 17724
rect 42466 17656 42524 17690
rect 42466 17622 42478 17656
rect 42512 17622 42524 17656
rect 42466 17588 42524 17622
rect 42466 17554 42478 17588
rect 42512 17554 42524 17588
rect 42466 17520 42524 17554
rect 42466 17486 42478 17520
rect 42512 17486 42524 17520
rect 42466 17452 42524 17486
rect 42466 17418 42478 17452
rect 42512 17418 42524 17452
rect 42466 17384 42524 17418
rect 42466 17350 42478 17384
rect 42512 17350 42524 17384
rect 42466 17316 42524 17350
rect 42466 17282 42478 17316
rect 42512 17282 42524 17316
rect 42466 17248 42524 17282
rect 42466 17214 42478 17248
rect 42512 17214 42524 17248
rect 42466 17180 42524 17214
rect 42466 17146 42478 17180
rect 42512 17146 42524 17180
rect 42466 17112 42524 17146
rect 42466 17078 42478 17112
rect 42512 17078 42524 17112
rect 42466 17044 42524 17078
rect 42466 17010 42478 17044
rect 42512 17010 42524 17044
rect 42466 16976 42524 17010
rect 42466 16942 42478 16976
rect 42512 16942 42524 16976
rect 42466 16908 42524 16942
rect 42466 16874 42478 16908
rect 42512 16874 42524 16908
rect 42466 16840 42524 16874
rect 45314 18812 45372 18846
rect 45314 18778 45326 18812
rect 45360 18778 45372 18812
rect 45314 18744 45372 18778
rect 45314 18710 45326 18744
rect 45360 18710 45372 18744
rect 45314 18676 45372 18710
rect 45314 18642 45326 18676
rect 45360 18642 45372 18676
rect 45314 18608 45372 18642
rect 45314 18574 45326 18608
rect 45360 18574 45372 18608
rect 45314 18540 45372 18574
rect 45314 18506 45326 18540
rect 45360 18506 45372 18540
rect 45314 18472 45372 18506
rect 45314 18438 45326 18472
rect 45360 18438 45372 18472
rect 45314 18404 45372 18438
rect 45314 18370 45326 18404
rect 45360 18370 45372 18404
rect 45314 18336 45372 18370
rect 45314 18302 45326 18336
rect 45360 18302 45372 18336
rect 45314 18268 45372 18302
rect 45314 18234 45326 18268
rect 45360 18234 45372 18268
rect 45314 18200 45372 18234
rect 45314 18166 45326 18200
rect 45360 18166 45372 18200
rect 45314 18132 45372 18166
rect 45314 18098 45326 18132
rect 45360 18098 45372 18132
rect 45314 18064 45372 18098
rect 45314 18030 45326 18064
rect 45360 18030 45372 18064
rect 45314 17996 45372 18030
rect 45314 17962 45326 17996
rect 45360 17962 45372 17996
rect 45314 17928 45372 17962
rect 45314 17894 45326 17928
rect 45360 17894 45372 17928
rect 45314 17860 45372 17894
rect 45314 17826 45326 17860
rect 45360 17826 45372 17860
rect 45314 17792 45372 17826
rect 45314 17758 45326 17792
rect 45360 17758 45372 17792
rect 45314 17724 45372 17758
rect 45314 17690 45326 17724
rect 45360 17690 45372 17724
rect 45314 17656 45372 17690
rect 45314 17622 45326 17656
rect 45360 17622 45372 17656
rect 45314 17588 45372 17622
rect 45314 17554 45326 17588
rect 45360 17554 45372 17588
rect 45314 17520 45372 17554
rect 45314 17486 45326 17520
rect 45360 17486 45372 17520
rect 45314 17452 45372 17486
rect 45314 17418 45326 17452
rect 45360 17418 45372 17452
rect 45314 17384 45372 17418
rect 45314 17350 45326 17384
rect 45360 17350 45372 17384
rect 45314 17316 45372 17350
rect 45314 17282 45326 17316
rect 45360 17282 45372 17316
rect 45314 17248 45372 17282
rect 45314 17214 45326 17248
rect 45360 17214 45372 17248
rect 45314 17180 45372 17214
rect 45314 17146 45326 17180
rect 45360 17146 45372 17180
rect 45314 17112 45372 17146
rect 45314 17078 45326 17112
rect 45360 17078 45372 17112
rect 45314 17044 45372 17078
rect 45314 17010 45326 17044
rect 45360 17010 45372 17044
rect 45314 16976 45372 17010
rect 45314 16942 45326 16976
rect 45360 16942 45372 16976
rect 45314 16908 45372 16942
rect 45314 16874 45326 16908
rect 45360 16874 45372 16908
rect 42466 16806 42478 16840
rect 42512 16806 42524 16840
rect 42466 16772 42524 16806
rect 42466 16738 42478 16772
rect 42512 16738 42524 16772
rect 45314 16840 45372 16874
rect 45314 16806 45326 16840
rect 45360 16806 45372 16840
rect 45314 16772 45372 16806
rect 42466 16670 42524 16738
rect 45314 16738 45326 16772
rect 45360 16738 45372 16772
rect 45314 16670 45372 16738
rect 42466 16658 45372 16670
rect 42466 16624 42576 16658
rect 42610 16624 42644 16658
rect 42678 16624 42712 16658
rect 42746 16624 42780 16658
rect 42814 16624 42848 16658
rect 42882 16624 42916 16658
rect 42950 16624 42984 16658
rect 43018 16624 43052 16658
rect 43086 16624 43120 16658
rect 43154 16624 43188 16658
rect 43222 16624 43256 16658
rect 43290 16624 43324 16658
rect 43358 16624 43392 16658
rect 43426 16624 43460 16658
rect 43494 16624 43528 16658
rect 43562 16624 43596 16658
rect 43630 16624 43664 16658
rect 43698 16624 43732 16658
rect 43766 16624 43800 16658
rect 43834 16624 43868 16658
rect 43902 16624 43936 16658
rect 43970 16624 44004 16658
rect 44038 16624 44072 16658
rect 44106 16624 44140 16658
rect 44174 16624 44208 16658
rect 44242 16624 44276 16658
rect 44310 16624 44344 16658
rect 44378 16624 44412 16658
rect 44446 16624 44480 16658
rect 44514 16624 44548 16658
rect 44582 16624 44616 16658
rect 44650 16624 44684 16658
rect 44718 16624 44752 16658
rect 44786 16624 44820 16658
rect 44854 16624 44888 16658
rect 44922 16624 44956 16658
rect 44990 16624 45024 16658
rect 45058 16624 45092 16658
rect 45126 16624 45160 16658
rect 45194 16624 45228 16658
rect 45262 16624 45372 16658
rect 42466 16612 45372 16624
rect -3126 15874 -3016 15908
rect -2982 15874 -2948 15908
rect -2914 15874 -2880 15908
rect -2846 15874 -2812 15908
rect -2778 15874 -2744 15908
rect -2710 15874 -2676 15908
rect -2642 15874 -2608 15908
rect -2574 15874 -2540 15908
rect -2506 15874 -2472 15908
rect -2438 15874 -2404 15908
rect -2370 15874 -2336 15908
rect -2302 15874 -2268 15908
rect -2234 15874 -2200 15908
rect -2166 15874 -2132 15908
rect -2098 15874 -2064 15908
rect -2030 15874 -1996 15908
rect -1962 15874 -1928 15908
rect -1894 15874 -1860 15908
rect -1826 15874 -1792 15908
rect -1758 15874 -1724 15908
rect -1690 15874 -1656 15908
rect -1622 15874 -1588 15908
rect -1554 15874 -1520 15908
rect -1486 15874 -1452 15908
rect -1418 15874 -1384 15908
rect -1350 15874 -1316 15908
rect -1282 15874 -1248 15908
rect -1214 15874 -1180 15908
rect -1146 15874 -1112 15908
rect -1078 15874 -1044 15908
rect -1010 15874 -976 15908
rect -942 15874 -908 15908
rect -874 15874 -840 15908
rect -806 15874 -772 15908
rect -738 15874 -704 15908
rect -670 15874 -636 15908
rect -602 15874 -568 15908
rect -534 15874 -500 15908
rect -466 15874 -432 15908
rect -398 15874 -364 15908
rect -330 15874 -220 15908
rect -3126 15862 -220 15874
rect 12848 14986 15290 14998
rect 12848 14952 12964 14986
rect 12998 14952 13032 14986
rect 13066 14952 13100 14986
rect 13134 14952 13168 14986
rect 13202 14952 13236 14986
rect 13270 14952 13304 14986
rect 13338 14952 13372 14986
rect 13406 14952 13440 14986
rect 13474 14952 13508 14986
rect 13542 14952 13576 14986
rect 13610 14952 13644 14986
rect 13678 14952 13712 14986
rect 13746 14952 13780 14986
rect 13814 14952 13848 14986
rect 13882 14952 13916 14986
rect 13950 14952 13984 14986
rect 14018 14952 14052 14986
rect 14086 14952 14120 14986
rect 14154 14952 14188 14986
rect 14222 14952 14256 14986
rect 14290 14952 14324 14986
rect 14358 14952 14392 14986
rect 14426 14952 14460 14986
rect 14494 14952 14528 14986
rect 14562 14952 14596 14986
rect 14630 14952 14664 14986
rect 14698 14952 14732 14986
rect 14766 14952 14800 14986
rect 14834 14952 14868 14986
rect 14902 14952 14936 14986
rect 14970 14952 15004 14986
rect 15038 14952 15072 14986
rect 15106 14952 15140 14986
rect 15174 14952 15290 14986
rect 12848 14940 15290 14952
rect 12848 14882 12906 14940
rect 12848 14848 12860 14882
rect 12894 14848 12906 14882
rect 15232 14882 15290 14940
rect 12848 14814 12906 14848
rect 12848 14780 12860 14814
rect 12894 14780 12906 14814
rect 12848 14746 12906 14780
rect 15232 14848 15244 14882
rect 15278 14848 15290 14882
rect 15232 14814 15290 14848
rect 15232 14780 15244 14814
rect 15278 14780 15290 14814
rect 12848 14712 12860 14746
rect 12894 14712 12906 14746
rect 12848 14678 12906 14712
rect 12848 14644 12860 14678
rect 12894 14644 12906 14678
rect 12848 14610 12906 14644
rect 12848 14576 12860 14610
rect 12894 14576 12906 14610
rect 12848 14542 12906 14576
rect 12848 14508 12860 14542
rect 12894 14508 12906 14542
rect 12848 14474 12906 14508
rect 12848 14440 12860 14474
rect 12894 14440 12906 14474
rect 12848 14406 12906 14440
rect 12848 14372 12860 14406
rect 12894 14372 12906 14406
rect 12848 14338 12906 14372
rect 12848 14304 12860 14338
rect 12894 14304 12906 14338
rect 12848 14270 12906 14304
rect 12848 14236 12860 14270
rect 12894 14236 12906 14270
rect 12848 14202 12906 14236
rect 12848 14168 12860 14202
rect 12894 14168 12906 14202
rect 12848 14134 12906 14168
rect 12848 14100 12860 14134
rect 12894 14100 12906 14134
rect 12848 14066 12906 14100
rect 12848 14032 12860 14066
rect 12894 14032 12906 14066
rect 12848 13998 12906 14032
rect 12848 13964 12860 13998
rect 12894 13964 12906 13998
rect 12848 13930 12906 13964
rect 12848 13896 12860 13930
rect 12894 13896 12906 13930
rect 12848 13862 12906 13896
rect 12848 13828 12860 13862
rect 12894 13828 12906 13862
rect 12848 13794 12906 13828
rect 12848 13760 12860 13794
rect 12894 13760 12906 13794
rect 12848 13726 12906 13760
rect 12848 13692 12860 13726
rect 12894 13692 12906 13726
rect 12848 13658 12906 13692
rect 12848 13624 12860 13658
rect 12894 13624 12906 13658
rect 12848 13590 12906 13624
rect 12848 13556 12860 13590
rect 12894 13556 12906 13590
rect 12848 13522 12906 13556
rect 12848 13488 12860 13522
rect 12894 13488 12906 13522
rect 12848 13454 12906 13488
rect 12848 13420 12860 13454
rect 12894 13420 12906 13454
rect 12848 13386 12906 13420
rect 12848 13352 12860 13386
rect 12894 13352 12906 13386
rect 12848 13318 12906 13352
rect 12848 13284 12860 13318
rect 12894 13284 12906 13318
rect 12848 13250 12906 13284
rect 12848 13216 12860 13250
rect 12894 13216 12906 13250
rect 12848 13182 12906 13216
rect 12848 13148 12860 13182
rect 12894 13148 12906 13182
rect 12848 13114 12906 13148
rect 12848 13080 12860 13114
rect 12894 13080 12906 13114
rect 12848 13046 12906 13080
rect 12848 13012 12860 13046
rect 12894 13012 12906 13046
rect 12848 12978 12906 13012
rect 12848 12944 12860 12978
rect 12894 12944 12906 12978
rect 12848 12910 12906 12944
rect 12848 12876 12860 12910
rect 12894 12876 12906 12910
rect 12848 12842 12906 12876
rect 12848 12808 12860 12842
rect 12894 12808 12906 12842
rect 12848 12774 12906 12808
rect 12848 12740 12860 12774
rect 12894 12740 12906 12774
rect 12848 12706 12906 12740
rect 12848 12672 12860 12706
rect 12894 12672 12906 12706
rect 12848 12638 12906 12672
rect 12848 12604 12860 12638
rect 12894 12604 12906 12638
rect 12848 12570 12906 12604
rect 12848 12536 12860 12570
rect 12894 12536 12906 12570
rect 12848 12502 12906 12536
rect 12848 12468 12860 12502
rect 12894 12468 12906 12502
rect 12848 12434 12906 12468
rect 12848 12400 12860 12434
rect 12894 12400 12906 12434
rect 12848 12366 12906 12400
rect 12848 12332 12860 12366
rect 12894 12332 12906 12366
rect 12848 12298 12906 12332
rect 12848 12264 12860 12298
rect 12894 12264 12906 12298
rect 12848 12230 12906 12264
rect 12848 12196 12860 12230
rect 12894 12196 12906 12230
rect 12848 12162 12906 12196
rect 12848 12128 12860 12162
rect 12894 12128 12906 12162
rect 12848 12094 12906 12128
rect 12848 12060 12860 12094
rect 12894 12060 12906 12094
rect 12848 12026 12906 12060
rect 12848 11992 12860 12026
rect 12894 11992 12906 12026
rect 12848 11958 12906 11992
rect 12848 11924 12860 11958
rect 12894 11924 12906 11958
rect 12848 11890 12906 11924
rect 12848 11856 12860 11890
rect 12894 11856 12906 11890
rect 12848 11822 12906 11856
rect 12848 11788 12860 11822
rect 12894 11788 12906 11822
rect 12848 11754 12906 11788
rect 15232 14746 15290 14780
rect 15232 14712 15244 14746
rect 15278 14712 15290 14746
rect 15232 14678 15290 14712
rect 15232 14644 15244 14678
rect 15278 14644 15290 14678
rect 15232 14610 15290 14644
rect 15232 14576 15244 14610
rect 15278 14576 15290 14610
rect 15232 14542 15290 14576
rect 15232 14508 15244 14542
rect 15278 14508 15290 14542
rect 15232 14474 15290 14508
rect 15232 14440 15244 14474
rect 15278 14440 15290 14474
rect 15232 14406 15290 14440
rect 15232 14372 15244 14406
rect 15278 14372 15290 14406
rect 15232 14338 15290 14372
rect 15232 14304 15244 14338
rect 15278 14304 15290 14338
rect 15232 14270 15290 14304
rect 15232 14236 15244 14270
rect 15278 14236 15290 14270
rect 15232 14202 15290 14236
rect 15232 14168 15244 14202
rect 15278 14168 15290 14202
rect 15232 14134 15290 14168
rect 15232 14100 15244 14134
rect 15278 14100 15290 14134
rect 15232 14066 15290 14100
rect 15232 14032 15244 14066
rect 15278 14032 15290 14066
rect 15232 13998 15290 14032
rect 15232 13964 15244 13998
rect 15278 13964 15290 13998
rect 15232 13930 15290 13964
rect 15232 13896 15244 13930
rect 15278 13896 15290 13930
rect 15232 13862 15290 13896
rect 15232 13828 15244 13862
rect 15278 13828 15290 13862
rect 15232 13794 15290 13828
rect 15232 13760 15244 13794
rect 15278 13760 15290 13794
rect 15232 13726 15290 13760
rect 15232 13692 15244 13726
rect 15278 13692 15290 13726
rect 15232 13658 15290 13692
rect 15232 13624 15244 13658
rect 15278 13624 15290 13658
rect 15232 13590 15290 13624
rect 15232 13556 15244 13590
rect 15278 13556 15290 13590
rect 15232 13522 15290 13556
rect 15232 13488 15244 13522
rect 15278 13488 15290 13522
rect 15232 13454 15290 13488
rect 15232 13420 15244 13454
rect 15278 13420 15290 13454
rect 15232 13386 15290 13420
rect 15232 13352 15244 13386
rect 15278 13352 15290 13386
rect 15232 13318 15290 13352
rect 15232 13284 15244 13318
rect 15278 13284 15290 13318
rect 15232 13250 15290 13284
rect 15232 13216 15244 13250
rect 15278 13216 15290 13250
rect 15232 13182 15290 13216
rect 15232 13148 15244 13182
rect 15278 13148 15290 13182
rect 15232 13114 15290 13148
rect 15232 13080 15244 13114
rect 15278 13080 15290 13114
rect 15232 13046 15290 13080
rect 15232 13012 15244 13046
rect 15278 13012 15290 13046
rect 15232 12978 15290 13012
rect 15232 12944 15244 12978
rect 15278 12944 15290 12978
rect 15232 12910 15290 12944
rect 15232 12876 15244 12910
rect 15278 12876 15290 12910
rect 15232 12842 15290 12876
rect 15232 12808 15244 12842
rect 15278 12808 15290 12842
rect 15232 12774 15290 12808
rect 15232 12740 15244 12774
rect 15278 12740 15290 12774
rect 15232 12706 15290 12740
rect 15232 12672 15244 12706
rect 15278 12672 15290 12706
rect 15232 12638 15290 12672
rect 15232 12604 15244 12638
rect 15278 12604 15290 12638
rect 15232 12570 15290 12604
rect 15232 12536 15244 12570
rect 15278 12536 15290 12570
rect 15232 12502 15290 12536
rect 15232 12468 15244 12502
rect 15278 12468 15290 12502
rect 15232 12434 15290 12468
rect 15232 12400 15244 12434
rect 15278 12400 15290 12434
rect 15232 12366 15290 12400
rect 15232 12332 15244 12366
rect 15278 12332 15290 12366
rect 15232 12298 15290 12332
rect 15232 12264 15244 12298
rect 15278 12264 15290 12298
rect 15232 12230 15290 12264
rect 15232 12196 15244 12230
rect 15278 12196 15290 12230
rect 15232 12162 15290 12196
rect 15232 12128 15244 12162
rect 15278 12128 15290 12162
rect 15232 12094 15290 12128
rect 15232 12060 15244 12094
rect 15278 12060 15290 12094
rect 15232 12026 15290 12060
rect 15232 11992 15244 12026
rect 15278 11992 15290 12026
rect 15232 11958 15290 11992
rect 15232 11924 15244 11958
rect 15278 11924 15290 11958
rect 15232 11890 15290 11924
rect 15232 11856 15244 11890
rect 15278 11856 15290 11890
rect 15232 11822 15290 11856
rect 15232 11788 15244 11822
rect 15278 11788 15290 11822
rect 12848 11720 12860 11754
rect 12894 11720 12906 11754
rect 12848 11686 12906 11720
rect 12848 11652 12860 11686
rect 12894 11652 12906 11686
rect 15232 11754 15290 11788
rect 15232 11720 15244 11754
rect 15278 11720 15290 11754
rect 15232 11686 15290 11720
rect 12848 11594 12906 11652
rect 15232 11652 15244 11686
rect 15278 11652 15290 11686
rect 15232 11594 15290 11652
rect 12848 11582 15290 11594
rect 12848 11548 12964 11582
rect 12998 11548 13032 11582
rect 13066 11548 13100 11582
rect 13134 11548 13168 11582
rect 13202 11548 13236 11582
rect 13270 11548 13304 11582
rect 13338 11548 13372 11582
rect 13406 11548 13440 11582
rect 13474 11548 13508 11582
rect 13542 11548 13576 11582
rect 13610 11548 13644 11582
rect 13678 11548 13712 11582
rect 13746 11548 13780 11582
rect 13814 11548 13848 11582
rect 13882 11548 13916 11582
rect 13950 11548 13984 11582
rect 14018 11548 14052 11582
rect 14086 11548 14120 11582
rect 14154 11548 14188 11582
rect 14222 11548 14256 11582
rect 14290 11548 14324 11582
rect 14358 11548 14392 11582
rect 14426 11548 14460 11582
rect 14494 11548 14528 11582
rect 14562 11548 14596 11582
rect 14630 11548 14664 11582
rect 14698 11548 14732 11582
rect 14766 11548 14800 11582
rect 14834 11548 14868 11582
rect 14902 11548 14936 11582
rect 14970 11548 15004 11582
rect 15038 11548 15072 11582
rect 15106 11548 15140 11582
rect 15174 11548 15290 11582
rect 12848 11536 15290 11548
rect 15418 14986 16802 14998
rect 15418 14952 15549 14986
rect 15583 14952 15617 14986
rect 15651 14952 15685 14986
rect 15719 14952 15753 14986
rect 15787 14952 15821 14986
rect 15855 14952 15889 14986
rect 15923 14952 15957 14986
rect 15991 14952 16025 14986
rect 16059 14952 16093 14986
rect 16127 14952 16161 14986
rect 16195 14952 16229 14986
rect 16263 14952 16297 14986
rect 16331 14952 16365 14986
rect 16399 14952 16433 14986
rect 16467 14952 16501 14986
rect 16535 14952 16569 14986
rect 16603 14952 16637 14986
rect 16671 14952 16802 14986
rect 15418 14940 16802 14952
rect 15418 14882 15476 14940
rect 15418 14848 15430 14882
rect 15464 14848 15476 14882
rect 16744 14882 16802 14940
rect 15418 14814 15476 14848
rect 15418 14780 15430 14814
rect 15464 14780 15476 14814
rect 15418 14746 15476 14780
rect 16744 14848 16756 14882
rect 16790 14848 16802 14882
rect 16744 14814 16802 14848
rect 16744 14780 16756 14814
rect 16790 14780 16802 14814
rect 15418 14712 15430 14746
rect 15464 14712 15476 14746
rect 15418 14678 15476 14712
rect 15418 14644 15430 14678
rect 15464 14644 15476 14678
rect 15418 14610 15476 14644
rect 15418 14576 15430 14610
rect 15464 14576 15476 14610
rect 15418 14542 15476 14576
rect 15418 14508 15430 14542
rect 15464 14508 15476 14542
rect 15418 14474 15476 14508
rect 15418 14440 15430 14474
rect 15464 14440 15476 14474
rect 15418 14406 15476 14440
rect 15418 14372 15430 14406
rect 15464 14372 15476 14406
rect 15418 14338 15476 14372
rect 15418 14304 15430 14338
rect 15464 14304 15476 14338
rect 15418 14270 15476 14304
rect 15418 14236 15430 14270
rect 15464 14236 15476 14270
rect 15418 14202 15476 14236
rect 15418 14168 15430 14202
rect 15464 14168 15476 14202
rect 15418 14134 15476 14168
rect 15418 14100 15430 14134
rect 15464 14100 15476 14134
rect 15418 14066 15476 14100
rect 15418 14032 15430 14066
rect 15464 14032 15476 14066
rect 15418 13998 15476 14032
rect 15418 13964 15430 13998
rect 15464 13964 15476 13998
rect 15418 13930 15476 13964
rect 15418 13896 15430 13930
rect 15464 13896 15476 13930
rect 15418 13862 15476 13896
rect 15418 13828 15430 13862
rect 15464 13828 15476 13862
rect 15418 13794 15476 13828
rect 15418 13760 15430 13794
rect 15464 13760 15476 13794
rect 15418 13726 15476 13760
rect 15418 13692 15430 13726
rect 15464 13692 15476 13726
rect 15418 13658 15476 13692
rect 15418 13624 15430 13658
rect 15464 13624 15476 13658
rect 15418 13590 15476 13624
rect 15418 13556 15430 13590
rect 15464 13556 15476 13590
rect 15418 13522 15476 13556
rect 15418 13488 15430 13522
rect 15464 13488 15476 13522
rect 15418 13454 15476 13488
rect 15418 13420 15430 13454
rect 15464 13420 15476 13454
rect 15418 13386 15476 13420
rect 15418 13352 15430 13386
rect 15464 13352 15476 13386
rect 15418 13318 15476 13352
rect 15418 13284 15430 13318
rect 15464 13284 15476 13318
rect 15418 13250 15476 13284
rect 15418 13216 15430 13250
rect 15464 13216 15476 13250
rect 15418 13182 15476 13216
rect 15418 13148 15430 13182
rect 15464 13148 15476 13182
rect 15418 13114 15476 13148
rect 15418 13080 15430 13114
rect 15464 13080 15476 13114
rect 15418 13046 15476 13080
rect 15418 13012 15430 13046
rect 15464 13012 15476 13046
rect 15418 12978 15476 13012
rect 15418 12944 15430 12978
rect 15464 12944 15476 12978
rect 15418 12910 15476 12944
rect 15418 12876 15430 12910
rect 15464 12876 15476 12910
rect 15418 12842 15476 12876
rect 15418 12808 15430 12842
rect 15464 12808 15476 12842
rect 15418 12774 15476 12808
rect 15418 12740 15430 12774
rect 15464 12740 15476 12774
rect 15418 12706 15476 12740
rect 15418 12672 15430 12706
rect 15464 12672 15476 12706
rect 15418 12638 15476 12672
rect 15418 12604 15430 12638
rect 15464 12604 15476 12638
rect 15418 12570 15476 12604
rect 15418 12536 15430 12570
rect 15464 12536 15476 12570
rect 15418 12502 15476 12536
rect 15418 12468 15430 12502
rect 15464 12468 15476 12502
rect 15418 12434 15476 12468
rect 15418 12400 15430 12434
rect 15464 12400 15476 12434
rect 15418 12366 15476 12400
rect 15418 12332 15430 12366
rect 15464 12332 15476 12366
rect 15418 12298 15476 12332
rect 15418 12264 15430 12298
rect 15464 12264 15476 12298
rect 15418 12230 15476 12264
rect 15418 12196 15430 12230
rect 15464 12196 15476 12230
rect 15418 12162 15476 12196
rect 15418 12128 15430 12162
rect 15464 12128 15476 12162
rect 15418 12094 15476 12128
rect 15418 12060 15430 12094
rect 15464 12060 15476 12094
rect 15418 12026 15476 12060
rect 15418 11992 15430 12026
rect 15464 11992 15476 12026
rect 15418 11958 15476 11992
rect 15418 11924 15430 11958
rect 15464 11924 15476 11958
rect 15418 11890 15476 11924
rect 15418 11856 15430 11890
rect 15464 11856 15476 11890
rect 15418 11822 15476 11856
rect 15418 11788 15430 11822
rect 15464 11788 15476 11822
rect 15418 11754 15476 11788
rect 16744 14746 16802 14780
rect 16744 14712 16756 14746
rect 16790 14712 16802 14746
rect 16744 14678 16802 14712
rect 16744 14644 16756 14678
rect 16790 14644 16802 14678
rect 16744 14610 16802 14644
rect 16744 14576 16756 14610
rect 16790 14576 16802 14610
rect 16744 14542 16802 14576
rect 16744 14508 16756 14542
rect 16790 14508 16802 14542
rect 16744 14474 16802 14508
rect 16744 14440 16756 14474
rect 16790 14440 16802 14474
rect 16744 14406 16802 14440
rect 16744 14372 16756 14406
rect 16790 14372 16802 14406
rect 16744 14338 16802 14372
rect 16744 14304 16756 14338
rect 16790 14304 16802 14338
rect 16744 14270 16802 14304
rect 16744 14236 16756 14270
rect 16790 14236 16802 14270
rect 16744 14202 16802 14236
rect 16744 14168 16756 14202
rect 16790 14168 16802 14202
rect 16744 14134 16802 14168
rect 16744 14100 16756 14134
rect 16790 14100 16802 14134
rect 16744 14066 16802 14100
rect 16744 14032 16756 14066
rect 16790 14032 16802 14066
rect 16744 13998 16802 14032
rect 16744 13964 16756 13998
rect 16790 13964 16802 13998
rect 16744 13930 16802 13964
rect 16744 13896 16756 13930
rect 16790 13896 16802 13930
rect 16744 13862 16802 13896
rect 16744 13828 16756 13862
rect 16790 13828 16802 13862
rect 16744 13794 16802 13828
rect 16744 13760 16756 13794
rect 16790 13760 16802 13794
rect 16744 13726 16802 13760
rect 16744 13692 16756 13726
rect 16790 13692 16802 13726
rect 16744 13658 16802 13692
rect 16744 13624 16756 13658
rect 16790 13624 16802 13658
rect 16744 13590 16802 13624
rect 16744 13556 16756 13590
rect 16790 13556 16802 13590
rect 16744 13522 16802 13556
rect 16744 13488 16756 13522
rect 16790 13488 16802 13522
rect 16744 13454 16802 13488
rect 16744 13420 16756 13454
rect 16790 13420 16802 13454
rect 16744 13386 16802 13420
rect 16744 13352 16756 13386
rect 16790 13352 16802 13386
rect 16744 13318 16802 13352
rect 16744 13284 16756 13318
rect 16790 13284 16802 13318
rect 16744 13250 16802 13284
rect 16744 13216 16756 13250
rect 16790 13216 16802 13250
rect 16744 13182 16802 13216
rect 16744 13148 16756 13182
rect 16790 13148 16802 13182
rect 16744 13114 16802 13148
rect 16744 13080 16756 13114
rect 16790 13080 16802 13114
rect 16744 13046 16802 13080
rect 16744 13012 16756 13046
rect 16790 13012 16802 13046
rect 16744 12978 16802 13012
rect 16744 12944 16756 12978
rect 16790 12944 16802 12978
rect 16744 12910 16802 12944
rect 16744 12876 16756 12910
rect 16790 12876 16802 12910
rect 16744 12842 16802 12876
rect 16744 12808 16756 12842
rect 16790 12808 16802 12842
rect 16744 12774 16802 12808
rect 16744 12740 16756 12774
rect 16790 12740 16802 12774
rect 16744 12706 16802 12740
rect 16744 12672 16756 12706
rect 16790 12672 16802 12706
rect 16744 12638 16802 12672
rect 16744 12604 16756 12638
rect 16790 12604 16802 12638
rect 16744 12570 16802 12604
rect 16744 12536 16756 12570
rect 16790 12536 16802 12570
rect 16744 12502 16802 12536
rect 16744 12468 16756 12502
rect 16790 12468 16802 12502
rect 16744 12434 16802 12468
rect 16744 12400 16756 12434
rect 16790 12400 16802 12434
rect 16744 12366 16802 12400
rect 16744 12332 16756 12366
rect 16790 12332 16802 12366
rect 16744 12298 16802 12332
rect 16744 12264 16756 12298
rect 16790 12264 16802 12298
rect 16744 12230 16802 12264
rect 16744 12196 16756 12230
rect 16790 12196 16802 12230
rect 16744 12162 16802 12196
rect 16744 12128 16756 12162
rect 16790 12128 16802 12162
rect 16744 12094 16802 12128
rect 16744 12060 16756 12094
rect 16790 12060 16802 12094
rect 16744 12026 16802 12060
rect 16744 11992 16756 12026
rect 16790 11992 16802 12026
rect 16744 11958 16802 11992
rect 16744 11924 16756 11958
rect 16790 11924 16802 11958
rect 16744 11890 16802 11924
rect 16744 11856 16756 11890
rect 16790 11856 16802 11890
rect 16744 11822 16802 11856
rect 16744 11788 16756 11822
rect 16790 11788 16802 11822
rect 15418 11720 15430 11754
rect 15464 11720 15476 11754
rect 15418 11686 15476 11720
rect 15418 11652 15430 11686
rect 15464 11652 15476 11686
rect 16744 11754 16802 11788
rect 16744 11720 16756 11754
rect 16790 11720 16802 11754
rect 16744 11686 16802 11720
rect 15418 11594 15476 11652
rect 16744 11652 16756 11686
rect 16790 11652 16802 11686
rect 16744 11594 16802 11652
rect 15418 11582 16802 11594
rect 15418 11548 15549 11582
rect 15583 11548 15617 11582
rect 15651 11548 15685 11582
rect 15719 11548 15753 11582
rect 15787 11548 15821 11582
rect 15855 11548 15889 11582
rect 15923 11548 15957 11582
rect 15991 11548 16025 11582
rect 16059 11548 16093 11582
rect 16127 11548 16161 11582
rect 16195 11548 16229 11582
rect 16263 11548 16297 11582
rect 16331 11548 16365 11582
rect 16399 11548 16433 11582
rect 16467 11548 16501 11582
rect 16535 11548 16569 11582
rect 16603 11548 16637 11582
rect 16671 11548 16802 11582
rect 15418 11536 16802 11548
rect 16928 14996 18312 15008
rect 16928 14962 17059 14996
rect 17093 14962 17127 14996
rect 17161 14962 17195 14996
rect 17229 14962 17263 14996
rect 17297 14962 17331 14996
rect 17365 14962 17399 14996
rect 17433 14962 17467 14996
rect 17501 14962 17535 14996
rect 17569 14962 17603 14996
rect 17637 14962 17671 14996
rect 17705 14962 17739 14996
rect 17773 14962 17807 14996
rect 17841 14962 17875 14996
rect 17909 14962 17943 14996
rect 17977 14962 18011 14996
rect 18045 14962 18079 14996
rect 18113 14962 18147 14996
rect 18181 14962 18312 14996
rect 16928 14950 18312 14962
rect 16928 14892 16986 14950
rect 16928 14858 16940 14892
rect 16974 14858 16986 14892
rect 18254 14892 18312 14950
rect 16928 14824 16986 14858
rect 16928 14790 16940 14824
rect 16974 14790 16986 14824
rect 16928 14756 16986 14790
rect 18254 14858 18266 14892
rect 18300 14858 18312 14892
rect 18254 14824 18312 14858
rect 18254 14790 18266 14824
rect 18300 14790 18312 14824
rect 16928 14722 16940 14756
rect 16974 14722 16986 14756
rect 16928 14688 16986 14722
rect 16928 14654 16940 14688
rect 16974 14654 16986 14688
rect 16928 14620 16986 14654
rect 16928 14586 16940 14620
rect 16974 14586 16986 14620
rect 16928 14552 16986 14586
rect 16928 14518 16940 14552
rect 16974 14518 16986 14552
rect 16928 14484 16986 14518
rect 16928 14450 16940 14484
rect 16974 14450 16986 14484
rect 16928 14416 16986 14450
rect 16928 14382 16940 14416
rect 16974 14382 16986 14416
rect 16928 14348 16986 14382
rect 16928 14314 16940 14348
rect 16974 14314 16986 14348
rect 16928 14280 16986 14314
rect 16928 14246 16940 14280
rect 16974 14246 16986 14280
rect 16928 14212 16986 14246
rect 16928 14178 16940 14212
rect 16974 14178 16986 14212
rect 16928 14144 16986 14178
rect 16928 14110 16940 14144
rect 16974 14110 16986 14144
rect 16928 14076 16986 14110
rect 16928 14042 16940 14076
rect 16974 14042 16986 14076
rect 16928 14008 16986 14042
rect 16928 13974 16940 14008
rect 16974 13974 16986 14008
rect 16928 13940 16986 13974
rect 16928 13906 16940 13940
rect 16974 13906 16986 13940
rect 16928 13872 16986 13906
rect 16928 13838 16940 13872
rect 16974 13838 16986 13872
rect 16928 13804 16986 13838
rect 16928 13770 16940 13804
rect 16974 13770 16986 13804
rect 16928 13736 16986 13770
rect 16928 13702 16940 13736
rect 16974 13702 16986 13736
rect 16928 13668 16986 13702
rect 16928 13634 16940 13668
rect 16974 13634 16986 13668
rect 16928 13600 16986 13634
rect 16928 13566 16940 13600
rect 16974 13566 16986 13600
rect 16928 13532 16986 13566
rect 16928 13498 16940 13532
rect 16974 13498 16986 13532
rect 16928 13464 16986 13498
rect 16928 13430 16940 13464
rect 16974 13430 16986 13464
rect 16928 13396 16986 13430
rect 16928 13362 16940 13396
rect 16974 13362 16986 13396
rect 16928 13328 16986 13362
rect 16928 13294 16940 13328
rect 16974 13294 16986 13328
rect 16928 13260 16986 13294
rect 16928 13226 16940 13260
rect 16974 13226 16986 13260
rect 16928 13192 16986 13226
rect 16928 13158 16940 13192
rect 16974 13158 16986 13192
rect 16928 13124 16986 13158
rect 16928 13090 16940 13124
rect 16974 13090 16986 13124
rect 16928 13056 16986 13090
rect 16928 13022 16940 13056
rect 16974 13022 16986 13056
rect 16928 12988 16986 13022
rect 16928 12954 16940 12988
rect 16974 12954 16986 12988
rect 16928 12920 16986 12954
rect 16928 12886 16940 12920
rect 16974 12886 16986 12920
rect 16928 12852 16986 12886
rect 16928 12818 16940 12852
rect 16974 12818 16986 12852
rect 16928 12784 16986 12818
rect 16928 12750 16940 12784
rect 16974 12750 16986 12784
rect 16928 12716 16986 12750
rect 16928 12682 16940 12716
rect 16974 12682 16986 12716
rect 16928 12648 16986 12682
rect 16928 12614 16940 12648
rect 16974 12614 16986 12648
rect 16928 12580 16986 12614
rect 16928 12546 16940 12580
rect 16974 12546 16986 12580
rect 16928 12512 16986 12546
rect 16928 12478 16940 12512
rect 16974 12478 16986 12512
rect 16928 12444 16986 12478
rect 16928 12410 16940 12444
rect 16974 12410 16986 12444
rect 16928 12376 16986 12410
rect 16928 12342 16940 12376
rect 16974 12342 16986 12376
rect 16928 12308 16986 12342
rect 16928 12274 16940 12308
rect 16974 12274 16986 12308
rect 16928 12240 16986 12274
rect 16928 12206 16940 12240
rect 16974 12206 16986 12240
rect 16928 12172 16986 12206
rect 16928 12138 16940 12172
rect 16974 12138 16986 12172
rect 16928 12104 16986 12138
rect 16928 12070 16940 12104
rect 16974 12070 16986 12104
rect 16928 12036 16986 12070
rect 16928 12002 16940 12036
rect 16974 12002 16986 12036
rect 16928 11968 16986 12002
rect 16928 11934 16940 11968
rect 16974 11934 16986 11968
rect 16928 11900 16986 11934
rect 16928 11866 16940 11900
rect 16974 11866 16986 11900
rect 16928 11832 16986 11866
rect 16928 11798 16940 11832
rect 16974 11798 16986 11832
rect 16928 11764 16986 11798
rect 18254 14756 18312 14790
rect 18254 14722 18266 14756
rect 18300 14722 18312 14756
rect 18254 14688 18312 14722
rect 18254 14654 18266 14688
rect 18300 14654 18312 14688
rect 18254 14620 18312 14654
rect 18254 14586 18266 14620
rect 18300 14586 18312 14620
rect 18254 14552 18312 14586
rect 18254 14518 18266 14552
rect 18300 14518 18312 14552
rect 18254 14484 18312 14518
rect 18254 14450 18266 14484
rect 18300 14450 18312 14484
rect 18254 14416 18312 14450
rect 18254 14382 18266 14416
rect 18300 14382 18312 14416
rect 18254 14348 18312 14382
rect 18254 14314 18266 14348
rect 18300 14314 18312 14348
rect 18254 14280 18312 14314
rect 18254 14246 18266 14280
rect 18300 14246 18312 14280
rect 18254 14212 18312 14246
rect 18254 14178 18266 14212
rect 18300 14178 18312 14212
rect 18254 14144 18312 14178
rect 18254 14110 18266 14144
rect 18300 14110 18312 14144
rect 18254 14076 18312 14110
rect 18254 14042 18266 14076
rect 18300 14042 18312 14076
rect 18254 14008 18312 14042
rect 18254 13974 18266 14008
rect 18300 13974 18312 14008
rect 18254 13940 18312 13974
rect 18254 13906 18266 13940
rect 18300 13906 18312 13940
rect 18254 13872 18312 13906
rect 18254 13838 18266 13872
rect 18300 13838 18312 13872
rect 18254 13804 18312 13838
rect 18254 13770 18266 13804
rect 18300 13770 18312 13804
rect 18254 13736 18312 13770
rect 18254 13702 18266 13736
rect 18300 13702 18312 13736
rect 18254 13668 18312 13702
rect 18254 13634 18266 13668
rect 18300 13634 18312 13668
rect 18254 13600 18312 13634
rect 18254 13566 18266 13600
rect 18300 13566 18312 13600
rect 18254 13532 18312 13566
rect 18254 13498 18266 13532
rect 18300 13498 18312 13532
rect 18254 13464 18312 13498
rect 18254 13430 18266 13464
rect 18300 13430 18312 13464
rect 18254 13396 18312 13430
rect 18254 13362 18266 13396
rect 18300 13362 18312 13396
rect 18254 13328 18312 13362
rect 18254 13294 18266 13328
rect 18300 13294 18312 13328
rect 18254 13260 18312 13294
rect 18254 13226 18266 13260
rect 18300 13226 18312 13260
rect 18254 13192 18312 13226
rect 18254 13158 18266 13192
rect 18300 13158 18312 13192
rect 18254 13124 18312 13158
rect 18254 13090 18266 13124
rect 18300 13090 18312 13124
rect 18254 13056 18312 13090
rect 18254 13022 18266 13056
rect 18300 13022 18312 13056
rect 18254 12988 18312 13022
rect 18254 12954 18266 12988
rect 18300 12954 18312 12988
rect 18254 12920 18312 12954
rect 18254 12886 18266 12920
rect 18300 12886 18312 12920
rect 18254 12852 18312 12886
rect 18254 12818 18266 12852
rect 18300 12818 18312 12852
rect 18254 12784 18312 12818
rect 18254 12750 18266 12784
rect 18300 12750 18312 12784
rect 18254 12716 18312 12750
rect 18254 12682 18266 12716
rect 18300 12682 18312 12716
rect 18254 12648 18312 12682
rect 18254 12614 18266 12648
rect 18300 12614 18312 12648
rect 18254 12580 18312 12614
rect 18254 12546 18266 12580
rect 18300 12546 18312 12580
rect 18254 12512 18312 12546
rect 18254 12478 18266 12512
rect 18300 12478 18312 12512
rect 18254 12444 18312 12478
rect 18254 12410 18266 12444
rect 18300 12410 18312 12444
rect 18254 12376 18312 12410
rect 18254 12342 18266 12376
rect 18300 12342 18312 12376
rect 18254 12308 18312 12342
rect 18254 12274 18266 12308
rect 18300 12274 18312 12308
rect 18254 12240 18312 12274
rect 18254 12206 18266 12240
rect 18300 12206 18312 12240
rect 18254 12172 18312 12206
rect 18254 12138 18266 12172
rect 18300 12138 18312 12172
rect 18254 12104 18312 12138
rect 18254 12070 18266 12104
rect 18300 12070 18312 12104
rect 18254 12036 18312 12070
rect 18254 12002 18266 12036
rect 18300 12002 18312 12036
rect 18254 11968 18312 12002
rect 18254 11934 18266 11968
rect 18300 11934 18312 11968
rect 18254 11900 18312 11934
rect 18254 11866 18266 11900
rect 18300 11866 18312 11900
rect 18254 11832 18312 11866
rect 18254 11798 18266 11832
rect 18300 11798 18312 11832
rect 16928 11730 16940 11764
rect 16974 11730 16986 11764
rect 16928 11696 16986 11730
rect 16928 11662 16940 11696
rect 16974 11662 16986 11696
rect 18254 11764 18312 11798
rect 18254 11730 18266 11764
rect 18300 11730 18312 11764
rect 18254 11696 18312 11730
rect 16928 11604 16986 11662
rect 18254 11662 18266 11696
rect 18300 11662 18312 11696
rect 18254 11604 18312 11662
rect 16928 11592 18312 11604
rect 16928 11558 17059 11592
rect 17093 11558 17127 11592
rect 17161 11558 17195 11592
rect 17229 11558 17263 11592
rect 17297 11558 17331 11592
rect 17365 11558 17399 11592
rect 17433 11558 17467 11592
rect 17501 11558 17535 11592
rect 17569 11558 17603 11592
rect 17637 11558 17671 11592
rect 17705 11558 17739 11592
rect 17773 11558 17807 11592
rect 17841 11558 17875 11592
rect 17909 11558 17943 11592
rect 17977 11558 18011 11592
rect 18045 11558 18079 11592
rect 18113 11558 18147 11592
rect 18181 11558 18312 11592
rect 16928 11546 18312 11558
rect 18392 14980 19776 14992
rect 18392 14946 18523 14980
rect 18557 14946 18591 14980
rect 18625 14946 18659 14980
rect 18693 14946 18727 14980
rect 18761 14946 18795 14980
rect 18829 14946 18863 14980
rect 18897 14946 18931 14980
rect 18965 14946 18999 14980
rect 19033 14946 19067 14980
rect 19101 14946 19135 14980
rect 19169 14946 19203 14980
rect 19237 14946 19271 14980
rect 19305 14946 19339 14980
rect 19373 14946 19407 14980
rect 19441 14946 19475 14980
rect 19509 14946 19543 14980
rect 19577 14946 19611 14980
rect 19645 14946 19776 14980
rect 18392 14934 19776 14946
rect 18392 14876 18450 14934
rect 18392 14842 18404 14876
rect 18438 14842 18450 14876
rect 19718 14876 19776 14934
rect 18392 14808 18450 14842
rect 18392 14774 18404 14808
rect 18438 14774 18450 14808
rect 18392 14740 18450 14774
rect 19718 14842 19730 14876
rect 19764 14842 19776 14876
rect 19718 14808 19776 14842
rect 19718 14774 19730 14808
rect 19764 14774 19776 14808
rect 18392 14706 18404 14740
rect 18438 14706 18450 14740
rect 18392 14672 18450 14706
rect 18392 14638 18404 14672
rect 18438 14638 18450 14672
rect 18392 14604 18450 14638
rect 18392 14570 18404 14604
rect 18438 14570 18450 14604
rect 18392 14536 18450 14570
rect 18392 14502 18404 14536
rect 18438 14502 18450 14536
rect 18392 14468 18450 14502
rect 18392 14434 18404 14468
rect 18438 14434 18450 14468
rect 18392 14400 18450 14434
rect 18392 14366 18404 14400
rect 18438 14366 18450 14400
rect 18392 14332 18450 14366
rect 18392 14298 18404 14332
rect 18438 14298 18450 14332
rect 18392 14264 18450 14298
rect 18392 14230 18404 14264
rect 18438 14230 18450 14264
rect 18392 14196 18450 14230
rect 18392 14162 18404 14196
rect 18438 14162 18450 14196
rect 18392 14128 18450 14162
rect 18392 14094 18404 14128
rect 18438 14094 18450 14128
rect 18392 14060 18450 14094
rect 18392 14026 18404 14060
rect 18438 14026 18450 14060
rect 18392 13992 18450 14026
rect 18392 13958 18404 13992
rect 18438 13958 18450 13992
rect 18392 13924 18450 13958
rect 18392 13890 18404 13924
rect 18438 13890 18450 13924
rect 18392 13856 18450 13890
rect 18392 13822 18404 13856
rect 18438 13822 18450 13856
rect 18392 13788 18450 13822
rect 18392 13754 18404 13788
rect 18438 13754 18450 13788
rect 18392 13720 18450 13754
rect 18392 13686 18404 13720
rect 18438 13686 18450 13720
rect 18392 13652 18450 13686
rect 18392 13618 18404 13652
rect 18438 13618 18450 13652
rect 18392 13584 18450 13618
rect 18392 13550 18404 13584
rect 18438 13550 18450 13584
rect 18392 13516 18450 13550
rect 18392 13482 18404 13516
rect 18438 13482 18450 13516
rect 18392 13448 18450 13482
rect 18392 13414 18404 13448
rect 18438 13414 18450 13448
rect 18392 13380 18450 13414
rect 18392 13346 18404 13380
rect 18438 13346 18450 13380
rect 18392 13312 18450 13346
rect 18392 13278 18404 13312
rect 18438 13278 18450 13312
rect 18392 13244 18450 13278
rect 18392 13210 18404 13244
rect 18438 13210 18450 13244
rect 18392 13176 18450 13210
rect 18392 13142 18404 13176
rect 18438 13142 18450 13176
rect 18392 13108 18450 13142
rect 18392 13074 18404 13108
rect 18438 13074 18450 13108
rect 18392 13040 18450 13074
rect 18392 13006 18404 13040
rect 18438 13006 18450 13040
rect 18392 12972 18450 13006
rect 18392 12938 18404 12972
rect 18438 12938 18450 12972
rect 18392 12904 18450 12938
rect 18392 12870 18404 12904
rect 18438 12870 18450 12904
rect 18392 12836 18450 12870
rect 18392 12802 18404 12836
rect 18438 12802 18450 12836
rect 18392 12768 18450 12802
rect 18392 12734 18404 12768
rect 18438 12734 18450 12768
rect 18392 12700 18450 12734
rect 18392 12666 18404 12700
rect 18438 12666 18450 12700
rect 18392 12632 18450 12666
rect 18392 12598 18404 12632
rect 18438 12598 18450 12632
rect 18392 12564 18450 12598
rect 18392 12530 18404 12564
rect 18438 12530 18450 12564
rect 18392 12496 18450 12530
rect 18392 12462 18404 12496
rect 18438 12462 18450 12496
rect 18392 12428 18450 12462
rect 18392 12394 18404 12428
rect 18438 12394 18450 12428
rect 18392 12360 18450 12394
rect 18392 12326 18404 12360
rect 18438 12326 18450 12360
rect 18392 12292 18450 12326
rect 18392 12258 18404 12292
rect 18438 12258 18450 12292
rect 18392 12224 18450 12258
rect 18392 12190 18404 12224
rect 18438 12190 18450 12224
rect 18392 12156 18450 12190
rect 18392 12122 18404 12156
rect 18438 12122 18450 12156
rect 18392 12088 18450 12122
rect 18392 12054 18404 12088
rect 18438 12054 18450 12088
rect 18392 12020 18450 12054
rect 18392 11986 18404 12020
rect 18438 11986 18450 12020
rect 18392 11952 18450 11986
rect 18392 11918 18404 11952
rect 18438 11918 18450 11952
rect 18392 11884 18450 11918
rect 18392 11850 18404 11884
rect 18438 11850 18450 11884
rect 18392 11816 18450 11850
rect 18392 11782 18404 11816
rect 18438 11782 18450 11816
rect 18392 11748 18450 11782
rect 19718 14740 19776 14774
rect 19718 14706 19730 14740
rect 19764 14706 19776 14740
rect 19718 14672 19776 14706
rect 19718 14638 19730 14672
rect 19764 14638 19776 14672
rect 19718 14604 19776 14638
rect 19718 14570 19730 14604
rect 19764 14570 19776 14604
rect 19718 14536 19776 14570
rect 19718 14502 19730 14536
rect 19764 14502 19776 14536
rect 19718 14468 19776 14502
rect 19718 14434 19730 14468
rect 19764 14434 19776 14468
rect 19718 14400 19776 14434
rect 19718 14366 19730 14400
rect 19764 14366 19776 14400
rect 19718 14332 19776 14366
rect 19718 14298 19730 14332
rect 19764 14298 19776 14332
rect 19718 14264 19776 14298
rect 19718 14230 19730 14264
rect 19764 14230 19776 14264
rect 19718 14196 19776 14230
rect 19718 14162 19730 14196
rect 19764 14162 19776 14196
rect 19718 14128 19776 14162
rect 19718 14094 19730 14128
rect 19764 14094 19776 14128
rect 19718 14060 19776 14094
rect 19718 14026 19730 14060
rect 19764 14026 19776 14060
rect 19718 13992 19776 14026
rect 19718 13958 19730 13992
rect 19764 13958 19776 13992
rect 19718 13924 19776 13958
rect 19718 13890 19730 13924
rect 19764 13890 19776 13924
rect 19718 13856 19776 13890
rect 19718 13822 19730 13856
rect 19764 13822 19776 13856
rect 19718 13788 19776 13822
rect 19718 13754 19730 13788
rect 19764 13754 19776 13788
rect 19718 13720 19776 13754
rect 19718 13686 19730 13720
rect 19764 13686 19776 13720
rect 19718 13652 19776 13686
rect 19718 13618 19730 13652
rect 19764 13618 19776 13652
rect 19718 13584 19776 13618
rect 19718 13550 19730 13584
rect 19764 13550 19776 13584
rect 19718 13516 19776 13550
rect 19718 13482 19730 13516
rect 19764 13482 19776 13516
rect 19718 13448 19776 13482
rect 19718 13414 19730 13448
rect 19764 13414 19776 13448
rect 19718 13380 19776 13414
rect 19718 13346 19730 13380
rect 19764 13346 19776 13380
rect 19718 13312 19776 13346
rect 19718 13278 19730 13312
rect 19764 13278 19776 13312
rect 19718 13244 19776 13278
rect 19718 13210 19730 13244
rect 19764 13210 19776 13244
rect 19718 13176 19776 13210
rect 19718 13142 19730 13176
rect 19764 13142 19776 13176
rect 19718 13108 19776 13142
rect 19718 13074 19730 13108
rect 19764 13074 19776 13108
rect 19718 13040 19776 13074
rect 19718 13006 19730 13040
rect 19764 13006 19776 13040
rect 19718 12972 19776 13006
rect 19718 12938 19730 12972
rect 19764 12938 19776 12972
rect 19718 12904 19776 12938
rect 19718 12870 19730 12904
rect 19764 12870 19776 12904
rect 19718 12836 19776 12870
rect 19718 12802 19730 12836
rect 19764 12802 19776 12836
rect 19718 12768 19776 12802
rect 19718 12734 19730 12768
rect 19764 12734 19776 12768
rect 19718 12700 19776 12734
rect 19718 12666 19730 12700
rect 19764 12666 19776 12700
rect 19718 12632 19776 12666
rect 19718 12598 19730 12632
rect 19764 12598 19776 12632
rect 19718 12564 19776 12598
rect 19718 12530 19730 12564
rect 19764 12530 19776 12564
rect 19718 12496 19776 12530
rect 19718 12462 19730 12496
rect 19764 12462 19776 12496
rect 19718 12428 19776 12462
rect 19718 12394 19730 12428
rect 19764 12394 19776 12428
rect 19718 12360 19776 12394
rect 19718 12326 19730 12360
rect 19764 12326 19776 12360
rect 19718 12292 19776 12326
rect 19718 12258 19730 12292
rect 19764 12258 19776 12292
rect 19718 12224 19776 12258
rect 19718 12190 19730 12224
rect 19764 12190 19776 12224
rect 19718 12156 19776 12190
rect 19718 12122 19730 12156
rect 19764 12122 19776 12156
rect 19718 12088 19776 12122
rect 19718 12054 19730 12088
rect 19764 12054 19776 12088
rect 19718 12020 19776 12054
rect 19718 11986 19730 12020
rect 19764 11986 19776 12020
rect 19718 11952 19776 11986
rect 19718 11918 19730 11952
rect 19764 11918 19776 11952
rect 19718 11884 19776 11918
rect 19718 11850 19730 11884
rect 19764 11850 19776 11884
rect 19718 11816 19776 11850
rect 19718 11782 19730 11816
rect 19764 11782 19776 11816
rect 18392 11714 18404 11748
rect 18438 11714 18450 11748
rect 18392 11680 18450 11714
rect 18392 11646 18404 11680
rect 18438 11646 18450 11680
rect 19718 11748 19776 11782
rect 19718 11714 19730 11748
rect 19764 11714 19776 11748
rect 19718 11680 19776 11714
rect 18392 11588 18450 11646
rect 19718 11646 19730 11680
rect 19764 11646 19776 11680
rect 19718 11588 19776 11646
rect 18392 11576 19776 11588
rect 18392 11542 18523 11576
rect 18557 11542 18591 11576
rect 18625 11542 18659 11576
rect 18693 11542 18727 11576
rect 18761 11542 18795 11576
rect 18829 11542 18863 11576
rect 18897 11542 18931 11576
rect 18965 11542 18999 11576
rect 19033 11542 19067 11576
rect 19101 11542 19135 11576
rect 19169 11542 19203 11576
rect 19237 11542 19271 11576
rect 19305 11542 19339 11576
rect 19373 11542 19407 11576
rect 19441 11542 19475 11576
rect 19509 11542 19543 11576
rect 19577 11542 19611 11576
rect 19645 11542 19776 11576
rect 18392 11530 19776 11542
rect 14808 11466 17250 11478
rect 14808 11432 14924 11466
rect 14958 11432 14992 11466
rect 15026 11432 15060 11466
rect 15094 11432 15128 11466
rect 15162 11432 15196 11466
rect 15230 11432 15264 11466
rect 15298 11432 15332 11466
rect 15366 11432 15400 11466
rect 15434 11432 15468 11466
rect 15502 11432 15536 11466
rect 15570 11432 15604 11466
rect 15638 11432 15672 11466
rect 15706 11432 15740 11466
rect 15774 11432 15808 11466
rect 15842 11432 15876 11466
rect 15910 11432 15944 11466
rect 15978 11432 16012 11466
rect 16046 11432 16080 11466
rect 16114 11432 16148 11466
rect 16182 11432 16216 11466
rect 16250 11432 16284 11466
rect 16318 11432 16352 11466
rect 16386 11432 16420 11466
rect 16454 11432 16488 11466
rect 16522 11432 16556 11466
rect 16590 11432 16624 11466
rect 16658 11432 16692 11466
rect 16726 11432 16760 11466
rect 16794 11432 16828 11466
rect 16862 11432 16896 11466
rect 16930 11432 16964 11466
rect 16998 11432 17032 11466
rect 17066 11432 17100 11466
rect 17134 11432 17250 11466
rect 14808 11420 17250 11432
rect 14808 11362 14866 11420
rect 14808 11328 14820 11362
rect 14854 11328 14866 11362
rect 17192 11362 17250 11420
rect 14808 11294 14866 11328
rect 14808 11260 14820 11294
rect 14854 11260 14866 11294
rect 14808 11226 14866 11260
rect 17192 11328 17204 11362
rect 17238 11328 17250 11362
rect 17192 11294 17250 11328
rect 17192 11260 17204 11294
rect 17238 11260 17250 11294
rect 14808 11192 14820 11226
rect 14854 11192 14866 11226
rect 14808 11158 14866 11192
rect 14808 11124 14820 11158
rect 14854 11124 14866 11158
rect 14808 11090 14866 11124
rect 14808 11056 14820 11090
rect 14854 11056 14866 11090
rect 14808 11022 14866 11056
rect 14808 10988 14820 11022
rect 14854 10988 14866 11022
rect 14808 10954 14866 10988
rect 14808 10920 14820 10954
rect 14854 10920 14866 10954
rect 14808 10886 14866 10920
rect 14808 10852 14820 10886
rect 14854 10852 14866 10886
rect 14808 10818 14866 10852
rect 14808 10784 14820 10818
rect 14854 10784 14866 10818
rect 14808 10750 14866 10784
rect 14808 10716 14820 10750
rect 14854 10716 14866 10750
rect 14808 10682 14866 10716
rect 14808 10648 14820 10682
rect 14854 10648 14866 10682
rect 14808 10614 14866 10648
rect 14808 10580 14820 10614
rect 14854 10580 14866 10614
rect 14808 10546 14866 10580
rect 14808 10512 14820 10546
rect 14854 10512 14866 10546
rect 14808 10478 14866 10512
rect 14808 10444 14820 10478
rect 14854 10444 14866 10478
rect 14808 10410 14866 10444
rect 14808 10376 14820 10410
rect 14854 10376 14866 10410
rect 14808 10342 14866 10376
rect 14808 10308 14820 10342
rect 14854 10308 14866 10342
rect 14808 10274 14866 10308
rect 14808 10240 14820 10274
rect 14854 10240 14866 10274
rect 14808 10206 14866 10240
rect 14808 10172 14820 10206
rect 14854 10172 14866 10206
rect 14808 10138 14866 10172
rect 14808 10104 14820 10138
rect 14854 10104 14866 10138
rect 14808 10070 14866 10104
rect 14808 10036 14820 10070
rect 14854 10036 14866 10070
rect 14808 10002 14866 10036
rect 14808 9968 14820 10002
rect 14854 9968 14866 10002
rect 14808 9934 14866 9968
rect 14808 9900 14820 9934
rect 14854 9900 14866 9934
rect 14808 9866 14866 9900
rect 14808 9832 14820 9866
rect 14854 9832 14866 9866
rect 14808 9798 14866 9832
rect 14808 9764 14820 9798
rect 14854 9764 14866 9798
rect 14808 9730 14866 9764
rect 14808 9696 14820 9730
rect 14854 9696 14866 9730
rect 14808 9662 14866 9696
rect 14808 9628 14820 9662
rect 14854 9628 14866 9662
rect 14808 9594 14866 9628
rect 14808 9560 14820 9594
rect 14854 9560 14866 9594
rect 14808 9526 14866 9560
rect 14808 9492 14820 9526
rect 14854 9492 14866 9526
rect 14808 9458 14866 9492
rect 14808 9424 14820 9458
rect 14854 9424 14866 9458
rect 14808 9390 14866 9424
rect 14808 9356 14820 9390
rect 14854 9356 14866 9390
rect 14808 9322 14866 9356
rect 14808 9288 14820 9322
rect 14854 9288 14866 9322
rect 14808 9254 14866 9288
rect 14808 9220 14820 9254
rect 14854 9220 14866 9254
rect 14808 9186 14866 9220
rect 14808 9152 14820 9186
rect 14854 9152 14866 9186
rect 14808 9118 14866 9152
rect 14808 9084 14820 9118
rect 14854 9084 14866 9118
rect 14808 9050 14866 9084
rect 14808 9016 14820 9050
rect 14854 9016 14866 9050
rect 14808 8982 14866 9016
rect 14808 8948 14820 8982
rect 14854 8948 14866 8982
rect 14808 8914 14866 8948
rect 14808 8880 14820 8914
rect 14854 8880 14866 8914
rect 14808 8846 14866 8880
rect 14808 8812 14820 8846
rect 14854 8812 14866 8846
rect 14808 8778 14866 8812
rect 14808 8744 14820 8778
rect 14854 8744 14866 8778
rect 14808 8710 14866 8744
rect 14808 8676 14820 8710
rect 14854 8676 14866 8710
rect 14808 8642 14866 8676
rect 14808 8608 14820 8642
rect 14854 8608 14866 8642
rect 14808 8574 14866 8608
rect 14808 8540 14820 8574
rect 14854 8540 14866 8574
rect 14808 8506 14866 8540
rect 14808 8472 14820 8506
rect 14854 8472 14866 8506
rect 14808 8438 14866 8472
rect 14808 8404 14820 8438
rect 14854 8404 14866 8438
rect 14808 8370 14866 8404
rect 14808 8336 14820 8370
rect 14854 8336 14866 8370
rect 14808 8302 14866 8336
rect 14808 8268 14820 8302
rect 14854 8268 14866 8302
rect 14808 8234 14866 8268
rect 17192 11226 17250 11260
rect 17192 11192 17204 11226
rect 17238 11192 17250 11226
rect 17192 11158 17250 11192
rect 17192 11124 17204 11158
rect 17238 11124 17250 11158
rect 17192 11090 17250 11124
rect 17192 11056 17204 11090
rect 17238 11056 17250 11090
rect 17192 11022 17250 11056
rect 17192 10988 17204 11022
rect 17238 10988 17250 11022
rect 17192 10954 17250 10988
rect 17192 10920 17204 10954
rect 17238 10920 17250 10954
rect 17192 10886 17250 10920
rect 17192 10852 17204 10886
rect 17238 10852 17250 10886
rect 17192 10818 17250 10852
rect 17192 10784 17204 10818
rect 17238 10784 17250 10818
rect 17192 10750 17250 10784
rect 17192 10716 17204 10750
rect 17238 10716 17250 10750
rect 17192 10682 17250 10716
rect 17192 10648 17204 10682
rect 17238 10648 17250 10682
rect 17192 10614 17250 10648
rect 17192 10580 17204 10614
rect 17238 10580 17250 10614
rect 17192 10546 17250 10580
rect 17192 10512 17204 10546
rect 17238 10512 17250 10546
rect 17192 10478 17250 10512
rect 17192 10444 17204 10478
rect 17238 10444 17250 10478
rect 17192 10410 17250 10444
rect 17192 10376 17204 10410
rect 17238 10376 17250 10410
rect 17192 10342 17250 10376
rect 17192 10308 17204 10342
rect 17238 10308 17250 10342
rect 17192 10274 17250 10308
rect 17192 10240 17204 10274
rect 17238 10240 17250 10274
rect 17192 10206 17250 10240
rect 17192 10172 17204 10206
rect 17238 10172 17250 10206
rect 17192 10138 17250 10172
rect 17192 10104 17204 10138
rect 17238 10104 17250 10138
rect 17192 10070 17250 10104
rect 17192 10036 17204 10070
rect 17238 10036 17250 10070
rect 17192 10002 17250 10036
rect 17192 9968 17204 10002
rect 17238 9968 17250 10002
rect 17192 9934 17250 9968
rect 17192 9900 17204 9934
rect 17238 9900 17250 9934
rect 17192 9866 17250 9900
rect 17192 9832 17204 9866
rect 17238 9832 17250 9866
rect 17192 9798 17250 9832
rect 17192 9764 17204 9798
rect 17238 9764 17250 9798
rect 17192 9730 17250 9764
rect 17192 9696 17204 9730
rect 17238 9696 17250 9730
rect 17192 9662 17250 9696
rect 17192 9628 17204 9662
rect 17238 9628 17250 9662
rect 17192 9594 17250 9628
rect 17192 9560 17204 9594
rect 17238 9560 17250 9594
rect 17192 9526 17250 9560
rect 17192 9492 17204 9526
rect 17238 9492 17250 9526
rect 17192 9458 17250 9492
rect 17192 9424 17204 9458
rect 17238 9424 17250 9458
rect 17192 9390 17250 9424
rect 17192 9356 17204 9390
rect 17238 9356 17250 9390
rect 17192 9322 17250 9356
rect 17192 9288 17204 9322
rect 17238 9288 17250 9322
rect 17192 9254 17250 9288
rect 17192 9220 17204 9254
rect 17238 9220 17250 9254
rect 17192 9186 17250 9220
rect 17192 9152 17204 9186
rect 17238 9152 17250 9186
rect 17192 9118 17250 9152
rect 17192 9084 17204 9118
rect 17238 9084 17250 9118
rect 17192 9050 17250 9084
rect 17192 9016 17204 9050
rect 17238 9016 17250 9050
rect 17192 8982 17250 9016
rect 17192 8948 17204 8982
rect 17238 8948 17250 8982
rect 17192 8914 17250 8948
rect 17192 8880 17204 8914
rect 17238 8880 17250 8914
rect 17192 8846 17250 8880
rect 17192 8812 17204 8846
rect 17238 8812 17250 8846
rect 17192 8778 17250 8812
rect 17192 8744 17204 8778
rect 17238 8744 17250 8778
rect 17192 8710 17250 8744
rect 17192 8676 17204 8710
rect 17238 8676 17250 8710
rect 17192 8642 17250 8676
rect 17192 8608 17204 8642
rect 17238 8608 17250 8642
rect 17192 8574 17250 8608
rect 17192 8540 17204 8574
rect 17238 8540 17250 8574
rect 17192 8506 17250 8540
rect 17192 8472 17204 8506
rect 17238 8472 17250 8506
rect 17192 8438 17250 8472
rect 17192 8404 17204 8438
rect 17238 8404 17250 8438
rect 17192 8370 17250 8404
rect 17192 8336 17204 8370
rect 17238 8336 17250 8370
rect 17192 8302 17250 8336
rect 17192 8268 17204 8302
rect 17238 8268 17250 8302
rect 14808 8200 14820 8234
rect 14854 8200 14866 8234
rect 14808 8166 14866 8200
rect 14808 8132 14820 8166
rect 14854 8132 14866 8166
rect 17192 8234 17250 8268
rect 17192 8200 17204 8234
rect 17238 8200 17250 8234
rect 17192 8166 17250 8200
rect 14808 8074 14866 8132
rect 17192 8132 17204 8166
rect 17238 8132 17250 8166
rect 17192 8074 17250 8132
rect 14808 8062 17250 8074
rect 14808 8028 14924 8062
rect 14958 8028 14992 8062
rect 15026 8028 15060 8062
rect 15094 8028 15128 8062
rect 15162 8028 15196 8062
rect 15230 8028 15264 8062
rect 15298 8028 15332 8062
rect 15366 8028 15400 8062
rect 15434 8028 15468 8062
rect 15502 8028 15536 8062
rect 15570 8028 15604 8062
rect 15638 8028 15672 8062
rect 15706 8028 15740 8062
rect 15774 8028 15808 8062
rect 15842 8028 15876 8062
rect 15910 8028 15944 8062
rect 15978 8028 16012 8062
rect 16046 8028 16080 8062
rect 16114 8028 16148 8062
rect 16182 8028 16216 8062
rect 16250 8028 16284 8062
rect 16318 8028 16352 8062
rect 16386 8028 16420 8062
rect 16454 8028 16488 8062
rect 16522 8028 16556 8062
rect 16590 8028 16624 8062
rect 16658 8028 16692 8062
rect 16726 8028 16760 8062
rect 16794 8028 16828 8062
rect 16862 8028 16896 8062
rect 16930 8028 16964 8062
rect 16998 8028 17032 8062
rect 17066 8028 17100 8062
rect 17134 8028 17250 8062
rect 14808 8016 17250 8028
rect 17332 11440 19774 11452
rect 17332 11406 17448 11440
rect 17482 11406 17516 11440
rect 17550 11406 17584 11440
rect 17618 11406 17652 11440
rect 17686 11406 17720 11440
rect 17754 11406 17788 11440
rect 17822 11406 17856 11440
rect 17890 11406 17924 11440
rect 17958 11406 17992 11440
rect 18026 11406 18060 11440
rect 18094 11406 18128 11440
rect 18162 11406 18196 11440
rect 18230 11406 18264 11440
rect 18298 11406 18332 11440
rect 18366 11406 18400 11440
rect 18434 11406 18468 11440
rect 18502 11406 18536 11440
rect 18570 11406 18604 11440
rect 18638 11406 18672 11440
rect 18706 11406 18740 11440
rect 18774 11406 18808 11440
rect 18842 11406 18876 11440
rect 18910 11406 18944 11440
rect 18978 11406 19012 11440
rect 19046 11406 19080 11440
rect 19114 11406 19148 11440
rect 19182 11406 19216 11440
rect 19250 11406 19284 11440
rect 19318 11406 19352 11440
rect 19386 11406 19420 11440
rect 19454 11406 19488 11440
rect 19522 11406 19556 11440
rect 19590 11406 19624 11440
rect 19658 11406 19774 11440
rect 17332 11394 19774 11406
rect 17332 11336 17390 11394
rect 17332 11302 17344 11336
rect 17378 11302 17390 11336
rect 19716 11336 19774 11394
rect 17332 11268 17390 11302
rect 17332 11234 17344 11268
rect 17378 11234 17390 11268
rect 17332 11200 17390 11234
rect 19716 11302 19728 11336
rect 19762 11302 19774 11336
rect 19716 11268 19774 11302
rect 19716 11234 19728 11268
rect 19762 11234 19774 11268
rect 17332 11166 17344 11200
rect 17378 11166 17390 11200
rect 17332 11132 17390 11166
rect 17332 11098 17344 11132
rect 17378 11098 17390 11132
rect 17332 11064 17390 11098
rect 17332 11030 17344 11064
rect 17378 11030 17390 11064
rect 17332 10996 17390 11030
rect 17332 10962 17344 10996
rect 17378 10962 17390 10996
rect 17332 10928 17390 10962
rect 17332 10894 17344 10928
rect 17378 10894 17390 10928
rect 17332 10860 17390 10894
rect 17332 10826 17344 10860
rect 17378 10826 17390 10860
rect 17332 10792 17390 10826
rect 17332 10758 17344 10792
rect 17378 10758 17390 10792
rect 17332 10724 17390 10758
rect 17332 10690 17344 10724
rect 17378 10690 17390 10724
rect 17332 10656 17390 10690
rect 17332 10622 17344 10656
rect 17378 10622 17390 10656
rect 17332 10588 17390 10622
rect 17332 10554 17344 10588
rect 17378 10554 17390 10588
rect 17332 10520 17390 10554
rect 17332 10486 17344 10520
rect 17378 10486 17390 10520
rect 17332 10452 17390 10486
rect 17332 10418 17344 10452
rect 17378 10418 17390 10452
rect 17332 10384 17390 10418
rect 17332 10350 17344 10384
rect 17378 10350 17390 10384
rect 17332 10316 17390 10350
rect 17332 10282 17344 10316
rect 17378 10282 17390 10316
rect 17332 10248 17390 10282
rect 17332 10214 17344 10248
rect 17378 10214 17390 10248
rect 17332 10180 17390 10214
rect 17332 10146 17344 10180
rect 17378 10146 17390 10180
rect 17332 10112 17390 10146
rect 17332 10078 17344 10112
rect 17378 10078 17390 10112
rect 17332 10044 17390 10078
rect 17332 10010 17344 10044
rect 17378 10010 17390 10044
rect 17332 9976 17390 10010
rect 17332 9942 17344 9976
rect 17378 9942 17390 9976
rect 17332 9908 17390 9942
rect 17332 9874 17344 9908
rect 17378 9874 17390 9908
rect 17332 9840 17390 9874
rect 17332 9806 17344 9840
rect 17378 9806 17390 9840
rect 17332 9772 17390 9806
rect 17332 9738 17344 9772
rect 17378 9738 17390 9772
rect 17332 9704 17390 9738
rect 17332 9670 17344 9704
rect 17378 9670 17390 9704
rect 17332 9636 17390 9670
rect 17332 9602 17344 9636
rect 17378 9602 17390 9636
rect 17332 9568 17390 9602
rect 17332 9534 17344 9568
rect 17378 9534 17390 9568
rect 17332 9500 17390 9534
rect 17332 9466 17344 9500
rect 17378 9466 17390 9500
rect 17332 9432 17390 9466
rect 17332 9398 17344 9432
rect 17378 9398 17390 9432
rect 17332 9364 17390 9398
rect 17332 9330 17344 9364
rect 17378 9330 17390 9364
rect 17332 9296 17390 9330
rect 17332 9262 17344 9296
rect 17378 9262 17390 9296
rect 17332 9228 17390 9262
rect 17332 9194 17344 9228
rect 17378 9194 17390 9228
rect 17332 9160 17390 9194
rect 17332 9126 17344 9160
rect 17378 9126 17390 9160
rect 17332 9092 17390 9126
rect 17332 9058 17344 9092
rect 17378 9058 17390 9092
rect 17332 9024 17390 9058
rect 17332 8990 17344 9024
rect 17378 8990 17390 9024
rect 17332 8956 17390 8990
rect 17332 8922 17344 8956
rect 17378 8922 17390 8956
rect 17332 8888 17390 8922
rect 17332 8854 17344 8888
rect 17378 8854 17390 8888
rect 17332 8820 17390 8854
rect 17332 8786 17344 8820
rect 17378 8786 17390 8820
rect 17332 8752 17390 8786
rect 17332 8718 17344 8752
rect 17378 8718 17390 8752
rect 17332 8684 17390 8718
rect 17332 8650 17344 8684
rect 17378 8650 17390 8684
rect 17332 8616 17390 8650
rect 17332 8582 17344 8616
rect 17378 8582 17390 8616
rect 17332 8548 17390 8582
rect 17332 8514 17344 8548
rect 17378 8514 17390 8548
rect 17332 8480 17390 8514
rect 17332 8446 17344 8480
rect 17378 8446 17390 8480
rect 17332 8412 17390 8446
rect 17332 8378 17344 8412
rect 17378 8378 17390 8412
rect 17332 8344 17390 8378
rect 17332 8310 17344 8344
rect 17378 8310 17390 8344
rect 17332 8276 17390 8310
rect 17332 8242 17344 8276
rect 17378 8242 17390 8276
rect 17332 8208 17390 8242
rect 19716 11200 19774 11234
rect 19716 11166 19728 11200
rect 19762 11166 19774 11200
rect 19716 11132 19774 11166
rect 19716 11098 19728 11132
rect 19762 11098 19774 11132
rect 19716 11064 19774 11098
rect 19716 11030 19728 11064
rect 19762 11030 19774 11064
rect 19716 10996 19774 11030
rect 19716 10962 19728 10996
rect 19762 10962 19774 10996
rect 19716 10928 19774 10962
rect 19716 10894 19728 10928
rect 19762 10894 19774 10928
rect 19716 10860 19774 10894
rect 19716 10826 19728 10860
rect 19762 10826 19774 10860
rect 19716 10792 19774 10826
rect 19716 10758 19728 10792
rect 19762 10758 19774 10792
rect 19716 10724 19774 10758
rect 19716 10690 19728 10724
rect 19762 10690 19774 10724
rect 19716 10656 19774 10690
rect 19716 10622 19728 10656
rect 19762 10622 19774 10656
rect 19716 10588 19774 10622
rect 19716 10554 19728 10588
rect 19762 10554 19774 10588
rect 19716 10520 19774 10554
rect 19716 10486 19728 10520
rect 19762 10486 19774 10520
rect 19716 10452 19774 10486
rect 19716 10418 19728 10452
rect 19762 10418 19774 10452
rect 19716 10384 19774 10418
rect 19716 10350 19728 10384
rect 19762 10350 19774 10384
rect 19716 10316 19774 10350
rect 19716 10282 19728 10316
rect 19762 10282 19774 10316
rect 19716 10248 19774 10282
rect 19716 10214 19728 10248
rect 19762 10214 19774 10248
rect 19716 10180 19774 10214
rect 19716 10146 19728 10180
rect 19762 10146 19774 10180
rect 19716 10112 19774 10146
rect 19716 10078 19728 10112
rect 19762 10078 19774 10112
rect 19716 10044 19774 10078
rect 19716 10010 19728 10044
rect 19762 10010 19774 10044
rect 19716 9976 19774 10010
rect 19716 9942 19728 9976
rect 19762 9942 19774 9976
rect 19716 9908 19774 9942
rect 19716 9874 19728 9908
rect 19762 9874 19774 9908
rect 19716 9840 19774 9874
rect 19716 9806 19728 9840
rect 19762 9806 19774 9840
rect 19716 9772 19774 9806
rect 19716 9738 19728 9772
rect 19762 9738 19774 9772
rect 19716 9704 19774 9738
rect 19716 9670 19728 9704
rect 19762 9670 19774 9704
rect 19716 9636 19774 9670
rect 19716 9602 19728 9636
rect 19762 9602 19774 9636
rect 19716 9568 19774 9602
rect 19716 9534 19728 9568
rect 19762 9534 19774 9568
rect 19716 9500 19774 9534
rect 19716 9466 19728 9500
rect 19762 9466 19774 9500
rect 19716 9432 19774 9466
rect 19716 9398 19728 9432
rect 19762 9398 19774 9432
rect 19716 9364 19774 9398
rect 19716 9330 19728 9364
rect 19762 9330 19774 9364
rect 19716 9296 19774 9330
rect 19716 9262 19728 9296
rect 19762 9262 19774 9296
rect 19716 9228 19774 9262
rect 19716 9194 19728 9228
rect 19762 9194 19774 9228
rect 19716 9160 19774 9194
rect 19716 9126 19728 9160
rect 19762 9126 19774 9160
rect 19716 9092 19774 9126
rect 19716 9058 19728 9092
rect 19762 9058 19774 9092
rect 19716 9024 19774 9058
rect 19716 8990 19728 9024
rect 19762 8990 19774 9024
rect 19716 8956 19774 8990
rect 19716 8922 19728 8956
rect 19762 8922 19774 8956
rect 19716 8888 19774 8922
rect 19716 8854 19728 8888
rect 19762 8854 19774 8888
rect 19716 8820 19774 8854
rect 19716 8786 19728 8820
rect 19762 8786 19774 8820
rect 19716 8752 19774 8786
rect 19716 8718 19728 8752
rect 19762 8718 19774 8752
rect 19716 8684 19774 8718
rect 19716 8650 19728 8684
rect 19762 8650 19774 8684
rect 19716 8616 19774 8650
rect 19716 8582 19728 8616
rect 19762 8582 19774 8616
rect 19716 8548 19774 8582
rect 19716 8514 19728 8548
rect 19762 8514 19774 8548
rect 19716 8480 19774 8514
rect 19716 8446 19728 8480
rect 19762 8446 19774 8480
rect 19716 8412 19774 8446
rect 19716 8378 19728 8412
rect 19762 8378 19774 8412
rect 19716 8344 19774 8378
rect 19716 8310 19728 8344
rect 19762 8310 19774 8344
rect 19716 8276 19774 8310
rect 19716 8242 19728 8276
rect 19762 8242 19774 8276
rect 17332 8174 17344 8208
rect 17378 8174 17390 8208
rect 17332 8140 17390 8174
rect 17332 8106 17344 8140
rect 17378 8106 17390 8140
rect 19716 8208 19774 8242
rect 19716 8174 19728 8208
rect 19762 8174 19774 8208
rect 19716 8140 19774 8174
rect 17332 8048 17390 8106
rect 19716 8106 19728 8140
rect 19762 8106 19774 8140
rect 19716 8048 19774 8106
rect 17332 8036 19774 8048
rect 17332 8002 17448 8036
rect 17482 8002 17516 8036
rect 17550 8002 17584 8036
rect 17618 8002 17652 8036
rect 17686 8002 17720 8036
rect 17754 8002 17788 8036
rect 17822 8002 17856 8036
rect 17890 8002 17924 8036
rect 17958 8002 17992 8036
rect 18026 8002 18060 8036
rect 18094 8002 18128 8036
rect 18162 8002 18196 8036
rect 18230 8002 18264 8036
rect 18298 8002 18332 8036
rect 18366 8002 18400 8036
rect 18434 8002 18468 8036
rect 18502 8002 18536 8036
rect 18570 8002 18604 8036
rect 18638 8002 18672 8036
rect 18706 8002 18740 8036
rect 18774 8002 18808 8036
rect 18842 8002 18876 8036
rect 18910 8002 18944 8036
rect 18978 8002 19012 8036
rect 19046 8002 19080 8036
rect 19114 8002 19148 8036
rect 19182 8002 19216 8036
rect 19250 8002 19284 8036
rect 19318 8002 19352 8036
rect 19386 8002 19420 8036
rect 19454 8002 19488 8036
rect 19522 8002 19556 8036
rect 19590 8002 19624 8036
rect 19658 8002 19774 8036
rect 17332 7990 19774 8002
rect 22978 13490 24440 13502
rect 22978 13456 23114 13490
rect 23148 13456 23182 13490
rect 23216 13456 23250 13490
rect 23284 13456 23318 13490
rect 23352 13456 23386 13490
rect 23420 13456 23454 13490
rect 23488 13456 23522 13490
rect 23556 13456 23590 13490
rect 23624 13456 23658 13490
rect 23692 13456 23726 13490
rect 23760 13456 23794 13490
rect 23828 13456 23862 13490
rect 23896 13456 23930 13490
rect 23964 13456 23998 13490
rect 24032 13456 24066 13490
rect 24100 13456 24134 13490
rect 24168 13456 24202 13490
rect 24236 13456 24270 13490
rect 24304 13456 24440 13490
rect 22978 13444 24440 13456
rect 22978 13371 23036 13444
rect 22978 13337 22990 13371
rect 23024 13337 23036 13371
rect 24382 13371 24440 13444
rect 22978 13303 23036 13337
rect 24382 13337 24394 13371
rect 24428 13337 24440 13371
rect 22978 13269 22990 13303
rect 23024 13269 23036 13303
rect 22978 13235 23036 13269
rect 22978 13201 22990 13235
rect 23024 13201 23036 13235
rect 22978 13167 23036 13201
rect 22978 13133 22990 13167
rect 23024 13133 23036 13167
rect 22978 13099 23036 13133
rect 22978 13065 22990 13099
rect 23024 13065 23036 13099
rect 22978 13031 23036 13065
rect 22978 12997 22990 13031
rect 23024 12997 23036 13031
rect 22978 12963 23036 12997
rect 22978 12929 22990 12963
rect 23024 12929 23036 12963
rect 22978 12895 23036 12929
rect 22978 12861 22990 12895
rect 23024 12861 23036 12895
rect 22978 12827 23036 12861
rect 22978 12793 22990 12827
rect 23024 12793 23036 12827
rect 22978 12759 23036 12793
rect 22978 12725 22990 12759
rect 23024 12725 23036 12759
rect 22978 12691 23036 12725
rect 22978 12657 22990 12691
rect 23024 12657 23036 12691
rect 22978 12623 23036 12657
rect 22978 12589 22990 12623
rect 23024 12589 23036 12623
rect 22978 12555 23036 12589
rect 22978 12521 22990 12555
rect 23024 12521 23036 12555
rect 22978 12487 23036 12521
rect 22978 12453 22990 12487
rect 23024 12453 23036 12487
rect 22978 12419 23036 12453
rect 22978 12385 22990 12419
rect 23024 12385 23036 12419
rect 22978 12351 23036 12385
rect 22978 12317 22990 12351
rect 23024 12317 23036 12351
rect 22978 12283 23036 12317
rect 24382 13303 24440 13337
rect 24382 13269 24394 13303
rect 24428 13269 24440 13303
rect 24382 13235 24440 13269
rect 24382 13201 24394 13235
rect 24428 13201 24440 13235
rect 24382 13167 24440 13201
rect 24382 13133 24394 13167
rect 24428 13133 24440 13167
rect 24382 13099 24440 13133
rect 24382 13065 24394 13099
rect 24428 13065 24440 13099
rect 24382 13031 24440 13065
rect 24382 12997 24394 13031
rect 24428 12997 24440 13031
rect 24382 12963 24440 12997
rect 24382 12929 24394 12963
rect 24428 12929 24440 12963
rect 24382 12895 24440 12929
rect 24382 12861 24394 12895
rect 24428 12861 24440 12895
rect 24382 12827 24440 12861
rect 24382 12793 24394 12827
rect 24428 12793 24440 12827
rect 24382 12759 24440 12793
rect 24382 12725 24394 12759
rect 24428 12725 24440 12759
rect 24382 12691 24440 12725
rect 24382 12657 24394 12691
rect 24428 12657 24440 12691
rect 24382 12623 24440 12657
rect 24382 12589 24394 12623
rect 24428 12589 24440 12623
rect 24382 12555 24440 12589
rect 24382 12521 24394 12555
rect 24428 12521 24440 12555
rect 24382 12487 24440 12521
rect 24382 12453 24394 12487
rect 24428 12453 24440 12487
rect 24382 12419 24440 12453
rect 24382 12385 24394 12419
rect 24428 12385 24440 12419
rect 24382 12351 24440 12385
rect 24382 12317 24394 12351
rect 24428 12317 24440 12351
rect 22978 12249 22990 12283
rect 23024 12249 23036 12283
rect 24382 12283 24440 12317
rect 22978 12176 23036 12249
rect 24382 12249 24394 12283
rect 24428 12249 24440 12283
rect 24382 12176 24440 12249
rect 22978 12164 24440 12176
rect 22978 12130 23114 12164
rect 23148 12130 23182 12164
rect 23216 12130 23250 12164
rect 23284 12130 23318 12164
rect 23352 12130 23386 12164
rect 23420 12130 23454 12164
rect 23488 12130 23522 12164
rect 23556 12130 23590 12164
rect 23624 12130 23658 12164
rect 23692 12130 23726 12164
rect 23760 12130 23794 12164
rect 23828 12130 23862 12164
rect 23896 12130 23930 12164
rect 23964 12130 23998 12164
rect 24032 12130 24066 12164
rect 24100 12130 24134 12164
rect 24168 12130 24202 12164
rect 24236 12130 24270 12164
rect 24304 12130 24440 12164
rect 22978 12118 24440 12130
rect 24538 13484 26000 13496
rect 24538 13450 24674 13484
rect 24708 13450 24742 13484
rect 24776 13450 24810 13484
rect 24844 13450 24878 13484
rect 24912 13450 24946 13484
rect 24980 13450 25014 13484
rect 25048 13450 25082 13484
rect 25116 13450 25150 13484
rect 25184 13450 25218 13484
rect 25252 13450 25286 13484
rect 25320 13450 25354 13484
rect 25388 13450 25422 13484
rect 25456 13450 25490 13484
rect 25524 13450 25558 13484
rect 25592 13450 25626 13484
rect 25660 13450 25694 13484
rect 25728 13450 25762 13484
rect 25796 13450 25830 13484
rect 25864 13450 26000 13484
rect 24538 13438 26000 13450
rect 24538 13376 24596 13438
rect 24538 13342 24550 13376
rect 24584 13342 24596 13376
rect 25942 13376 26000 13438
rect 24538 13308 24596 13342
rect 24538 13274 24550 13308
rect 24584 13274 24596 13308
rect 25942 13342 25954 13376
rect 25988 13342 26000 13376
rect 25942 13308 26000 13342
rect 24538 13240 24596 13274
rect 24538 13206 24550 13240
rect 24584 13206 24596 13240
rect 24538 13172 24596 13206
rect 24538 13138 24550 13172
rect 24584 13138 24596 13172
rect 24538 13104 24596 13138
rect 24538 13070 24550 13104
rect 24584 13070 24596 13104
rect 24538 13036 24596 13070
rect 24538 13002 24550 13036
rect 24584 13002 24596 13036
rect 24538 12968 24596 13002
rect 24538 12934 24550 12968
rect 24584 12934 24596 12968
rect 24538 12900 24596 12934
rect 24538 12866 24550 12900
rect 24584 12866 24596 12900
rect 24538 12832 24596 12866
rect 24538 12798 24550 12832
rect 24584 12798 24596 12832
rect 24538 12764 24596 12798
rect 24538 12730 24550 12764
rect 24584 12730 24596 12764
rect 24538 12696 24596 12730
rect 24538 12662 24550 12696
rect 24584 12662 24596 12696
rect 24538 12628 24596 12662
rect 24538 12594 24550 12628
rect 24584 12594 24596 12628
rect 24538 12560 24596 12594
rect 24538 12526 24550 12560
rect 24584 12526 24596 12560
rect 24538 12492 24596 12526
rect 24538 12458 24550 12492
rect 24584 12458 24596 12492
rect 24538 12424 24596 12458
rect 24538 12390 24550 12424
rect 24584 12390 24596 12424
rect 24538 12356 24596 12390
rect 24538 12322 24550 12356
rect 24584 12322 24596 12356
rect 24538 12288 24596 12322
rect 25942 13274 25954 13308
rect 25988 13274 26000 13308
rect 25942 13240 26000 13274
rect 25942 13206 25954 13240
rect 25988 13206 26000 13240
rect 25942 13172 26000 13206
rect 25942 13138 25954 13172
rect 25988 13138 26000 13172
rect 25942 13104 26000 13138
rect 25942 13070 25954 13104
rect 25988 13070 26000 13104
rect 25942 13036 26000 13070
rect 25942 13002 25954 13036
rect 25988 13002 26000 13036
rect 25942 12968 26000 13002
rect 25942 12934 25954 12968
rect 25988 12934 26000 12968
rect 25942 12900 26000 12934
rect 25942 12866 25954 12900
rect 25988 12866 26000 12900
rect 25942 12832 26000 12866
rect 25942 12798 25954 12832
rect 25988 12798 26000 12832
rect 25942 12764 26000 12798
rect 25942 12730 25954 12764
rect 25988 12730 26000 12764
rect 25942 12696 26000 12730
rect 25942 12662 25954 12696
rect 25988 12662 26000 12696
rect 25942 12628 26000 12662
rect 25942 12594 25954 12628
rect 25988 12594 26000 12628
rect 25942 12560 26000 12594
rect 25942 12526 25954 12560
rect 25988 12526 26000 12560
rect 25942 12492 26000 12526
rect 25942 12458 25954 12492
rect 25988 12458 26000 12492
rect 25942 12424 26000 12458
rect 25942 12390 25954 12424
rect 25988 12390 26000 12424
rect 25942 12356 26000 12390
rect 25942 12322 25954 12356
rect 25988 12322 26000 12356
rect 24538 12254 24550 12288
rect 24584 12254 24596 12288
rect 24538 12220 24596 12254
rect 25942 12288 26000 12322
rect 25942 12254 25954 12288
rect 25988 12254 26000 12288
rect 24538 12186 24550 12220
rect 24584 12186 24596 12220
rect 24538 12152 24596 12186
rect 24538 12118 24550 12152
rect 24584 12118 24596 12152
rect 24538 12084 24596 12118
rect 24538 12050 24550 12084
rect 24584 12050 24596 12084
rect 24538 12016 24596 12050
rect 24538 11982 24550 12016
rect 24584 11982 24596 12016
rect 24538 11948 24596 11982
rect 24538 11914 24550 11948
rect 24584 11914 24596 11948
rect 24538 11880 24596 11914
rect 24538 11846 24550 11880
rect 24584 11846 24596 11880
rect 24538 11812 24596 11846
rect 24538 11778 24550 11812
rect 24584 11778 24596 11812
rect 24538 11744 24596 11778
rect 24538 11710 24550 11744
rect 24584 11710 24596 11744
rect 24538 11676 24596 11710
rect 24538 11642 24550 11676
rect 24584 11642 24596 11676
rect 24538 11608 24596 11642
rect 24538 11574 24550 11608
rect 24584 11574 24596 11608
rect 24538 11540 24596 11574
rect 24538 11506 24550 11540
rect 24584 11506 24596 11540
rect 24538 11472 24596 11506
rect 24538 11438 24550 11472
rect 24584 11438 24596 11472
rect 24538 11404 24596 11438
rect 24538 11370 24550 11404
rect 24584 11370 24596 11404
rect 24538 11336 24596 11370
rect 24538 11302 24550 11336
rect 24584 11302 24596 11336
rect 24538 11268 24596 11302
rect 24538 11234 24550 11268
rect 24584 11234 24596 11268
rect 25942 12220 26000 12254
rect 25942 12186 25954 12220
rect 25988 12186 26000 12220
rect 25942 12152 26000 12186
rect 25942 12118 25954 12152
rect 25988 12118 26000 12152
rect 25942 12084 26000 12118
rect 25942 12050 25954 12084
rect 25988 12050 26000 12084
rect 25942 12016 26000 12050
rect 25942 11982 25954 12016
rect 25988 11982 26000 12016
rect 25942 11948 26000 11982
rect 25942 11914 25954 11948
rect 25988 11914 26000 11948
rect 25942 11880 26000 11914
rect 25942 11846 25954 11880
rect 25988 11846 26000 11880
rect 25942 11812 26000 11846
rect 25942 11778 25954 11812
rect 25988 11778 26000 11812
rect 25942 11744 26000 11778
rect 25942 11710 25954 11744
rect 25988 11710 26000 11744
rect 25942 11676 26000 11710
rect 25942 11642 25954 11676
rect 25988 11642 26000 11676
rect 25942 11608 26000 11642
rect 25942 11574 25954 11608
rect 25988 11574 26000 11608
rect 25942 11540 26000 11574
rect 25942 11506 25954 11540
rect 25988 11506 26000 11540
rect 25942 11472 26000 11506
rect 25942 11438 25954 11472
rect 25988 11438 26000 11472
rect 25942 11404 26000 11438
rect 25942 11370 25954 11404
rect 25988 11370 26000 11404
rect 25942 11336 26000 11370
rect 25942 11302 25954 11336
rect 25988 11302 26000 11336
rect 25942 11268 26000 11302
rect 24538 11200 24596 11234
rect 24538 11166 24550 11200
rect 24584 11166 24596 11200
rect 25942 11234 25954 11268
rect 25988 11234 26000 11268
rect 25942 11200 26000 11234
rect 24538 11132 24596 11166
rect 24538 11098 24550 11132
rect 24584 11098 24596 11132
rect 24538 11064 24596 11098
rect 24538 11030 24550 11064
rect 24584 11030 24596 11064
rect 24538 10996 24596 11030
rect 24538 10962 24550 10996
rect 24584 10962 24596 10996
rect 24538 10928 24596 10962
rect 24538 10894 24550 10928
rect 24584 10894 24596 10928
rect 24538 10860 24596 10894
rect 24538 10826 24550 10860
rect 24584 10826 24596 10860
rect 24538 10792 24596 10826
rect 24538 10758 24550 10792
rect 24584 10758 24596 10792
rect 24538 10724 24596 10758
rect 24538 10690 24550 10724
rect 24584 10690 24596 10724
rect 24538 10656 24596 10690
rect 24538 10622 24550 10656
rect 24584 10622 24596 10656
rect 24538 10588 24596 10622
rect 24538 10554 24550 10588
rect 24584 10554 24596 10588
rect 24538 10520 24596 10554
rect 24538 10486 24550 10520
rect 24584 10486 24596 10520
rect 24538 10452 24596 10486
rect 24538 10418 24550 10452
rect 24584 10418 24596 10452
rect 24538 10384 24596 10418
rect 24538 10350 24550 10384
rect 24584 10350 24596 10384
rect 24538 10316 24596 10350
rect 24538 10282 24550 10316
rect 24584 10282 24596 10316
rect 24538 10248 24596 10282
rect 24538 10214 24550 10248
rect 24584 10214 24596 10248
rect 24538 10180 24596 10214
rect 25942 11166 25954 11200
rect 25988 11166 26000 11200
rect 25942 11132 26000 11166
rect 25942 11098 25954 11132
rect 25988 11098 26000 11132
rect 25942 11064 26000 11098
rect 25942 11030 25954 11064
rect 25988 11030 26000 11064
rect 25942 10996 26000 11030
rect 25942 10962 25954 10996
rect 25988 10962 26000 10996
rect 25942 10928 26000 10962
rect 25942 10894 25954 10928
rect 25988 10894 26000 10928
rect 25942 10860 26000 10894
rect 25942 10826 25954 10860
rect 25988 10826 26000 10860
rect 25942 10792 26000 10826
rect 25942 10758 25954 10792
rect 25988 10758 26000 10792
rect 25942 10724 26000 10758
rect 25942 10690 25954 10724
rect 25988 10690 26000 10724
rect 25942 10656 26000 10690
rect 25942 10622 25954 10656
rect 25988 10622 26000 10656
rect 25942 10588 26000 10622
rect 25942 10554 25954 10588
rect 25988 10554 26000 10588
rect 25942 10520 26000 10554
rect 25942 10486 25954 10520
rect 25988 10486 26000 10520
rect 25942 10452 26000 10486
rect 25942 10418 25954 10452
rect 25988 10418 26000 10452
rect 25942 10384 26000 10418
rect 25942 10350 25954 10384
rect 25988 10350 26000 10384
rect 25942 10316 26000 10350
rect 25942 10282 25954 10316
rect 25988 10282 26000 10316
rect 25942 10248 26000 10282
rect 25942 10214 25954 10248
rect 25988 10214 26000 10248
rect 24538 10146 24550 10180
rect 24584 10146 24596 10180
rect 24538 10112 24596 10146
rect 25942 10180 26000 10214
rect 25942 10146 25954 10180
rect 25988 10146 26000 10180
rect 24538 10078 24550 10112
rect 24584 10078 24596 10112
rect 24538 10044 24596 10078
rect 24538 10010 24550 10044
rect 24584 10010 24596 10044
rect 24538 9976 24596 10010
rect 24538 9942 24550 9976
rect 24584 9942 24596 9976
rect 24538 9908 24596 9942
rect 24538 9874 24550 9908
rect 24584 9874 24596 9908
rect 24538 9840 24596 9874
rect 24538 9806 24550 9840
rect 24584 9806 24596 9840
rect 24538 9772 24596 9806
rect 24538 9738 24550 9772
rect 24584 9738 24596 9772
rect 24538 9704 24596 9738
rect 24538 9670 24550 9704
rect 24584 9670 24596 9704
rect 24538 9636 24596 9670
rect 24538 9602 24550 9636
rect 24584 9602 24596 9636
rect 24538 9568 24596 9602
rect 24538 9534 24550 9568
rect 24584 9534 24596 9568
rect 24538 9500 24596 9534
rect 24538 9466 24550 9500
rect 24584 9466 24596 9500
rect 24538 9432 24596 9466
rect 24538 9398 24550 9432
rect 24584 9398 24596 9432
rect 24538 9364 24596 9398
rect 24538 9330 24550 9364
rect 24584 9330 24596 9364
rect 24538 9296 24596 9330
rect 24538 9262 24550 9296
rect 24584 9262 24596 9296
rect 24538 9228 24596 9262
rect 24538 9194 24550 9228
rect 24584 9194 24596 9228
rect 24538 9160 24596 9194
rect 24538 9126 24550 9160
rect 24584 9126 24596 9160
rect 25942 10112 26000 10146
rect 25942 10078 25954 10112
rect 25988 10078 26000 10112
rect 25942 10044 26000 10078
rect 25942 10010 25954 10044
rect 25988 10010 26000 10044
rect 25942 9976 26000 10010
rect 25942 9942 25954 9976
rect 25988 9942 26000 9976
rect 25942 9908 26000 9942
rect 25942 9874 25954 9908
rect 25988 9874 26000 9908
rect 25942 9840 26000 9874
rect 25942 9806 25954 9840
rect 25988 9806 26000 9840
rect 25942 9772 26000 9806
rect 25942 9738 25954 9772
rect 25988 9738 26000 9772
rect 25942 9704 26000 9738
rect 25942 9670 25954 9704
rect 25988 9670 26000 9704
rect 25942 9636 26000 9670
rect 25942 9602 25954 9636
rect 25988 9602 26000 9636
rect 25942 9568 26000 9602
rect 25942 9534 25954 9568
rect 25988 9534 26000 9568
rect 25942 9500 26000 9534
rect 25942 9466 25954 9500
rect 25988 9466 26000 9500
rect 25942 9432 26000 9466
rect 25942 9398 25954 9432
rect 25988 9398 26000 9432
rect 25942 9364 26000 9398
rect 25942 9330 25954 9364
rect 25988 9330 26000 9364
rect 25942 9296 26000 9330
rect 25942 9262 25954 9296
rect 25988 9262 26000 9296
rect 25942 9228 26000 9262
rect 25942 9194 25954 9228
rect 25988 9194 26000 9228
rect 25942 9160 26000 9194
rect 24538 9092 24596 9126
rect 24538 9058 24550 9092
rect 24584 9058 24596 9092
rect 25942 9126 25954 9160
rect 25988 9126 26000 9160
rect 25942 9092 26000 9126
rect 24538 8996 24596 9058
rect 25942 9058 25954 9092
rect 25988 9058 26000 9092
rect 25942 8996 26000 9058
rect 24538 8984 26000 8996
rect 24538 8950 24674 8984
rect 24708 8950 24742 8984
rect 24776 8950 24810 8984
rect 24844 8950 24878 8984
rect 24912 8950 24946 8984
rect 24980 8950 25014 8984
rect 25048 8950 25082 8984
rect 25116 8950 25150 8984
rect 25184 8950 25218 8984
rect 25252 8950 25286 8984
rect 25320 8950 25354 8984
rect 25388 8950 25422 8984
rect 25456 8950 25490 8984
rect 25524 8950 25558 8984
rect 25592 8950 25626 8984
rect 25660 8950 25694 8984
rect 25728 8950 25762 8984
rect 25796 8950 25830 8984
rect 25864 8950 26000 8984
rect 24538 8938 26000 8950
<< psubdiffcont >>
rect 24559 16716 24593 16750
rect 24627 16716 24661 16750
rect 24695 16716 24729 16750
rect 24763 16716 24797 16750
rect 24831 16716 24865 16750
rect 24899 16716 24933 16750
rect 24967 16716 25001 16750
rect 25035 16716 25069 16750
rect 25103 16716 25137 16750
rect 25171 16716 25205 16750
rect 25239 16716 25273 16750
rect 25307 16716 25341 16750
rect 25375 16716 25409 16750
rect 25443 16716 25477 16750
rect 25511 16716 25545 16750
rect 25579 16716 25613 16750
rect 25647 16716 25681 16750
rect 25715 16716 25749 16750
rect 25783 16716 25817 16750
rect 25851 16716 25885 16750
rect 25919 16716 25953 16750
rect 25987 16716 26021 16750
rect 26055 16716 26089 16750
rect 26123 16716 26157 16750
rect 26191 16716 26225 16750
rect 26259 16716 26293 16750
rect 26327 16716 26361 16750
rect 26395 16716 26429 16750
rect 26463 16716 26497 16750
rect 26531 16716 26565 16750
rect 26599 16716 26633 16750
rect 26667 16716 26701 16750
rect 26735 16716 26769 16750
rect 26803 16716 26837 16750
rect 26871 16716 26905 16750
rect 26939 16716 26973 16750
rect 27007 16716 27041 16750
rect 27075 16716 27109 16750
rect 27143 16716 27177 16750
rect 27211 16716 27245 16750
rect 27279 16716 27313 16750
rect 27347 16716 27381 16750
rect 27415 16716 27449 16750
rect 27483 16716 27517 16750
rect 27551 16716 27585 16750
rect 24460 16612 24494 16646
rect 24460 16544 24494 16578
rect 27650 16612 27684 16646
rect 24460 16476 24494 16510
rect 24460 16408 24494 16442
rect 24460 16340 24494 16374
rect 24460 16272 24494 16306
rect 27650 16544 27684 16578
rect 27650 16476 27684 16510
rect 27650 16408 27684 16442
rect 27650 16340 27684 16374
rect 24460 16204 24494 16238
rect 27650 16272 27684 16306
rect 24460 16136 24494 16170
rect 24460 16068 24494 16102
rect 24460 16000 24494 16034
rect 27650 16204 27684 16238
rect 27650 16136 27684 16170
rect 27650 16068 27684 16102
rect 27650 16000 27684 16034
rect 24460 15932 24494 15966
rect 27650 15932 27684 15966
rect 24460 15864 24494 15898
rect 23144 15760 23178 15794
rect 23240 15783 23274 15817
rect 23330 15783 23364 15817
rect 23420 15783 23454 15817
rect 23510 15783 23544 15817
rect 23600 15783 23634 15817
rect 23690 15783 23724 15817
rect 23780 15783 23814 15817
rect 23870 15783 23904 15817
rect 23960 15783 23994 15817
rect 24050 15783 24084 15817
rect 24140 15783 24174 15817
rect 24230 15783 24264 15817
rect 24331 15760 24365 15794
rect 23144 15670 23178 15704
rect 23144 15580 23178 15614
rect -7630 15432 -7596 15466
rect -7562 15432 -7528 15466
rect -7494 15432 -7460 15466
rect -7426 15432 -7392 15466
rect -7358 15432 -7324 15466
rect -7290 15432 -7256 15466
rect -7222 15432 -7188 15466
rect -7154 15432 -7120 15466
rect -7086 15432 -7052 15466
rect -7018 15432 -6984 15466
rect -6950 15432 -6916 15466
rect -6882 15432 -6848 15466
rect -6814 15432 -6780 15466
rect -6746 15432 -6712 15466
rect -6678 15432 -6644 15466
rect -6610 15432 -6576 15466
rect -6542 15432 -6508 15466
rect -6474 15432 -6440 15466
rect -6406 15432 -6372 15466
rect -6338 15432 -6304 15466
rect -6270 15432 -6236 15466
rect -6202 15432 -6168 15466
rect -6134 15432 -6100 15466
rect -6066 15432 -6032 15466
rect -5998 15432 -5964 15466
rect -5930 15432 -5896 15466
rect -5862 15432 -5828 15466
rect -5794 15432 -5760 15466
rect -5726 15432 -5692 15466
rect -5658 15432 -5624 15466
rect -5590 15432 -5556 15466
rect -5522 15432 -5488 15466
rect -5454 15432 -5420 15466
rect -5386 15432 -5352 15466
rect -5318 15432 -5284 15466
rect -5250 15432 -5216 15466
rect -5182 15432 -5148 15466
rect -5114 15432 -5080 15466
rect -5046 15432 -5012 15466
rect -4978 15432 -4944 15466
rect -4910 15432 -4876 15466
rect -4842 15432 -4808 15466
rect -4774 15432 -4740 15466
rect -4706 15432 -4672 15466
rect -7843 15274 -7809 15308
rect -7843 15206 -7809 15240
rect -7843 15138 -7809 15172
rect -7843 15070 -7809 15104
rect -7843 15002 -7809 15036
rect -4503 15234 -4469 15268
rect -4503 15166 -4469 15200
rect -4503 15098 -4469 15132
rect -4503 15030 -4469 15064
rect 23144 15490 23178 15524
rect 23144 15400 23178 15434
rect 23144 15310 23178 15344
rect 23144 15220 23178 15254
rect 23144 15130 23178 15164
rect 23144 15040 23178 15074
rect -7843 14934 -7809 14968
rect -7843 14866 -7809 14900
rect -4503 14962 -4469 14996
rect -4503 14894 -4469 14928
rect -7843 14798 -7809 14832
rect -7843 14730 -7809 14764
rect -7843 14662 -7809 14696
rect -7843 14594 -7809 14628
rect -7843 14526 -7809 14560
rect -7843 14458 -7809 14492
rect -7843 14390 -7809 14424
rect -7843 14322 -7809 14356
rect -7843 14254 -7809 14288
rect -7843 14186 -7809 14220
rect -7843 14118 -7809 14152
rect -7843 14050 -7809 14084
rect -7843 13982 -7809 14016
rect -7843 13914 -7809 13948
rect -7843 13846 -7809 13880
rect -7843 13778 -7809 13812
rect -7843 13710 -7809 13744
rect -7843 13642 -7809 13676
rect -7843 13574 -7809 13608
rect -7843 13506 -7809 13540
rect -7843 13438 -7809 13472
rect -7843 13370 -7809 13404
rect -7843 13302 -7809 13336
rect -7843 13234 -7809 13268
rect -7843 13166 -7809 13200
rect -7843 13098 -7809 13132
rect -7843 13030 -7809 13064
rect -7843 12962 -7809 12996
rect -7843 12894 -7809 12928
rect -7843 12826 -7809 12860
rect -4503 14826 -4469 14860
rect -4503 14758 -4469 14792
rect -4503 14690 -4469 14724
rect -4503 14622 -4469 14656
rect -4503 14554 -4469 14588
rect -4503 14486 -4469 14520
rect -4503 14418 -4469 14452
rect -4503 14350 -4469 14384
rect -4503 14282 -4469 14316
rect -4503 14214 -4469 14248
rect -4503 14146 -4469 14180
rect -4503 14078 -4469 14112
rect -4503 14010 -4469 14044
rect -4503 13942 -4469 13976
rect -4503 13874 -4469 13908
rect -4503 13806 -4469 13840
rect -4503 13738 -4469 13772
rect -4503 13670 -4469 13704
rect -4503 13602 -4469 13636
rect -4503 13534 -4469 13568
rect -4503 13466 -4469 13500
rect -4503 13398 -4469 13432
rect -4503 13330 -4469 13364
rect -4503 13262 -4469 13296
rect -4503 13194 -4469 13228
rect -4503 13126 -4469 13160
rect -4503 13058 -4469 13092
rect -4503 12990 -4469 13024
rect -4503 12922 -4469 12956
rect -4503 12854 -4469 12888
rect -7843 12758 -7809 12792
rect -7843 12690 -7809 12724
rect -7843 12622 -7809 12656
rect -4503 12786 -4469 12820
rect -4503 12718 -4469 12752
rect -4503 12650 -4469 12684
rect -7843 12554 -7809 12588
rect -7843 12486 -7809 12520
rect -7843 12418 -7809 12452
rect -7843 12350 -7809 12384
rect -4503 12582 -4469 12616
rect -4503 12514 -4469 12548
rect -4503 12446 -4469 12480
rect -4503 12378 -4469 12412
rect -4503 12310 -4469 12344
rect -3896 15001 -3862 15035
rect -3828 15001 -3794 15035
rect -4010 14880 -3976 14914
rect -4010 14812 -3976 14846
rect -4010 14744 -3976 14778
rect -4010 14676 -3976 14710
rect -4010 14608 -3976 14642
rect -4010 14540 -3976 14574
rect -4010 14472 -3976 14506
rect -4010 14404 -3976 14438
rect -4010 14336 -3976 14370
rect -4010 14268 -3976 14302
rect -4010 14200 -3976 14234
rect -4010 14132 -3976 14166
rect -4010 14064 -3976 14098
rect -4010 13996 -3976 14030
rect -4010 13928 -3976 13962
rect -4010 13860 -3976 13894
rect -4010 13792 -3976 13826
rect -4010 13724 -3976 13758
rect -4010 13656 -3976 13690
rect -4010 13588 -3976 13622
rect -4010 13520 -3976 13554
rect -4010 13452 -3976 13486
rect -4010 13384 -3976 13418
rect -4010 13316 -3976 13350
rect -4010 13248 -3976 13282
rect -4010 13180 -3976 13214
rect -4010 13112 -3976 13146
rect -4010 13044 -3976 13078
rect -4010 12976 -3976 13010
rect -4010 12908 -3976 12942
rect -4010 12840 -3976 12874
rect -4010 12772 -3976 12806
rect -4010 12704 -3976 12738
rect -4010 12636 -3976 12670
rect -4010 12568 -3976 12602
rect -4010 12500 -3976 12534
rect -4010 12432 -3976 12466
rect -3714 14880 -3680 14914
rect -3714 14812 -3680 14846
rect -3714 14744 -3680 14778
rect -3714 14676 -3680 14710
rect -3714 14608 -3680 14642
rect -3714 14540 -3680 14574
rect -3714 14472 -3680 14506
rect -3714 14404 -3680 14438
rect -3714 14336 -3680 14370
rect -3714 14268 -3680 14302
rect -3714 14200 -3680 14234
rect -3714 14132 -3680 14166
rect -3714 14064 -3680 14098
rect -3714 13996 -3680 14030
rect -3714 13928 -3680 13962
rect -3714 13860 -3680 13894
rect -3714 13792 -3680 13826
rect -3714 13724 -3680 13758
rect -3714 13656 -3680 13690
rect -3714 13588 -3680 13622
rect -3714 13520 -3680 13554
rect -3714 13452 -3680 13486
rect -3714 13384 -3680 13418
rect -3714 13316 -3680 13350
rect -3714 13248 -3680 13282
rect -3714 13180 -3680 13214
rect -3714 13112 -3680 13146
rect -3714 13044 -3680 13078
rect -3714 12976 -3680 13010
rect -3714 12908 -3680 12942
rect -3714 12840 -3680 12874
rect -3714 12772 -3680 12806
rect -3714 12704 -3680 12738
rect -3714 12636 -3680 12670
rect -3714 12568 -3680 12602
rect -3714 12500 -3680 12534
rect -3714 12432 -3680 12466
rect -3896 12311 -3862 12345
rect -3828 12311 -3794 12345
rect -7570 12202 -7536 12236
rect -7502 12202 -7468 12236
rect -7434 12202 -7400 12236
rect -7366 12202 -7332 12236
rect -7298 12202 -7264 12236
rect -7230 12202 -7196 12236
rect -7162 12202 -7128 12236
rect -7094 12202 -7060 12236
rect -7026 12202 -6992 12236
rect -6958 12202 -6924 12236
rect -6890 12202 -6856 12236
rect -6822 12202 -6788 12236
rect -6754 12202 -6720 12236
rect -6686 12202 -6652 12236
rect -6618 12202 -6584 12236
rect -6550 12202 -6516 12236
rect -6482 12202 -6448 12236
rect -6414 12202 -6380 12236
rect -6346 12202 -6312 12236
rect -6278 12202 -6244 12236
rect -6210 12202 -6176 12236
rect -6142 12202 -6108 12236
rect -6074 12202 -6040 12236
rect -6006 12202 -5972 12236
rect -5938 12202 -5904 12236
rect -5870 12202 -5836 12236
rect -5802 12202 -5768 12236
rect -5734 12202 -5700 12236
rect -5666 12202 -5632 12236
rect -5598 12202 -5564 12236
rect -5530 12202 -5496 12236
rect -5462 12202 -5428 12236
rect -5394 12202 -5360 12236
rect -5326 12202 -5292 12236
rect -5258 12202 -5224 12236
rect -5190 12202 -5156 12236
rect -5122 12202 -5088 12236
rect -5054 12202 -5020 12236
rect -4986 12202 -4952 12236
rect -4918 12202 -4884 12236
rect -4850 12202 -4816 12236
rect -4782 12202 -4748 12236
rect -4714 12202 -4680 12236
rect -4646 12202 -4612 12236
rect 23144 14950 23178 14984
rect 23144 14860 23178 14894
rect 23144 14770 23178 14804
rect 24331 15670 24365 15704
rect 24331 15580 24365 15614
rect 24331 15490 24365 15524
rect 24331 15400 24365 15434
rect 24331 15310 24365 15344
rect 24331 15220 24365 15254
rect 24331 15130 24365 15164
rect 24460 15796 24494 15830
rect 24460 15728 24494 15762
rect 24460 15660 24494 15694
rect 27650 15864 27684 15898
rect 27650 15796 27684 15830
rect 27650 15728 27684 15762
rect 24460 15592 24494 15626
rect 27650 15660 27684 15694
rect 24460 15524 24494 15558
rect 24460 15456 24494 15490
rect 24460 15388 24494 15422
rect 24460 15320 24494 15354
rect 27650 15592 27684 15626
rect 27650 15524 27684 15558
rect 27650 15456 27684 15490
rect 27650 15388 27684 15422
rect 37962 16182 37996 16216
rect 38030 16182 38064 16216
rect 38098 16182 38132 16216
rect 38166 16182 38200 16216
rect 38234 16182 38268 16216
rect 38302 16182 38336 16216
rect 38370 16182 38404 16216
rect 38438 16182 38472 16216
rect 38506 16182 38540 16216
rect 38574 16182 38608 16216
rect 38642 16182 38676 16216
rect 38710 16182 38744 16216
rect 38778 16182 38812 16216
rect 38846 16182 38880 16216
rect 38914 16182 38948 16216
rect 38982 16182 39016 16216
rect 39050 16182 39084 16216
rect 39118 16182 39152 16216
rect 39186 16182 39220 16216
rect 39254 16182 39288 16216
rect 39322 16182 39356 16216
rect 39390 16182 39424 16216
rect 39458 16182 39492 16216
rect 39526 16182 39560 16216
rect 39594 16182 39628 16216
rect 39662 16182 39696 16216
rect 39730 16182 39764 16216
rect 39798 16182 39832 16216
rect 39866 16182 39900 16216
rect 39934 16182 39968 16216
rect 40002 16182 40036 16216
rect 40070 16182 40104 16216
rect 40138 16182 40172 16216
rect 40206 16182 40240 16216
rect 40274 16182 40308 16216
rect 40342 16182 40376 16216
rect 40410 16182 40444 16216
rect 40478 16182 40512 16216
rect 40546 16182 40580 16216
rect 40614 16182 40648 16216
rect 40682 16182 40716 16216
rect 40750 16182 40784 16216
rect 40818 16182 40852 16216
rect 40886 16182 40920 16216
rect 37749 16024 37783 16058
rect 37749 15956 37783 15990
rect 37749 15888 37783 15922
rect 37749 15820 37783 15854
rect 37749 15752 37783 15786
rect 41089 15984 41123 16018
rect 41089 15916 41123 15950
rect 41089 15848 41123 15882
rect 41089 15780 41123 15814
rect 37749 15684 37783 15718
rect 37749 15616 37783 15650
rect 41089 15712 41123 15746
rect 41089 15644 41123 15678
rect 37749 15548 37783 15582
rect 37749 15480 37783 15514
rect 37749 15412 37783 15446
rect 24460 15252 24494 15286
rect 27650 15320 27684 15354
rect 27650 15252 27684 15286
rect 24559 15148 24593 15182
rect 24627 15148 24661 15182
rect 24695 15148 24729 15182
rect 24763 15148 24797 15182
rect 24831 15148 24865 15182
rect 24899 15148 24933 15182
rect 24967 15148 25001 15182
rect 25035 15148 25069 15182
rect 25103 15148 25137 15182
rect 25171 15148 25205 15182
rect 25239 15148 25273 15182
rect 25307 15148 25341 15182
rect 25375 15148 25409 15182
rect 25443 15148 25477 15182
rect 25511 15148 25545 15182
rect 25579 15148 25613 15182
rect 25647 15148 25681 15182
rect 25715 15148 25749 15182
rect 25783 15148 25817 15182
rect 25851 15148 25885 15182
rect 25919 15148 25953 15182
rect 25987 15148 26021 15182
rect 26055 15148 26089 15182
rect 26123 15148 26157 15182
rect 26191 15148 26225 15182
rect 26259 15148 26293 15182
rect 26327 15148 26361 15182
rect 26395 15148 26429 15182
rect 26463 15148 26497 15182
rect 26531 15148 26565 15182
rect 26599 15148 26633 15182
rect 26667 15148 26701 15182
rect 26735 15148 26769 15182
rect 26803 15148 26837 15182
rect 26871 15148 26905 15182
rect 26939 15148 26973 15182
rect 27007 15148 27041 15182
rect 27075 15148 27109 15182
rect 27143 15148 27177 15182
rect 27211 15148 27245 15182
rect 27279 15148 27313 15182
rect 27347 15148 27381 15182
rect 27415 15148 27449 15182
rect 27483 15148 27517 15182
rect 27551 15148 27585 15182
rect 28960 15358 28994 15392
rect 29028 15358 29062 15392
rect 29096 15358 29130 15392
rect 29164 15358 29198 15392
rect 29232 15358 29266 15392
rect 29300 15358 29334 15392
rect 29368 15358 29402 15392
rect 29436 15358 29470 15392
rect 29504 15358 29538 15392
rect 29572 15358 29606 15392
rect 29640 15358 29674 15392
rect 28834 15241 28868 15275
rect 28834 15173 28868 15207
rect 24331 15040 24365 15074
rect 24331 14950 24365 14984
rect 24331 14860 24365 14894
rect 24331 14770 24365 14804
rect 23144 14680 23178 14714
rect 24331 14680 24365 14714
rect 20497 14566 20531 14600
rect 20565 14566 20599 14600
rect 20633 14566 20667 14600
rect 20701 14566 20735 14600
rect 20769 14566 20803 14600
rect 20837 14566 20871 14600
rect 20905 14566 20939 14600
rect 20973 14566 21007 14600
rect 21041 14566 21075 14600
rect 21109 14566 21143 14600
rect 21177 14566 21211 14600
rect 21245 14566 21279 14600
rect 21313 14566 21347 14600
rect 21381 14566 21415 14600
rect 21449 14566 21483 14600
rect 21517 14566 21551 14600
rect 20382 14440 20416 14474
rect 23240 14596 23274 14630
rect 23330 14596 23364 14630
rect 23420 14596 23454 14630
rect 23510 14596 23544 14630
rect 23600 14596 23634 14630
rect 23690 14596 23724 14630
rect 23780 14596 23814 14630
rect 23870 14596 23904 14630
rect 23960 14596 23994 14630
rect 24050 14596 24084 14630
rect 24140 14596 24174 14630
rect 24230 14596 24264 14630
rect 28834 15105 28868 15139
rect 28834 15037 28868 15071
rect 28834 14969 28868 15003
rect 28834 14901 28868 14935
rect 28834 14833 28868 14867
rect 28834 14765 28868 14799
rect 28834 14697 28868 14731
rect 28834 14629 28868 14663
rect 20382 14372 20416 14406
rect 20382 14304 20416 14338
rect 20382 14236 20416 14270
rect 20382 14168 20416 14202
rect 20382 14100 20416 14134
rect 20382 14032 20416 14066
rect 20382 13964 20416 13998
rect 20382 13896 20416 13930
rect 20382 13828 20416 13862
rect 20382 13760 20416 13794
rect 20382 13692 20416 13726
rect 20382 13624 20416 13658
rect 20382 13556 20416 13590
rect 20382 13488 20416 13522
rect 20382 13420 20416 13454
rect 20382 13352 20416 13386
rect 20382 13284 20416 13318
rect 20382 13216 20416 13250
rect 20382 13148 20416 13182
rect 20382 13080 20416 13114
rect 20382 13012 20416 13046
rect 20382 12944 20416 12978
rect 20382 12876 20416 12910
rect 20382 12808 20416 12842
rect 20382 12740 20416 12774
rect 20382 12672 20416 12706
rect 20382 12604 20416 12638
rect 20382 12536 20416 12570
rect 20382 12468 20416 12502
rect 20382 12400 20416 12434
rect 20382 12332 20416 12366
rect 20382 12264 20416 12298
rect 20382 12196 20416 12230
rect 20382 12128 20416 12162
rect 20382 12060 20416 12094
rect 20382 11992 20416 12026
rect 20382 11924 20416 11958
rect 20382 11856 20416 11890
rect 20382 11788 20416 11822
rect 20382 11720 20416 11754
rect 20382 11652 20416 11686
rect 20382 11584 20416 11618
rect 20382 11516 20416 11550
rect 12816 11242 12850 11276
rect 12912 11265 12946 11299
rect 13002 11265 13036 11299
rect 13092 11265 13126 11299
rect 13182 11265 13216 11299
rect 13272 11265 13306 11299
rect 13362 11265 13396 11299
rect 13452 11265 13486 11299
rect 13542 11265 13576 11299
rect 13632 11265 13666 11299
rect 13722 11265 13756 11299
rect 13812 11265 13846 11299
rect 13902 11265 13936 11299
rect 14003 11242 14037 11276
rect 12816 11152 12850 11186
rect 12816 11062 12850 11096
rect 12816 10972 12850 11006
rect 12816 10882 12850 10916
rect 12816 10792 12850 10826
rect 12816 10702 12850 10736
rect 12816 10612 12850 10646
rect 12816 10522 12850 10556
rect 12816 10432 12850 10466
rect 12816 10342 12850 10376
rect 12816 10252 12850 10286
rect 14003 11152 14037 11186
rect 14003 11062 14037 11096
rect 14003 10972 14037 11006
rect 14003 10882 14037 10916
rect 14003 10792 14037 10826
rect 14003 10702 14037 10736
rect 14003 10612 14037 10646
rect 14003 10522 14037 10556
rect 14003 10432 14037 10466
rect 14003 10342 14037 10376
rect 14003 10252 14037 10286
rect 12816 10162 12850 10196
rect 14003 10162 14037 10196
rect 12912 10078 12946 10112
rect 13002 10078 13036 10112
rect 13092 10078 13126 10112
rect 13182 10078 13216 10112
rect 13272 10078 13306 10112
rect 13362 10078 13396 10112
rect 13452 10078 13486 10112
rect 13542 10078 13576 10112
rect 13632 10078 13666 10112
rect 13722 10078 13756 10112
rect 13812 10078 13846 10112
rect 13902 10078 13936 10112
rect 12816 9752 12850 9786
rect 12912 9775 12946 9809
rect 13002 9775 13036 9809
rect 13092 9775 13126 9809
rect 13182 9775 13216 9809
rect 13272 9775 13306 9809
rect 13362 9775 13396 9809
rect 13452 9775 13486 9809
rect 13542 9775 13576 9809
rect 13632 9775 13666 9809
rect 13722 9775 13756 9809
rect 13812 9775 13846 9809
rect 13902 9775 13936 9809
rect 14003 9752 14037 9786
rect 12816 9662 12850 9696
rect 12816 9572 12850 9606
rect 12816 9482 12850 9516
rect 12816 9392 12850 9426
rect 12816 9302 12850 9336
rect 12816 9212 12850 9246
rect 12816 9122 12850 9156
rect 12816 9032 12850 9066
rect 12816 8942 12850 8976
rect 12816 8852 12850 8886
rect 12816 8762 12850 8796
rect 14003 9662 14037 9696
rect 14003 9572 14037 9606
rect 14003 9482 14037 9516
rect 14003 9392 14037 9426
rect 14003 9302 14037 9336
rect 14003 9212 14037 9246
rect 14003 9122 14037 9156
rect 14003 9032 14037 9066
rect 14003 8942 14037 8976
rect 14003 8852 14037 8886
rect 14003 8762 14037 8796
rect 12816 8672 12850 8706
rect 14003 8672 14037 8706
rect 12912 8588 12946 8622
rect 13002 8588 13036 8622
rect 13092 8588 13126 8622
rect 13182 8588 13216 8622
rect 13272 8588 13306 8622
rect 13362 8588 13396 8622
rect 13452 8588 13486 8622
rect 13542 8588 13576 8622
rect 13632 8588 13666 8622
rect 13722 8588 13756 8622
rect 13812 8588 13846 8622
rect 13902 8588 13936 8622
rect 12806 8342 12840 8376
rect 12902 8365 12936 8399
rect 12992 8365 13026 8399
rect 13082 8365 13116 8399
rect 13172 8365 13206 8399
rect 13262 8365 13296 8399
rect 13352 8365 13386 8399
rect 13442 8365 13476 8399
rect 13532 8365 13566 8399
rect 13622 8365 13656 8399
rect 13712 8365 13746 8399
rect 13802 8365 13836 8399
rect 13892 8365 13926 8399
rect 13993 8342 14027 8376
rect 12806 8252 12840 8286
rect 12806 8162 12840 8196
rect 12806 8072 12840 8106
rect 12806 7982 12840 8016
rect 12806 7892 12840 7926
rect 12806 7802 12840 7836
rect 12806 7712 12840 7746
rect 12806 7622 12840 7656
rect 12806 7532 12840 7566
rect 12806 7442 12840 7476
rect 12806 7352 12840 7386
rect 13993 8252 14027 8286
rect 13993 8162 14027 8196
rect 13993 8072 14027 8106
rect 13993 7982 14027 8016
rect 20382 11448 20416 11482
rect 20382 11380 20416 11414
rect 20382 11312 20416 11346
rect 20382 11244 20416 11278
rect 20382 11176 20416 11210
rect 20382 11108 20416 11142
rect 20382 11040 20416 11074
rect 20382 10972 20416 11006
rect 20382 10904 20416 10938
rect 20382 10836 20416 10870
rect 20382 10768 20416 10802
rect 20382 10700 20416 10734
rect 20382 10632 20416 10666
rect 20382 10564 20416 10598
rect 20382 10496 20416 10530
rect 20382 10428 20416 10462
rect 20382 10360 20416 10394
rect 20382 10292 20416 10326
rect 20382 10224 20416 10258
rect 20382 10156 20416 10190
rect 20382 10088 20416 10122
rect 20382 10020 20416 10054
rect 20382 9952 20416 9986
rect 20382 9884 20416 9918
rect 20382 9816 20416 9850
rect 20382 9748 20416 9782
rect 20382 9680 20416 9714
rect 20382 9612 20416 9646
rect 20382 9544 20416 9578
rect 20382 9476 20416 9510
rect 20382 9408 20416 9442
rect 20382 9340 20416 9374
rect 20382 9272 20416 9306
rect 20382 9204 20416 9238
rect 20382 9136 20416 9170
rect 20382 9068 20416 9102
rect 20382 9000 20416 9034
rect 20382 8932 20416 8966
rect 20382 8864 20416 8898
rect 20382 8796 20416 8830
rect 20382 8728 20416 8762
rect 20382 8660 20416 8694
rect 20382 8592 20416 8626
rect 20382 8524 20416 8558
rect 20382 8456 20416 8490
rect 20382 8388 20416 8422
rect 20382 8320 20416 8354
rect 20382 8252 20416 8286
rect 20382 8184 20416 8218
rect 20382 8116 20416 8150
rect 20382 8048 20416 8082
rect 13993 7892 14027 7926
rect 13993 7802 14027 7836
rect 20382 7980 20416 8014
rect 20382 7912 20416 7946
rect 20382 7844 20416 7878
rect 20382 7776 20416 7810
rect 13993 7712 14027 7746
rect 13993 7622 14027 7656
rect 13993 7532 14027 7566
rect 13993 7442 14027 7476
rect 13993 7352 14027 7386
rect 12806 7262 12840 7296
rect 13993 7262 14027 7296
rect 12902 7178 12936 7212
rect 12992 7178 13026 7212
rect 13082 7178 13116 7212
rect 13172 7178 13206 7212
rect 13262 7178 13296 7212
rect 13352 7178 13386 7212
rect 13442 7178 13476 7212
rect 13532 7178 13566 7212
rect 13622 7178 13656 7212
rect 13712 7178 13746 7212
rect 13802 7178 13836 7212
rect 13892 7178 13926 7212
rect 16206 7206 16240 7240
rect 16274 7206 16308 7240
rect 16342 7206 16376 7240
rect 16410 7206 16444 7240
rect 16478 7206 16512 7240
rect 16546 7206 16580 7240
rect 16614 7206 16648 7240
rect 16682 7206 16716 7240
rect 16750 7206 16784 7240
rect 16818 7206 16852 7240
rect 16886 7206 16920 7240
rect 12806 6992 12840 7026
rect 12902 7015 12936 7049
rect 12992 7015 13026 7049
rect 13082 7015 13116 7049
rect 13172 7015 13206 7049
rect 13262 7015 13296 7049
rect 13352 7015 13386 7049
rect 13442 7015 13476 7049
rect 13532 7015 13566 7049
rect 13622 7015 13656 7049
rect 13712 7015 13746 7049
rect 13802 7015 13836 7049
rect 13892 7015 13926 7049
rect 13993 6992 14027 7026
rect 12806 6902 12840 6936
rect 12806 6812 12840 6846
rect 12806 6722 12840 6756
rect 12806 6632 12840 6666
rect 12806 6542 12840 6576
rect 12806 6452 12840 6486
rect 12806 6362 12840 6396
rect 12806 6272 12840 6306
rect 12806 6182 12840 6216
rect 12806 6092 12840 6126
rect 12806 6002 12840 6036
rect 13993 6902 14027 6936
rect 13993 6812 14027 6846
rect 13993 6722 14027 6756
rect 13993 6632 14027 6666
rect 13993 6542 14027 6576
rect 13993 6452 14027 6486
rect 13993 6362 14027 6396
rect 13993 6272 14027 6306
rect 13993 6182 14027 6216
rect 13993 6092 14027 6126
rect 13993 6002 14027 6036
rect 12806 5912 12840 5946
rect 13993 5912 14027 5946
rect 12902 5828 12936 5862
rect 12992 5828 13026 5862
rect 13082 5828 13116 5862
rect 13172 5828 13206 5862
rect 13262 5828 13296 5862
rect 13352 5828 13386 5862
rect 13442 5828 13476 5862
rect 13532 5828 13566 5862
rect 13622 5828 13656 5862
rect 13712 5828 13746 5862
rect 13802 5828 13836 5862
rect 13892 5828 13926 5862
rect 14456 7022 14490 7056
rect 14552 7045 14586 7079
rect 14642 7045 14676 7079
rect 14732 7045 14766 7079
rect 14822 7045 14856 7079
rect 14912 7045 14946 7079
rect 15002 7045 15036 7079
rect 15092 7045 15126 7079
rect 15182 7045 15216 7079
rect 15272 7045 15306 7079
rect 15362 7045 15396 7079
rect 15452 7045 15486 7079
rect 15542 7045 15576 7079
rect 15643 7022 15677 7056
rect 14456 6932 14490 6966
rect 14456 6842 14490 6876
rect 14456 6752 14490 6786
rect 14456 6662 14490 6696
rect 14456 6572 14490 6606
rect 14456 6482 14490 6516
rect 14456 6392 14490 6426
rect 14456 6302 14490 6336
rect 14456 6212 14490 6246
rect 14456 6122 14490 6156
rect 14456 6032 14490 6066
rect 15643 6932 15677 6966
rect 15643 6842 15677 6876
rect 15643 6752 15677 6786
rect 15643 6662 15677 6696
rect 15643 6572 15677 6606
rect 15643 6482 15677 6516
rect 15643 6392 15677 6426
rect 15643 6302 15677 6336
rect 15643 6212 15677 6246
rect 15643 6122 15677 6156
rect 15643 6032 15677 6066
rect 14456 5942 14490 5976
rect 15643 5942 15677 5976
rect 14552 5858 14586 5892
rect 14642 5858 14676 5892
rect 14732 5858 14766 5892
rect 14822 5858 14856 5892
rect 14912 5858 14946 5892
rect 15002 5858 15036 5892
rect 15092 5858 15126 5892
rect 15182 5858 15216 5892
rect 15272 5858 15306 5892
rect 15362 5858 15396 5892
rect 15452 5858 15486 5892
rect 15542 5858 15576 5892
rect 16080 7085 16114 7119
rect 16080 7017 16114 7051
rect 16080 6949 16114 6983
rect 16080 6881 16114 6915
rect 16080 6813 16114 6847
rect 16080 6745 16114 6779
rect 16080 6677 16114 6711
rect 16080 6609 16114 6643
rect 16080 6541 16114 6575
rect 16080 6473 16114 6507
rect 16080 6405 16114 6439
rect 16080 6337 16114 6371
rect 16080 6269 16114 6303
rect 16080 6201 16114 6235
rect 16080 6133 16114 6167
rect 16080 6065 16114 6099
rect 16080 5997 16114 6031
rect 16080 5929 16114 5963
rect 16080 5861 16114 5895
rect 16080 5793 16114 5827
rect 12806 5642 12840 5676
rect 12902 5665 12936 5699
rect 12992 5665 13026 5699
rect 13082 5665 13116 5699
rect 13172 5665 13206 5699
rect 13262 5665 13296 5699
rect 13352 5665 13386 5699
rect 13442 5665 13476 5699
rect 13532 5665 13566 5699
rect 13622 5665 13656 5699
rect 13712 5665 13746 5699
rect 13802 5665 13836 5699
rect 13892 5665 13926 5699
rect 13993 5642 14027 5676
rect 12806 5552 12840 5586
rect 12806 5462 12840 5496
rect 12806 5372 12840 5406
rect 12806 5282 12840 5316
rect 12806 5192 12840 5226
rect 12806 5102 12840 5136
rect 12806 5012 12840 5046
rect 12806 4922 12840 4956
rect 12806 4832 12840 4866
rect 12806 4742 12840 4776
rect 12806 4652 12840 4686
rect 13993 5552 14027 5586
rect 13993 5462 14027 5496
rect 13993 5372 14027 5406
rect 13993 5282 14027 5316
rect 13993 5192 14027 5226
rect 13993 5102 14027 5136
rect 13993 5012 14027 5046
rect 13993 4922 14027 4956
rect 13993 4832 14027 4866
rect 13993 4742 14027 4776
rect 13993 4652 14027 4686
rect 12806 4562 12840 4596
rect 13993 4562 14027 4596
rect 12902 4478 12936 4512
rect 12992 4478 13026 4512
rect 13082 4478 13116 4512
rect 13172 4478 13206 4512
rect 13262 4478 13296 4512
rect 13352 4478 13386 4512
rect 13442 4478 13476 4512
rect 13532 4478 13566 4512
rect 13622 4478 13656 4512
rect 13712 4478 13746 4512
rect 13802 4478 13836 4512
rect 13892 4478 13926 4512
rect 14456 5662 14490 5696
rect 14552 5685 14586 5719
rect 14642 5685 14676 5719
rect 14732 5685 14766 5719
rect 14822 5685 14856 5719
rect 14912 5685 14946 5719
rect 15002 5685 15036 5719
rect 15092 5685 15126 5719
rect 15182 5685 15216 5719
rect 15272 5685 15306 5719
rect 15362 5685 15396 5719
rect 15452 5685 15486 5719
rect 15542 5685 15576 5719
rect 15643 5662 15677 5696
rect 14456 5572 14490 5606
rect 14456 5482 14490 5516
rect 14456 5392 14490 5426
rect 14456 5302 14490 5336
rect 14456 5212 14490 5246
rect 14456 5122 14490 5156
rect 14456 5032 14490 5066
rect 14456 4942 14490 4976
rect 14456 4852 14490 4886
rect 14456 4762 14490 4796
rect 14456 4672 14490 4706
rect 15643 5572 15677 5606
rect 15643 5482 15677 5516
rect 15643 5392 15677 5426
rect 15643 5302 15677 5336
rect 15643 5212 15677 5246
rect 15643 5122 15677 5156
rect 15643 5032 15677 5066
rect 15643 4942 15677 4976
rect 15643 4852 15677 4886
rect 15643 4762 15677 4796
rect 15643 4672 15677 4706
rect 14456 4582 14490 4616
rect 15643 4582 15677 4616
rect 14552 4498 14586 4532
rect 14642 4498 14676 4532
rect 14732 4498 14766 4532
rect 14822 4498 14856 4532
rect 14912 4498 14946 4532
rect 15002 4498 15036 4532
rect 15092 4498 15126 4532
rect 15182 4498 15216 4532
rect 15272 4498 15306 4532
rect 15362 4498 15396 4532
rect 15452 4498 15486 4532
rect 15542 4498 15576 4532
rect 16080 5725 16114 5759
rect 16080 5657 16114 5691
rect 16080 5589 16114 5623
rect 16080 5521 16114 5555
rect 16080 5453 16114 5487
rect 16080 5385 16114 5419
rect 16080 5317 16114 5351
rect 16080 5249 16114 5283
rect 16080 5181 16114 5215
rect 16080 5113 16114 5147
rect 16080 5045 16114 5079
rect 16080 4977 16114 5011
rect 16080 4909 16114 4943
rect 16080 4841 16114 4875
rect 16080 4773 16114 4807
rect 16080 4705 16114 4739
rect 16080 4637 16114 4671
rect 17012 7085 17046 7119
rect 17012 7017 17046 7051
rect 17012 6949 17046 6983
rect 17012 6881 17046 6915
rect 17012 6813 17046 6847
rect 17012 6745 17046 6779
rect 17012 6677 17046 6711
rect 17012 6609 17046 6643
rect 17012 6541 17046 6575
rect 17012 6473 17046 6507
rect 17012 6405 17046 6439
rect 17012 6337 17046 6371
rect 17012 6269 17046 6303
rect 17012 6201 17046 6235
rect 17012 6133 17046 6167
rect 17012 6065 17046 6099
rect 17012 5997 17046 6031
rect 17012 5929 17046 5963
rect 17012 5861 17046 5895
rect 17012 5793 17046 5827
rect 17012 5725 17046 5759
rect 17012 5657 17046 5691
rect 17012 5589 17046 5623
rect 17012 5521 17046 5555
rect 17012 5453 17046 5487
rect 17012 5385 17046 5419
rect 17012 5317 17046 5351
rect 17012 5249 17046 5283
rect 17012 5181 17046 5215
rect 17012 5113 17046 5147
rect 17012 5045 17046 5079
rect 17012 4977 17046 5011
rect 17012 4909 17046 4943
rect 17012 4841 17046 4875
rect 17012 4773 17046 4807
rect 17012 4705 17046 4739
rect 17012 4637 17046 4671
rect 16206 4516 16240 4550
rect 16274 4516 16308 4550
rect 16342 4516 16376 4550
rect 16410 4516 16444 4550
rect 16478 4516 16512 4550
rect 16546 4516 16580 4550
rect 16614 4516 16648 4550
rect 16682 4516 16716 4550
rect 16750 4516 16784 4550
rect 16818 4516 16852 4550
rect 16886 4516 16920 4550
rect 20382 7708 20416 7742
rect 20382 7640 20416 7674
rect 20382 7572 20416 7606
rect 20382 7504 20416 7538
rect 20382 7436 20416 7470
rect 20382 7368 20416 7402
rect 20382 7300 20416 7334
rect 20382 7232 20416 7266
rect 20382 7164 20416 7198
rect 20382 7096 20416 7130
rect 20382 7028 20416 7062
rect 20382 6960 20416 6994
rect 20382 6892 20416 6926
rect 20382 6824 20416 6858
rect 20382 6756 20416 6790
rect 20382 6688 20416 6722
rect 20382 6620 20416 6654
rect 20382 6552 20416 6586
rect 20382 6484 20416 6518
rect 20382 6416 20416 6450
rect 20382 6348 20416 6382
rect 20382 6280 20416 6314
rect 20382 6212 20416 6246
rect 20382 6144 20416 6178
rect 20382 6076 20416 6110
rect 20382 6008 20416 6042
rect 20382 5940 20416 5974
rect 20382 5872 20416 5906
rect 20382 5804 20416 5838
rect 20382 5736 20416 5770
rect 20382 5668 20416 5702
rect 20382 5600 20416 5634
rect 20382 5532 20416 5566
rect 20382 5464 20416 5498
rect 20382 5396 20416 5430
rect 20382 5328 20416 5362
rect 20382 5260 20416 5294
rect 20382 5192 20416 5226
rect 20382 5124 20416 5158
rect 20382 5056 20416 5090
rect 20382 4988 20416 5022
rect 20382 4920 20416 4954
rect 20382 4852 20416 4886
rect 20382 4784 20416 4818
rect 20382 4716 20416 4750
rect 21632 14440 21666 14474
rect 21632 14372 21666 14406
rect 21632 14304 21666 14338
rect 21632 14236 21666 14270
rect 21632 14168 21666 14202
rect 21632 14100 21666 14134
rect 21632 14032 21666 14066
rect 21632 13964 21666 13998
rect 21632 13896 21666 13930
rect 21632 13828 21666 13862
rect 21632 13760 21666 13794
rect 21632 13692 21666 13726
rect 21632 13624 21666 13658
rect 28834 14561 28868 14595
rect 28834 14493 28868 14527
rect 28834 14425 28868 14459
rect 28834 14357 28868 14391
rect 28834 14289 28868 14323
rect 28834 14221 28868 14255
rect 28834 14153 28868 14187
rect 28834 14085 28868 14119
rect 28834 14017 28868 14051
rect 28834 13949 28868 13983
rect 28834 13881 28868 13915
rect 28834 13813 28868 13847
rect 28834 13745 28868 13779
rect 29766 15241 29800 15275
rect 29766 15173 29800 15207
rect 29766 15105 29800 15139
rect 29766 15037 29800 15071
rect 29766 14969 29800 15003
rect 29766 14901 29800 14935
rect 29766 14833 29800 14867
rect 29766 14765 29800 14799
rect 29766 14697 29800 14731
rect 29766 14629 29800 14663
rect 29766 14561 29800 14595
rect 29766 14493 29800 14527
rect 29766 14425 29800 14459
rect 29766 14357 29800 14391
rect 29766 14289 29800 14323
rect 29766 14221 29800 14255
rect 29766 14153 29800 14187
rect 29766 14085 29800 14119
rect 29766 14017 29800 14051
rect 29766 13949 29800 13983
rect 29766 13881 29800 13915
rect 29766 13813 29800 13847
rect 29766 13745 29800 13779
rect 28960 13628 28994 13662
rect 29028 13628 29062 13662
rect 29096 13628 29130 13662
rect 29164 13628 29198 13662
rect 29232 13628 29266 13662
rect 29300 13628 29334 13662
rect 29368 13628 29402 13662
rect 29436 13628 29470 13662
rect 29504 13628 29538 13662
rect 29572 13628 29606 13662
rect 29640 13628 29674 13662
rect 37749 15344 37783 15378
rect 37749 15276 37783 15310
rect 37749 15208 37783 15242
rect 37749 15140 37783 15174
rect 37749 15072 37783 15106
rect 37749 15004 37783 15038
rect 37749 14936 37783 14970
rect 37749 14868 37783 14902
rect 37749 14800 37783 14834
rect 37749 14732 37783 14766
rect 37749 14664 37783 14698
rect 37749 14596 37783 14630
rect 37749 14528 37783 14562
rect 37749 14460 37783 14494
rect 37749 14392 37783 14426
rect 37749 14324 37783 14358
rect 37749 14256 37783 14290
rect 37749 14188 37783 14222
rect 37749 14120 37783 14154
rect 37749 14052 37783 14086
rect 37749 13984 37783 14018
rect 37749 13916 37783 13950
rect 37749 13848 37783 13882
rect 37749 13780 37783 13814
rect 37749 13712 37783 13746
rect 37749 13644 37783 13678
rect 21632 13556 21666 13590
rect 21632 13488 21666 13522
rect 37749 13576 37783 13610
rect 41089 15576 41123 15610
rect 41089 15508 41123 15542
rect 41089 15440 41123 15474
rect 41089 15372 41123 15406
rect 41089 15304 41123 15338
rect 41089 15236 41123 15270
rect 41089 15168 41123 15202
rect 41089 15100 41123 15134
rect 41089 15032 41123 15066
rect 41089 14964 41123 14998
rect 41089 14896 41123 14930
rect 41089 14828 41123 14862
rect 41089 14760 41123 14794
rect 41089 14692 41123 14726
rect 41089 14624 41123 14658
rect 41089 14556 41123 14590
rect 41089 14488 41123 14522
rect 41089 14420 41123 14454
rect 41089 14352 41123 14386
rect 41089 14284 41123 14318
rect 41089 14216 41123 14250
rect 41089 14148 41123 14182
rect 41089 14080 41123 14114
rect 41089 14012 41123 14046
rect 41089 13944 41123 13978
rect 41089 13876 41123 13910
rect 41089 13808 41123 13842
rect 41089 13740 41123 13774
rect 41089 13672 41123 13706
rect 41089 13604 41123 13638
rect 37749 13508 37783 13542
rect 21632 13420 21666 13454
rect 21632 13352 21666 13386
rect 21632 13284 21666 13318
rect 21632 13216 21666 13250
rect 21632 13148 21666 13182
rect 21632 13080 21666 13114
rect 21632 13012 21666 13046
rect 21632 12944 21666 12978
rect 21632 12876 21666 12910
rect 21632 12808 21666 12842
rect 21632 12740 21666 12774
rect 21632 12672 21666 12706
rect 21632 12604 21666 12638
rect 21632 12536 21666 12570
rect 21632 12468 21666 12502
rect 21632 12400 21666 12434
rect 21632 12332 21666 12366
rect 21632 12264 21666 12298
rect 21632 12196 21666 12230
rect 21632 12128 21666 12162
rect 21632 12060 21666 12094
rect 21632 11992 21666 12026
rect 21632 11924 21666 11958
rect 21632 11856 21666 11890
rect 21632 11788 21666 11822
rect 21632 11720 21666 11754
rect 21632 11652 21666 11686
rect 21632 11584 21666 11618
rect 21632 11516 21666 11550
rect 21632 11448 21666 11482
rect 21632 11380 21666 11414
rect 21632 11312 21666 11346
rect 21632 11244 21666 11278
rect 21632 11176 21666 11210
rect 21632 11108 21666 11142
rect 21632 11040 21666 11074
rect 21632 10972 21666 11006
rect 21632 10904 21666 10938
rect 21632 10836 21666 10870
rect 21632 10768 21666 10802
rect 21632 10700 21666 10734
rect 21632 10632 21666 10666
rect 21632 10564 21666 10598
rect 21632 10496 21666 10530
rect 21632 10428 21666 10462
rect 21632 10360 21666 10394
rect 21632 10292 21666 10326
rect 21632 10224 21666 10258
rect 21632 10156 21666 10190
rect 21632 10088 21666 10122
rect 21632 10020 21666 10054
rect 21632 9952 21666 9986
rect 21632 9884 21666 9918
rect 21632 9816 21666 9850
rect 21632 9748 21666 9782
rect 21632 9680 21666 9714
rect 21632 9612 21666 9646
rect 21632 9544 21666 9578
rect 21632 9476 21666 9510
rect 21632 9408 21666 9442
rect 21632 9340 21666 9374
rect 21632 9272 21666 9306
rect 21632 9204 21666 9238
rect 21632 9136 21666 9170
rect 21632 9068 21666 9102
rect 21632 9000 21666 9034
rect 21632 8932 21666 8966
rect 26524 13440 26558 13474
rect 26592 13440 26626 13474
rect 26660 13440 26694 13474
rect 26728 13440 26762 13474
rect 26796 13440 26830 13474
rect 26864 13440 26898 13474
rect 26932 13440 26966 13474
rect 27000 13440 27034 13474
rect 27068 13440 27102 13474
rect 27136 13440 27170 13474
rect 27204 13440 27238 13474
rect 26398 13329 26432 13363
rect 26398 13261 26432 13295
rect 26398 13193 26432 13227
rect 26398 13125 26432 13159
rect 26398 13057 26432 13091
rect 26398 12989 26432 13023
rect 26398 12921 26432 12955
rect 26398 12853 26432 12887
rect 26398 12785 26432 12819
rect 26398 12717 26432 12751
rect 26398 12649 26432 12683
rect 26398 12581 26432 12615
rect 26398 12513 26432 12547
rect 26398 12445 26432 12479
rect 26398 12377 26432 12411
rect 26398 12309 26432 12343
rect 26398 12241 26432 12275
rect 26398 12173 26432 12207
rect 26398 12105 26432 12139
rect 26398 12037 26432 12071
rect 26398 11969 26432 12003
rect 26398 11901 26432 11935
rect 26398 11833 26432 11867
rect 26398 11765 26432 11799
rect 26398 11697 26432 11731
rect 26398 11629 26432 11663
rect 26398 11561 26432 11595
rect 26398 11493 26432 11527
rect 26398 11425 26432 11459
rect 26398 11357 26432 11391
rect 26398 11289 26432 11323
rect 26398 11221 26432 11255
rect 26398 11153 26432 11187
rect 26398 11085 26432 11119
rect 26398 11017 26432 11051
rect 26398 10949 26432 10983
rect 26398 10881 26432 10915
rect 26398 10813 26432 10847
rect 26398 10745 26432 10779
rect 26398 10677 26432 10711
rect 26398 10609 26432 10643
rect 26398 10541 26432 10575
rect 26398 10473 26432 10507
rect 26398 10405 26432 10439
rect 26398 10337 26432 10371
rect 26398 10269 26432 10303
rect 26398 10201 26432 10235
rect 26398 10133 26432 10167
rect 26398 10065 26432 10099
rect 26398 9997 26432 10031
rect 26398 9929 26432 9963
rect 26398 9861 26432 9895
rect 26398 9793 26432 9827
rect 26398 9725 26432 9759
rect 26398 9657 26432 9691
rect 26398 9589 26432 9623
rect 26398 9521 26432 9555
rect 26398 9453 26432 9487
rect 26398 9385 26432 9419
rect 26398 9317 26432 9351
rect 26398 9249 26432 9283
rect 26398 9181 26432 9215
rect 26398 9113 26432 9147
rect 26398 9045 26432 9079
rect 26398 8977 26432 9011
rect 21632 8864 21666 8898
rect 21632 8796 21666 8830
rect 21632 8728 21666 8762
rect 21632 8660 21666 8694
rect 21632 8592 21666 8626
rect 21632 8524 21666 8558
rect 21632 8456 21666 8490
rect 21632 8388 21666 8422
rect 21632 8320 21666 8354
rect 21632 8252 21666 8286
rect 21632 8184 21666 8218
rect 21632 8116 21666 8150
rect 21632 8048 21666 8082
rect 26398 8909 26432 8943
rect 26398 8841 26432 8875
rect 26398 8773 26432 8807
rect 26398 8705 26432 8739
rect 26398 8637 26432 8671
rect 26398 8569 26432 8603
rect 26398 8501 26432 8535
rect 26398 8433 26432 8467
rect 26398 8365 26432 8399
rect 26398 8297 26432 8331
rect 26398 8229 26432 8263
rect 26398 8161 26432 8195
rect 26398 8093 26432 8127
rect 21632 7980 21666 8014
rect 21632 7912 21666 7946
rect 21632 7844 21666 7878
rect 21632 7776 21666 7810
rect 21632 7708 21666 7742
rect 21632 7640 21666 7674
rect 21632 7572 21666 7606
rect 21632 7504 21666 7538
rect 21632 7436 21666 7470
rect 21632 7368 21666 7402
rect 21632 7300 21666 7334
rect 21632 7232 21666 7266
rect 21632 7164 21666 7198
rect 21632 7096 21666 7130
rect 21632 7028 21666 7062
rect 21632 6960 21666 6994
rect 21632 6892 21666 6926
rect 21632 6824 21666 6858
rect 21632 6756 21666 6790
rect 21632 6688 21666 6722
rect 21632 6620 21666 6654
rect 21632 6552 21666 6586
rect 21632 6484 21666 6518
rect 21632 6416 21666 6450
rect 21632 6348 21666 6382
rect 21632 6280 21666 6314
rect 21632 6212 21666 6246
rect 21632 6144 21666 6178
rect 21632 6076 21666 6110
rect 21632 6008 21666 6042
rect 21632 5940 21666 5974
rect 21632 5872 21666 5906
rect 21632 5804 21666 5838
rect 21632 5736 21666 5770
rect 21632 5668 21666 5702
rect 21632 5600 21666 5634
rect 21632 5532 21666 5566
rect 21632 5464 21666 5498
rect 21632 5396 21666 5430
rect 21632 5328 21666 5362
rect 21632 5260 21666 5294
rect 21632 5192 21666 5226
rect 21632 5124 21666 5158
rect 21632 5056 21666 5090
rect 21632 4988 21666 5022
rect 21632 4920 21666 4954
rect 21632 4852 21666 4886
rect 21632 4784 21666 4818
rect 21632 4716 21666 4750
rect 20497 4590 20531 4624
rect 20565 4590 20599 4624
rect 20633 4590 20667 4624
rect 20701 4590 20735 4624
rect 20769 4590 20803 4624
rect 20837 4590 20871 4624
rect 20905 4590 20939 4624
rect 20973 4590 21007 4624
rect 21041 4590 21075 4624
rect 21109 4590 21143 4624
rect 21177 4590 21211 4624
rect 21245 4590 21279 4624
rect 21313 4590 21347 4624
rect 21381 4590 21415 4624
rect 21449 4590 21483 4624
rect 21517 4590 21551 4624
rect 26398 8025 26432 8059
rect 26398 7957 26432 7991
rect 26398 7889 26432 7923
rect 26398 7821 26432 7855
rect 26398 7753 26432 7787
rect 26398 7685 26432 7719
rect 26398 7617 26432 7651
rect 26398 7549 26432 7583
rect 26398 7481 26432 7515
rect 26398 7413 26432 7447
rect 26398 7345 26432 7379
rect 26398 7277 26432 7311
rect 26398 7209 26432 7243
rect 26398 7141 26432 7175
rect 26398 7073 26432 7107
rect 26398 7005 26432 7039
rect 26398 6937 26432 6971
rect 26398 6869 26432 6903
rect 26398 6801 26432 6835
rect 26398 6733 26432 6767
rect 26398 6665 26432 6699
rect 26398 6597 26432 6631
rect 26398 6529 26432 6563
rect 26398 6461 26432 6495
rect 26398 6393 26432 6427
rect 26398 6325 26432 6359
rect 26398 6257 26432 6291
rect 26398 6189 26432 6223
rect 26398 6121 26432 6155
rect 26398 6053 26432 6087
rect 26398 5985 26432 6019
rect 26398 5917 26432 5951
rect 26398 5849 26432 5883
rect 26398 5781 26432 5815
rect 26398 5713 26432 5747
rect 26398 5645 26432 5679
rect 26398 5577 26432 5611
rect 26398 5509 26432 5543
rect 26398 5441 26432 5475
rect 26398 5373 26432 5407
rect 26398 5305 26432 5339
rect 26398 5237 26432 5271
rect 26398 5169 26432 5203
rect 26398 5101 26432 5135
rect 26398 5033 26432 5067
rect 26398 4965 26432 4999
rect 26398 4897 26432 4931
rect 26398 4829 26432 4863
rect 26398 4761 26432 4795
rect 26398 4693 26432 4727
rect 26398 4625 26432 4659
rect 26398 4557 26432 4591
rect 26398 4489 26432 4523
rect 26398 4421 26432 4455
rect 26398 4353 26432 4387
rect 26398 4285 26432 4319
rect 26398 4217 26432 4251
rect 26398 4149 26432 4183
rect 26398 4081 26432 4115
rect 26398 4013 26432 4047
rect 26398 3945 26432 3979
rect 26398 3877 26432 3911
rect 26398 3809 26432 3843
rect 26398 3741 26432 3775
rect 26398 3673 26432 3707
rect 26398 3605 26432 3639
rect 26398 3537 26432 3571
rect 26398 3469 26432 3503
rect 26398 3401 26432 3435
rect 26398 3333 26432 3367
rect 26398 3265 26432 3299
rect 26398 3197 26432 3231
rect 26398 3129 26432 3163
rect 26398 3061 26432 3095
rect 27330 13329 27364 13363
rect 27330 13261 27364 13295
rect 27330 13193 27364 13227
rect 27330 13125 27364 13159
rect 27330 13057 27364 13091
rect 27330 12989 27364 13023
rect 27330 12921 27364 12955
rect 27330 12853 27364 12887
rect 27330 12785 27364 12819
rect 27330 12717 27364 12751
rect 27330 12649 27364 12683
rect 27330 12581 27364 12615
rect 27330 12513 27364 12547
rect 27330 12445 27364 12479
rect 27330 12377 27364 12411
rect 27330 12309 27364 12343
rect 27330 12241 27364 12275
rect 27330 12173 27364 12207
rect 27330 12105 27364 12139
rect 27330 12037 27364 12071
rect 27330 11969 27364 12003
rect 27330 11901 27364 11935
rect 27330 11833 27364 11867
rect 27330 11765 27364 11799
rect 27330 11697 27364 11731
rect 27330 11629 27364 11663
rect 27330 11561 27364 11595
rect 27330 11493 27364 11527
rect 27330 11425 27364 11459
rect 27330 11357 27364 11391
rect 27330 11289 27364 11323
rect 27330 11221 27364 11255
rect 27330 11153 27364 11187
rect 27330 11085 27364 11119
rect 27330 11017 27364 11051
rect 27330 10949 27364 10983
rect 27330 10881 27364 10915
rect 27330 10813 27364 10847
rect 27330 10745 27364 10779
rect 27330 10677 27364 10711
rect 27330 10609 27364 10643
rect 27330 10541 27364 10575
rect 27330 10473 27364 10507
rect 27330 10405 27364 10439
rect 27330 10337 27364 10371
rect 27330 10269 27364 10303
rect 27330 10201 27364 10235
rect 27330 10133 27364 10167
rect 27330 10065 27364 10099
rect 27330 9997 27364 10031
rect 27330 9929 27364 9963
rect 27330 9861 27364 9895
rect 27330 9793 27364 9827
rect 27330 9725 27364 9759
rect 27330 9657 27364 9691
rect 27330 9589 27364 9623
rect 27330 9521 27364 9555
rect 27330 9453 27364 9487
rect 27330 9385 27364 9419
rect 27330 9317 27364 9351
rect 27330 9249 27364 9283
rect 27330 9181 27364 9215
rect 27330 9113 27364 9147
rect 27330 9045 27364 9079
rect 27330 8977 27364 9011
rect 27330 8909 27364 8943
rect 27330 8841 27364 8875
rect 27330 8773 27364 8807
rect 27330 8705 27364 8739
rect 27330 8637 27364 8671
rect 27330 8569 27364 8603
rect 27330 8501 27364 8535
rect 27330 8433 27364 8467
rect 27330 8365 27364 8399
rect 27330 8297 27364 8331
rect 27330 8229 27364 8263
rect 27330 8161 27364 8195
rect 27330 8093 27364 8127
rect 27330 8025 27364 8059
rect 27330 7957 27364 7991
rect 27330 7889 27364 7923
rect 27330 7821 27364 7855
rect 27330 7753 27364 7787
rect 27330 7685 27364 7719
rect 27330 7617 27364 7651
rect 27330 7549 27364 7583
rect 27330 7481 27364 7515
rect 27330 7413 27364 7447
rect 27330 7345 27364 7379
rect 27330 7277 27364 7311
rect 27330 7209 27364 7243
rect 27330 7141 27364 7175
rect 27330 7073 27364 7107
rect 27330 7005 27364 7039
rect 27330 6937 27364 6971
rect 27330 6869 27364 6903
rect 27330 6801 27364 6835
rect 27330 6733 27364 6767
rect 27330 6665 27364 6699
rect 27330 6597 27364 6631
rect 27330 6529 27364 6563
rect 27330 6461 27364 6495
rect 27330 6393 27364 6427
rect 27330 6325 27364 6359
rect 27686 13424 27720 13458
rect 27754 13424 27788 13458
rect 27822 13424 27856 13458
rect 27890 13424 27924 13458
rect 27958 13424 27992 13458
rect 28026 13424 28060 13458
rect 28094 13424 28128 13458
rect 28162 13424 28196 13458
rect 28230 13424 28264 13458
rect 28298 13424 28332 13458
rect 28366 13424 28400 13458
rect 28434 13424 28468 13458
rect 28502 13424 28536 13458
rect 28570 13424 28604 13458
rect 28638 13424 28672 13458
rect 28706 13424 28740 13458
rect 28774 13424 28808 13458
rect 28842 13424 28876 13458
rect 28910 13424 28944 13458
rect 28978 13424 29012 13458
rect 29046 13424 29080 13458
rect 29114 13424 29148 13458
rect 29182 13424 29216 13458
rect 29250 13424 29284 13458
rect 29318 13424 29352 13458
rect 29386 13424 29420 13458
rect 29454 13424 29488 13458
rect 29522 13424 29556 13458
rect 29590 13424 29624 13458
rect 29658 13424 29692 13458
rect 27570 13313 27604 13347
rect 27570 13245 27604 13279
rect 27570 13177 27604 13211
rect 27570 13109 27604 13143
rect 27570 13041 27604 13075
rect 27570 12973 27604 13007
rect 27570 12905 27604 12939
rect 27570 12837 27604 12871
rect 27570 12769 27604 12803
rect 27570 12701 27604 12735
rect 27570 12633 27604 12667
rect 27570 12565 27604 12599
rect 27570 12497 27604 12531
rect 27570 12429 27604 12463
rect 27570 12361 27604 12395
rect 27570 12293 27604 12327
rect 27570 12225 27604 12259
rect 27570 12157 27604 12191
rect 27570 12089 27604 12123
rect 27570 12021 27604 12055
rect 27570 11953 27604 11987
rect 27570 11885 27604 11919
rect 27570 11817 27604 11851
rect 27570 11749 27604 11783
rect 27570 11681 27604 11715
rect 27570 11613 27604 11647
rect 27570 11545 27604 11579
rect 27570 11477 27604 11511
rect 27570 11409 27604 11443
rect 27570 11341 27604 11375
rect 27570 11273 27604 11307
rect 27570 11205 27604 11239
rect 27570 11137 27604 11171
rect 27570 11069 27604 11103
rect 27570 11001 27604 11035
rect 27570 10933 27604 10967
rect 27570 10865 27604 10899
rect 27570 10797 27604 10831
rect 27570 10729 27604 10763
rect 27570 10661 27604 10695
rect 27570 10593 27604 10627
rect 27570 10525 27604 10559
rect 27570 10457 27604 10491
rect 27570 10389 27604 10423
rect 27570 10321 27604 10355
rect 27570 10253 27604 10287
rect 27570 10185 27604 10219
rect 27570 10117 27604 10151
rect 27570 10049 27604 10083
rect 27570 9981 27604 10015
rect 27570 9913 27604 9947
rect 27570 9845 27604 9879
rect 27570 9777 27604 9811
rect 27570 9709 27604 9743
rect 27570 9641 27604 9675
rect 27570 9573 27604 9607
rect 27570 9505 27604 9539
rect 27570 9437 27604 9471
rect 27570 9369 27604 9403
rect 27570 9301 27604 9335
rect 27570 9233 27604 9267
rect 27570 9165 27604 9199
rect 27570 9097 27604 9131
rect 27570 9029 27604 9063
rect 27570 8961 27604 8995
rect 27570 8893 27604 8927
rect 27570 8825 27604 8859
rect 27570 8757 27604 8791
rect 27570 8689 27604 8723
rect 27570 8621 27604 8655
rect 27570 8553 27604 8587
rect 27570 8485 27604 8519
rect 27570 8417 27604 8451
rect 27570 8349 27604 8383
rect 27570 8281 27604 8315
rect 27570 8213 27604 8247
rect 27570 8145 27604 8179
rect 27570 8077 27604 8111
rect 27570 8009 27604 8043
rect 27570 7941 27604 7975
rect 27570 7873 27604 7907
rect 27570 7805 27604 7839
rect 27570 7737 27604 7771
rect 27570 7669 27604 7703
rect 27570 7601 27604 7635
rect 27570 7533 27604 7567
rect 27570 7465 27604 7499
rect 27570 7397 27604 7431
rect 27570 7329 27604 7363
rect 27570 7261 27604 7295
rect 27570 7193 27604 7227
rect 27570 7125 27604 7159
rect 27570 7057 27604 7091
rect 27570 6989 27604 7023
rect 27570 6921 27604 6955
rect 27570 6853 27604 6887
rect 27570 6785 27604 6819
rect 27570 6717 27604 6751
rect 27570 6649 27604 6683
rect 27570 6581 27604 6615
rect 27570 6513 27604 6547
rect 27570 6445 27604 6479
rect 29774 13313 29808 13347
rect 29774 13245 29808 13279
rect 29774 13177 29808 13211
rect 29774 13109 29808 13143
rect 29774 13041 29808 13075
rect 29774 12973 29808 13007
rect 29774 12905 29808 12939
rect 37749 13440 37783 13474
rect 37749 13372 37783 13406
rect 41089 13536 41123 13570
rect 41089 13468 41123 13502
rect 41089 13400 41123 13434
rect 37749 13304 37783 13338
rect 37749 13236 37783 13270
rect 37749 13168 37783 13202
rect 37749 13100 37783 13134
rect 41089 13332 41123 13366
rect 41089 13264 41123 13298
rect 41089 13196 41123 13230
rect 41089 13128 41123 13162
rect 41089 13060 41123 13094
rect 41696 15751 41730 15785
rect 41764 15751 41798 15785
rect 41582 15630 41616 15664
rect 41582 15562 41616 15596
rect 41582 15494 41616 15528
rect 41582 15426 41616 15460
rect 41582 15358 41616 15392
rect 41582 15290 41616 15324
rect 41582 15222 41616 15256
rect 41582 15154 41616 15188
rect 41582 15086 41616 15120
rect 41582 15018 41616 15052
rect 41582 14950 41616 14984
rect 41582 14882 41616 14916
rect 41582 14814 41616 14848
rect 41582 14746 41616 14780
rect 41582 14678 41616 14712
rect 41582 14610 41616 14644
rect 41582 14542 41616 14576
rect 41582 14474 41616 14508
rect 41582 14406 41616 14440
rect 41582 14338 41616 14372
rect 41582 14270 41616 14304
rect 41582 14202 41616 14236
rect 41582 14134 41616 14168
rect 41582 14066 41616 14100
rect 41582 13998 41616 14032
rect 41582 13930 41616 13964
rect 41582 13862 41616 13896
rect 41582 13794 41616 13828
rect 41582 13726 41616 13760
rect 41582 13658 41616 13692
rect 41582 13590 41616 13624
rect 41582 13522 41616 13556
rect 41582 13454 41616 13488
rect 41582 13386 41616 13420
rect 41582 13318 41616 13352
rect 41582 13250 41616 13284
rect 41582 13182 41616 13216
rect 41878 15630 41912 15664
rect 41878 15562 41912 15596
rect 41878 15494 41912 15528
rect 41878 15426 41912 15460
rect 41878 15358 41912 15392
rect 41878 15290 41912 15324
rect 41878 15222 41912 15256
rect 41878 15154 41912 15188
rect 41878 15086 41912 15120
rect 41878 15018 41912 15052
rect 41878 14950 41912 14984
rect 41878 14882 41912 14916
rect 41878 14814 41912 14848
rect 41878 14746 41912 14780
rect 41878 14678 41912 14712
rect 41878 14610 41912 14644
rect 41878 14542 41912 14576
rect 41878 14474 41912 14508
rect 41878 14406 41912 14440
rect 41878 14338 41912 14372
rect 41878 14270 41912 14304
rect 41878 14202 41912 14236
rect 41878 14134 41912 14168
rect 41878 14066 41912 14100
rect 41878 13998 41912 14032
rect 41878 13930 41912 13964
rect 41878 13862 41912 13896
rect 41878 13794 41912 13828
rect 41878 13726 41912 13760
rect 41878 13658 41912 13692
rect 41878 13590 41912 13624
rect 41878 13522 41912 13556
rect 41878 13454 41912 13488
rect 41878 13386 41912 13420
rect 41878 13318 41912 13352
rect 41878 13250 41912 13284
rect 41878 13182 41912 13216
rect 41696 13061 41730 13095
rect 41764 13061 41798 13095
rect 38022 12952 38056 12986
rect 38090 12952 38124 12986
rect 38158 12952 38192 12986
rect 38226 12952 38260 12986
rect 38294 12952 38328 12986
rect 38362 12952 38396 12986
rect 38430 12952 38464 12986
rect 38498 12952 38532 12986
rect 38566 12952 38600 12986
rect 38634 12952 38668 12986
rect 38702 12952 38736 12986
rect 38770 12952 38804 12986
rect 38838 12952 38872 12986
rect 38906 12952 38940 12986
rect 38974 12952 39008 12986
rect 39042 12952 39076 12986
rect 39110 12952 39144 12986
rect 39178 12952 39212 12986
rect 39246 12952 39280 12986
rect 39314 12952 39348 12986
rect 39382 12952 39416 12986
rect 39450 12952 39484 12986
rect 39518 12952 39552 12986
rect 39586 12952 39620 12986
rect 39654 12952 39688 12986
rect 39722 12952 39756 12986
rect 39790 12952 39824 12986
rect 39858 12952 39892 12986
rect 39926 12952 39960 12986
rect 39994 12952 40028 12986
rect 40062 12952 40096 12986
rect 40130 12952 40164 12986
rect 40198 12952 40232 12986
rect 40266 12952 40300 12986
rect 40334 12952 40368 12986
rect 40402 12952 40436 12986
rect 40470 12952 40504 12986
rect 40538 12952 40572 12986
rect 40606 12952 40640 12986
rect 40674 12952 40708 12986
rect 40742 12952 40776 12986
rect 40810 12952 40844 12986
rect 40878 12952 40912 12986
rect 40946 12952 40980 12986
rect 29774 12837 29808 12871
rect 29774 12769 29808 12803
rect 29774 12701 29808 12735
rect 29774 12633 29808 12667
rect 29774 12565 29808 12599
rect 29774 12497 29808 12531
rect 29774 12429 29808 12463
rect 29774 12361 29808 12395
rect 29774 12293 29808 12327
rect 29774 12225 29808 12259
rect 29774 12157 29808 12191
rect 29774 12089 29808 12123
rect 29774 12021 29808 12055
rect 29774 11953 29808 11987
rect 29774 11885 29808 11919
rect 29774 11817 29808 11851
rect 29774 11749 29808 11783
rect 29774 11681 29808 11715
rect 29774 11613 29808 11647
rect 29774 11545 29808 11579
rect 29774 11477 29808 11511
rect 29774 11409 29808 11443
rect 29774 11341 29808 11375
rect 29774 11273 29808 11307
rect 29774 11205 29808 11239
rect 29774 11137 29808 11171
rect 29774 11069 29808 11103
rect 29774 11001 29808 11035
rect 29774 10933 29808 10967
rect 29774 10865 29808 10899
rect 29774 10797 29808 10831
rect 29774 10729 29808 10763
rect 29774 10661 29808 10695
rect 29774 10593 29808 10627
rect 29774 10525 29808 10559
rect 29774 10457 29808 10491
rect 29774 10389 29808 10423
rect 29774 10321 29808 10355
rect 29774 10253 29808 10287
rect 29774 10185 29808 10219
rect 29774 10117 29808 10151
rect 29774 10049 29808 10083
rect 29774 9981 29808 10015
rect 29774 9913 29808 9947
rect 29774 9845 29808 9879
rect 29774 9777 29808 9811
rect 29774 9709 29808 9743
rect 29774 9641 29808 9675
rect 29774 9573 29808 9607
rect 29774 9505 29808 9539
rect 29774 9437 29808 9471
rect 29774 9369 29808 9403
rect 29774 9301 29808 9335
rect 29774 9233 29808 9267
rect 29774 9165 29808 9199
rect 29774 9097 29808 9131
rect 29774 9029 29808 9063
rect 29774 8961 29808 8995
rect 29774 8893 29808 8927
rect 29774 8825 29808 8859
rect 29774 8757 29808 8791
rect 29774 8689 29808 8723
rect 29774 8621 29808 8655
rect 29774 8553 29808 8587
rect 29774 8485 29808 8519
rect 29774 8417 29808 8451
rect 29774 8349 29808 8383
rect 29774 8281 29808 8315
rect 29774 8213 29808 8247
rect 29774 8145 29808 8179
rect 29774 8077 29808 8111
rect 29774 8009 29808 8043
rect 29774 7941 29808 7975
rect 29774 7873 29808 7907
rect 29774 7805 29808 7839
rect 29774 7737 29808 7771
rect 29774 7669 29808 7703
rect 29774 7601 29808 7635
rect 29774 7533 29808 7567
rect 29774 7465 29808 7499
rect 29774 7397 29808 7431
rect 29774 7329 29808 7363
rect 29774 7261 29808 7295
rect 29774 7193 29808 7227
rect 29774 7125 29808 7159
rect 29774 7057 29808 7091
rect 29774 6989 29808 7023
rect 29774 6921 29808 6955
rect 29774 6853 29808 6887
rect 29774 6785 29808 6819
rect 29774 6717 29808 6751
rect 29774 6649 29808 6683
rect 29774 6581 29808 6615
rect 29774 6513 29808 6547
rect 29774 6445 29808 6479
rect 27686 6334 27720 6368
rect 27754 6334 27788 6368
rect 27822 6334 27856 6368
rect 27890 6334 27924 6368
rect 27958 6334 27992 6368
rect 28026 6334 28060 6368
rect 28094 6334 28128 6368
rect 28162 6334 28196 6368
rect 28230 6334 28264 6368
rect 28298 6334 28332 6368
rect 28366 6334 28400 6368
rect 28434 6334 28468 6368
rect 28502 6334 28536 6368
rect 28570 6334 28604 6368
rect 28638 6334 28672 6368
rect 28706 6334 28740 6368
rect 28774 6334 28808 6368
rect 28842 6334 28876 6368
rect 28910 6334 28944 6368
rect 28978 6334 29012 6368
rect 29046 6334 29080 6368
rect 29114 6334 29148 6368
rect 29182 6334 29216 6368
rect 29250 6334 29284 6368
rect 29318 6334 29352 6368
rect 29386 6334 29420 6368
rect 29454 6334 29488 6368
rect 29522 6334 29556 6368
rect 29590 6334 29624 6368
rect 29658 6334 29692 6368
rect 27330 6257 27364 6291
rect 27330 6189 27364 6223
rect 27330 6121 27364 6155
rect 27330 6053 27364 6087
rect 27330 5985 27364 6019
rect 27330 5917 27364 5951
rect 27330 5849 27364 5883
rect 27330 5781 27364 5815
rect 27330 5713 27364 5747
rect 27330 5645 27364 5679
rect 27330 5577 27364 5611
rect 27330 5509 27364 5543
rect 27330 5441 27364 5475
rect 27330 5373 27364 5407
rect 27330 5305 27364 5339
rect 27330 5237 27364 5271
rect 27330 5169 27364 5203
rect 27330 5101 27364 5135
rect 27330 5033 27364 5067
rect 27330 4965 27364 4999
rect 27330 4897 27364 4931
rect 27330 4829 27364 4863
rect 27330 4761 27364 4795
rect 27330 4693 27364 4727
rect 27330 4625 27364 4659
rect 27330 4557 27364 4591
rect 27330 4489 27364 4523
rect 27330 4421 27364 4455
rect 27330 4353 27364 4387
rect 27330 4285 27364 4319
rect 27330 4217 27364 4251
rect 27330 4149 27364 4183
rect 27330 4081 27364 4115
rect 27330 4013 27364 4047
rect 27330 3945 27364 3979
rect 27330 3877 27364 3911
rect 27330 3809 27364 3843
rect 27330 3741 27364 3775
rect 27330 3673 27364 3707
rect 27330 3605 27364 3639
rect 27330 3537 27364 3571
rect 27330 3469 27364 3503
rect 27330 3401 27364 3435
rect 27330 3333 27364 3367
rect 27330 3265 27364 3299
rect 27330 3197 27364 3231
rect 27330 3129 27364 3163
rect 27330 3061 27364 3095
rect 26524 2950 26558 2984
rect 26592 2950 26626 2984
rect 26660 2950 26694 2984
rect 26728 2950 26762 2984
rect 26796 2950 26830 2984
rect 26864 2950 26898 2984
rect 26932 2950 26966 2984
rect 27000 2950 27034 2984
rect 27068 2950 27102 2984
rect 27136 2950 27170 2984
rect 27204 2950 27238 2984
<< nsubdiffcont >>
rect 23404 15636 23438 15670
rect 23494 15636 23528 15670
rect 23584 15636 23618 15670
rect 23674 15636 23708 15670
rect 23764 15636 23798 15670
rect 23854 15636 23888 15670
rect 23944 15636 23978 15670
rect 24034 15636 24068 15670
rect 24124 15636 24158 15670
rect 23292 15579 23326 15613
rect 24182 15560 24216 15594
rect 23292 15489 23326 15523
rect 23292 15399 23326 15433
rect 23292 15309 23326 15343
rect 23292 15219 23326 15253
rect 23292 15129 23326 15163
rect 23292 15039 23326 15073
rect 23292 14949 23326 14983
rect 23292 14859 23326 14893
rect 24182 15470 24216 15504
rect 24182 15380 24216 15414
rect 24182 15290 24216 15324
rect 24182 15200 24216 15234
rect 24182 15110 24216 15144
rect 24182 15020 24216 15054
rect 24182 14930 24216 14964
rect 24182 14840 24216 14874
rect 23370 14746 23404 14780
rect 23460 14746 23494 14780
rect 23550 14746 23584 14780
rect 23640 14746 23674 14780
rect 23730 14746 23764 14780
rect 23820 14746 23854 14780
rect 23910 14746 23944 14780
rect 24000 14746 24034 14780
rect 24090 14746 24124 14780
rect 13076 11118 13110 11152
rect 13166 11118 13200 11152
rect 13256 11118 13290 11152
rect 13346 11118 13380 11152
rect 13436 11118 13470 11152
rect 13526 11118 13560 11152
rect 13616 11118 13650 11152
rect 13706 11118 13740 11152
rect 13796 11118 13830 11152
rect 12964 11061 12998 11095
rect 13854 11042 13888 11076
rect 12964 10971 12998 11005
rect 12964 10881 12998 10915
rect 12964 10791 12998 10825
rect 12964 10701 12998 10735
rect 12964 10611 12998 10645
rect 12964 10521 12998 10555
rect 12964 10431 12998 10465
rect 12964 10341 12998 10375
rect 13854 10952 13888 10986
rect 13854 10862 13888 10896
rect 13854 10772 13888 10806
rect 13854 10682 13888 10716
rect 13854 10592 13888 10626
rect 13854 10502 13888 10536
rect 13854 10412 13888 10446
rect 13854 10322 13888 10356
rect 13042 10228 13076 10262
rect 13132 10228 13166 10262
rect 13222 10228 13256 10262
rect 13312 10228 13346 10262
rect 13402 10228 13436 10262
rect 13492 10228 13526 10262
rect 13582 10228 13616 10262
rect 13672 10228 13706 10262
rect 13762 10228 13796 10262
rect 13076 9628 13110 9662
rect 13166 9628 13200 9662
rect 13256 9628 13290 9662
rect 13346 9628 13380 9662
rect 13436 9628 13470 9662
rect 13526 9628 13560 9662
rect 13616 9628 13650 9662
rect 13706 9628 13740 9662
rect 13796 9628 13830 9662
rect 12964 9571 12998 9605
rect 13854 9552 13888 9586
rect 12964 9481 12998 9515
rect 12964 9391 12998 9425
rect 12964 9301 12998 9335
rect 12964 9211 12998 9245
rect 12964 9121 12998 9155
rect 12964 9031 12998 9065
rect 12964 8941 12998 8975
rect 12964 8851 12998 8885
rect 13854 9462 13888 9496
rect 13854 9372 13888 9406
rect 13854 9282 13888 9316
rect 13854 9192 13888 9226
rect 13854 9102 13888 9136
rect 13854 9012 13888 9046
rect 13854 8922 13888 8956
rect 13854 8832 13888 8866
rect 13042 8738 13076 8772
rect 13132 8738 13166 8772
rect 13222 8738 13256 8772
rect 13312 8738 13346 8772
rect 13402 8738 13436 8772
rect 13492 8738 13526 8772
rect 13582 8738 13616 8772
rect 13672 8738 13706 8772
rect 13762 8738 13796 8772
rect 13066 8218 13100 8252
rect 13156 8218 13190 8252
rect 13246 8218 13280 8252
rect 13336 8218 13370 8252
rect 13426 8218 13460 8252
rect 13516 8218 13550 8252
rect 13606 8218 13640 8252
rect 13696 8218 13730 8252
rect 13786 8218 13820 8252
rect 12954 8161 12988 8195
rect 13844 8142 13878 8176
rect 12954 8071 12988 8105
rect 12954 7981 12988 8015
rect 12954 7891 12988 7925
rect 12954 7801 12988 7835
rect 12954 7711 12988 7745
rect 12954 7621 12988 7655
rect 12954 7531 12988 7565
rect 12954 7441 12988 7475
rect 13844 8052 13878 8086
rect 13844 7962 13878 7996
rect 13844 7872 13878 7906
rect 13844 7782 13878 7816
rect 13844 7692 13878 7726
rect 13844 7602 13878 7636
rect 13844 7512 13878 7546
rect 13844 7422 13878 7456
rect 13032 7328 13066 7362
rect 13122 7328 13156 7362
rect 13212 7328 13246 7362
rect 13302 7328 13336 7362
rect 13392 7328 13426 7362
rect 13482 7328 13516 7362
rect 13572 7328 13606 7362
rect 13662 7328 13696 7362
rect 13752 7328 13786 7362
rect 13066 6868 13100 6902
rect 13156 6868 13190 6902
rect 13246 6868 13280 6902
rect 13336 6868 13370 6902
rect 13426 6868 13460 6902
rect 13516 6868 13550 6902
rect 13606 6868 13640 6902
rect 13696 6868 13730 6902
rect 13786 6868 13820 6902
rect 12954 6811 12988 6845
rect 13844 6792 13878 6826
rect 12954 6721 12988 6755
rect 12954 6631 12988 6665
rect 12954 6541 12988 6575
rect 12954 6451 12988 6485
rect 12954 6361 12988 6395
rect 12954 6271 12988 6305
rect 12954 6181 12988 6215
rect 12954 6091 12988 6125
rect 13844 6702 13878 6736
rect 13844 6612 13878 6646
rect 13844 6522 13878 6556
rect 13844 6432 13878 6466
rect 13844 6342 13878 6376
rect 13844 6252 13878 6286
rect 13844 6162 13878 6196
rect 13844 6072 13878 6106
rect 13032 5978 13066 6012
rect 13122 5978 13156 6012
rect 13212 5978 13246 6012
rect 13302 5978 13336 6012
rect 13392 5978 13426 6012
rect 13482 5978 13516 6012
rect 13572 5978 13606 6012
rect 13662 5978 13696 6012
rect 13752 5978 13786 6012
rect 14716 6898 14750 6932
rect 14806 6898 14840 6932
rect 14896 6898 14930 6932
rect 14986 6898 15020 6932
rect 15076 6898 15110 6932
rect 15166 6898 15200 6932
rect 15256 6898 15290 6932
rect 15346 6898 15380 6932
rect 15436 6898 15470 6932
rect 14604 6841 14638 6875
rect 15494 6822 15528 6856
rect 14604 6751 14638 6785
rect 14604 6661 14638 6695
rect 14604 6571 14638 6605
rect 14604 6481 14638 6515
rect 14604 6391 14638 6425
rect 14604 6301 14638 6335
rect 14604 6211 14638 6245
rect 14604 6121 14638 6155
rect 15494 6732 15528 6766
rect 15494 6642 15528 6676
rect 15494 6552 15528 6586
rect 15494 6462 15528 6496
rect 15494 6372 15528 6406
rect 15494 6282 15528 6316
rect 15494 6192 15528 6226
rect 15494 6102 15528 6136
rect 14682 6008 14716 6042
rect 14772 6008 14806 6042
rect 14862 6008 14896 6042
rect 14952 6008 14986 6042
rect 15042 6008 15076 6042
rect 15132 6008 15166 6042
rect 15222 6008 15256 6042
rect 15312 6008 15346 6042
rect 15402 6008 15436 6042
rect 13066 5518 13100 5552
rect 13156 5518 13190 5552
rect 13246 5518 13280 5552
rect 13336 5518 13370 5552
rect 13426 5518 13460 5552
rect 13516 5518 13550 5552
rect 13606 5518 13640 5552
rect 13696 5518 13730 5552
rect 13786 5518 13820 5552
rect 12954 5461 12988 5495
rect 13844 5442 13878 5476
rect 12954 5371 12988 5405
rect 12954 5281 12988 5315
rect 12954 5191 12988 5225
rect 12954 5101 12988 5135
rect 12954 5011 12988 5045
rect 12954 4921 12988 4955
rect 12954 4831 12988 4865
rect 12954 4741 12988 4775
rect 13844 5352 13878 5386
rect 13844 5262 13878 5296
rect 13844 5172 13878 5206
rect 13844 5082 13878 5116
rect 13844 4992 13878 5026
rect 13844 4902 13878 4936
rect 13844 4812 13878 4846
rect 13844 4722 13878 4756
rect 13032 4628 13066 4662
rect 13122 4628 13156 4662
rect 13212 4628 13246 4662
rect 13302 4628 13336 4662
rect 13392 4628 13426 4662
rect 13482 4628 13516 4662
rect 13572 4628 13606 4662
rect 13662 4628 13696 4662
rect 13752 4628 13786 4662
rect 14716 5538 14750 5572
rect 14806 5538 14840 5572
rect 14896 5538 14930 5572
rect 14986 5538 15020 5572
rect 15076 5538 15110 5572
rect 15166 5538 15200 5572
rect 15256 5538 15290 5572
rect 15346 5538 15380 5572
rect 15436 5538 15470 5572
rect 14604 5481 14638 5515
rect 15494 5462 15528 5496
rect 14604 5391 14638 5425
rect 14604 5301 14638 5335
rect 14604 5211 14638 5245
rect 14604 5121 14638 5155
rect 14604 5031 14638 5065
rect 14604 4941 14638 4975
rect 14604 4851 14638 4885
rect 14604 4761 14638 4795
rect 15494 5372 15528 5406
rect 15494 5282 15528 5316
rect 15494 5192 15528 5226
rect 15494 5102 15528 5136
rect 15494 5012 15528 5046
rect 15494 4922 15528 4956
rect 15494 4832 15528 4866
rect 15494 4742 15528 4776
rect 14682 4648 14716 4682
rect 14772 4648 14806 4682
rect 14862 4648 14896 4682
rect 14952 4648 14986 4682
rect 15042 4648 15076 4682
rect 15132 4648 15166 4682
rect 15222 4648 15256 4682
rect 15312 4648 15346 4682
rect 15402 4648 15436 4682
<< mvpsubdiffcont >>
rect 23135 17312 23169 17346
rect 23203 17312 23237 17346
rect 23271 17312 23305 17346
rect 23339 17312 23373 17346
rect 23407 17312 23441 17346
rect 23475 17312 23509 17346
rect 23543 17312 23577 17346
rect 23611 17312 23645 17346
rect 23679 17312 23713 17346
rect 23747 17312 23781 17346
rect 23815 17312 23849 17346
rect 23883 17312 23917 17346
rect 23951 17312 23985 17346
rect 24019 17312 24053 17346
rect 24087 17312 24121 17346
rect 24155 17312 24189 17346
rect 24223 17312 24257 17346
rect 23016 17197 23050 17231
rect 23016 17129 23050 17163
rect 24342 17197 24376 17231
rect 23016 17061 23050 17095
rect 23016 16993 23050 17027
rect 23016 16925 23050 16959
rect 23016 16857 23050 16891
rect 23016 16789 23050 16823
rect 23016 16721 23050 16755
rect 23016 16653 23050 16687
rect 23016 16585 23050 16619
rect 23016 16517 23050 16551
rect 23016 16449 23050 16483
rect 23016 16381 23050 16415
rect 23016 16313 23050 16347
rect 23016 16245 23050 16279
rect 23016 16177 23050 16211
rect 23016 16109 23050 16143
rect 24342 17129 24376 17163
rect 24342 17061 24376 17095
rect 24342 16993 24376 17027
rect 24342 16925 24376 16959
rect 24342 16857 24376 16891
rect 24342 16789 24376 16823
rect 24342 16721 24376 16755
rect 24342 16653 24376 16687
rect 24342 16585 24376 16619
rect 24342 16517 24376 16551
rect 24342 16449 24376 16483
rect 24342 16381 24376 16415
rect 24342 16313 24376 16347
rect 24342 16245 24376 16279
rect 24342 16177 24376 16211
rect 23016 16041 23050 16075
rect 24342 16109 24376 16143
rect 24342 16041 24376 16075
rect 23135 15926 23169 15960
rect 23203 15926 23237 15960
rect 23271 15926 23305 15960
rect 23339 15926 23373 15960
rect 23407 15926 23441 15960
rect 23475 15926 23509 15960
rect 23543 15926 23577 15960
rect 23611 15926 23645 15960
rect 23679 15926 23713 15960
rect 23747 15926 23781 15960
rect 23815 15926 23849 15960
rect 23883 15926 23917 15960
rect 23951 15926 23985 15960
rect 24019 15926 24053 15960
rect 24087 15926 24121 15960
rect 24155 15926 24189 15960
rect 24223 15926 24257 15960
rect -8832 11531 -8798 11565
rect -8764 11531 -8730 11565
rect -8696 11531 -8662 11565
rect -8628 11531 -8594 11565
rect -8560 11531 -8526 11565
rect -8492 11531 -8458 11565
rect -8424 11531 -8390 11565
rect -8356 11531 -8322 11565
rect -8288 11531 -8254 11565
rect -8220 11531 -8186 11565
rect -8152 11531 -8118 11565
rect -8084 11531 -8050 11565
rect -8016 11531 -7982 11565
rect -7948 11531 -7914 11565
rect -7880 11531 -7846 11565
rect -7812 11531 -7778 11565
rect -7744 11531 -7710 11565
rect -7676 11531 -7642 11565
rect -7608 11531 -7574 11565
rect -7540 11531 -7506 11565
rect -7472 11531 -7438 11565
rect -7404 11531 -7370 11565
rect -7336 11531 -7302 11565
rect -7268 11531 -7234 11565
rect -7200 11531 -7166 11565
rect -7132 11531 -7098 11565
rect -7064 11531 -7030 11565
rect -6996 11531 -6962 11565
rect -6928 11531 -6894 11565
rect -6860 11531 -6826 11565
rect -6792 11531 -6758 11565
rect -6724 11531 -6690 11565
rect -6656 11531 -6622 11565
rect -6588 11531 -6554 11565
rect -6520 11531 -6486 11565
rect -6452 11531 -6418 11565
rect -6384 11531 -6350 11565
rect -6316 11531 -6282 11565
rect -6248 11531 -6214 11565
rect -6180 11531 -6146 11565
rect -6112 11531 -6078 11565
rect -6044 11531 -6010 11565
rect -5976 11531 -5942 11565
rect -5908 11531 -5874 11565
rect -5840 11531 -5806 11565
rect -5772 11531 -5738 11565
rect -5704 11531 -5670 11565
rect -5636 11531 -5602 11565
rect -5568 11531 -5534 11565
rect -5500 11531 -5466 11565
rect -5432 11531 -5398 11565
rect -5364 11531 -5330 11565
rect -5296 11531 -5262 11565
rect -5228 11531 -5194 11565
rect -5160 11531 -5126 11565
rect -5092 11531 -5058 11565
rect -5024 11531 -4990 11565
rect -4956 11531 -4922 11565
rect -4888 11531 -4854 11565
rect -4820 11531 -4786 11565
rect -4752 11531 -4718 11565
rect -4684 11531 -4650 11565
rect -4616 11531 -4582 11565
rect -4548 11531 -4514 11565
rect -4480 11531 -4446 11565
rect -4412 11531 -4378 11565
rect -4344 11531 -4310 11565
rect -4276 11531 -4242 11565
rect -4208 11531 -4174 11565
rect -4140 11531 -4106 11565
rect -4072 11531 -4038 11565
rect -4004 11531 -3970 11565
rect -3936 11531 -3902 11565
rect -3868 11531 -3834 11565
rect -3800 11531 -3766 11565
rect -3732 11531 -3698 11565
rect -3664 11531 -3630 11565
rect -3596 11531 -3562 11565
rect -9081 11341 -9047 11375
rect -9081 11273 -9047 11307
rect -3355 11301 -3321 11335
rect -9081 11205 -9047 11239
rect -9081 11137 -9047 11171
rect -3355 11233 -3321 11267
rect -3355 11165 -3321 11199
rect -9081 11069 -9047 11103
rect -9081 11001 -9047 11035
rect -9081 10933 -9047 10967
rect -9081 10865 -9047 10899
rect -9081 10797 -9047 10831
rect -9081 10729 -9047 10763
rect -9081 10661 -9047 10695
rect -9081 10593 -9047 10627
rect -9081 10525 -9047 10559
rect -9081 10457 -9047 10491
rect -9081 10389 -9047 10423
rect -9081 10321 -9047 10355
rect -9081 10253 -9047 10287
rect -9081 10185 -9047 10219
rect -3355 11097 -3321 11131
rect -3355 11029 -3321 11063
rect -3355 10961 -3321 10995
rect -3355 10893 -3321 10927
rect -3355 10825 -3321 10859
rect -3355 10757 -3321 10791
rect -3355 10689 -3321 10723
rect -3355 10621 -3321 10655
rect -3355 10553 -3321 10587
rect -3355 10485 -3321 10519
rect -3355 10417 -3321 10451
rect -3355 10349 -3321 10383
rect -3355 10281 -3321 10315
rect -3355 10213 -3321 10247
rect -9081 10117 -9047 10151
rect -9081 10049 -9047 10083
rect -3355 10145 -3321 10179
rect -3355 10077 -3321 10111
rect -9081 9981 -9047 10015
rect -9081 9913 -9047 9947
rect -3355 10009 -3321 10043
rect -3355 9941 -3321 9975
rect -9081 9845 -9047 9879
rect -9081 9777 -9047 9811
rect -3355 9873 -3321 9907
rect -3355 9805 -3321 9839
rect -9081 9709 -9047 9743
rect -9081 9641 -9047 9675
rect -9081 9573 -9047 9607
rect -9081 9505 -9047 9539
rect -9081 9437 -9047 9471
rect -9081 9369 -9047 9403
rect -9081 9301 -9047 9335
rect -9081 9233 -9047 9267
rect -9081 9165 -9047 9199
rect -9081 9097 -9047 9131
rect -9081 9029 -9047 9063
rect -9081 8961 -9047 8995
rect -9081 8893 -9047 8927
rect -9081 8825 -9047 8859
rect -3355 9737 -3321 9771
rect -3355 9669 -3321 9703
rect -3355 9601 -3321 9635
rect -3355 9533 -3321 9567
rect -3355 9465 -3321 9499
rect -3355 9397 -3321 9431
rect -3355 9329 -3321 9363
rect -3355 9261 -3321 9295
rect -3355 9193 -3321 9227
rect -3355 9125 -3321 9159
rect -3355 9057 -3321 9091
rect -3355 8989 -3321 9023
rect -3355 8921 -3321 8955
rect -3355 8853 -3321 8887
rect -9081 8757 -9047 8791
rect -9081 8689 -9047 8723
rect -3355 8785 -3321 8819
rect -3355 8717 -3321 8751
rect -9081 8621 -9047 8655
rect -3355 8649 -3321 8683
rect -3355 8581 -3321 8615
rect -8813 8365 -8779 8399
rect -8745 8365 -8711 8399
rect -8677 8365 -8643 8399
rect -8609 8365 -8575 8399
rect -8541 8365 -8507 8399
rect -8473 8365 -8439 8399
rect -8405 8365 -8371 8399
rect -8337 8365 -8303 8399
rect -8269 8365 -8235 8399
rect -8201 8365 -8167 8399
rect -8133 8365 -8099 8399
rect -8065 8365 -8031 8399
rect -7997 8365 -7963 8399
rect -7929 8365 -7895 8399
rect -7861 8365 -7827 8399
rect -7793 8365 -7759 8399
rect -7725 8365 -7691 8399
rect -7657 8365 -7623 8399
rect -7589 8365 -7555 8399
rect -7521 8365 -7487 8399
rect -7453 8365 -7419 8399
rect -7385 8365 -7351 8399
rect -7317 8365 -7283 8399
rect -7249 8365 -7215 8399
rect -7181 8365 -7147 8399
rect -7113 8365 -7079 8399
rect -7045 8365 -7011 8399
rect -6977 8365 -6943 8399
rect -6909 8365 -6875 8399
rect -6841 8365 -6807 8399
rect -6773 8365 -6739 8399
rect -6705 8365 -6671 8399
rect -6637 8365 -6603 8399
rect -6569 8365 -6535 8399
rect -6501 8365 -6467 8399
rect -6433 8365 -6399 8399
rect -6365 8365 -6331 8399
rect -6297 8365 -6263 8399
rect -6229 8365 -6195 8399
rect -6161 8365 -6127 8399
rect -6093 8365 -6059 8399
rect -6025 8365 -5991 8399
rect -5957 8365 -5923 8399
rect -5889 8365 -5855 8399
rect -5821 8365 -5787 8399
rect -5753 8365 -5719 8399
rect -5685 8365 -5651 8399
rect -5617 8365 -5583 8399
rect -5549 8365 -5515 8399
rect -5481 8365 -5447 8399
rect -5413 8365 -5379 8399
rect -5345 8365 -5311 8399
rect -5277 8365 -5243 8399
rect -5209 8365 -5175 8399
rect -5141 8365 -5107 8399
rect -5073 8365 -5039 8399
rect -5005 8365 -4971 8399
rect -4937 8365 -4903 8399
rect -4869 8365 -4835 8399
rect -4801 8365 -4767 8399
rect -4733 8365 -4699 8399
rect -4665 8365 -4631 8399
rect -4597 8365 -4563 8399
rect -4529 8365 -4495 8399
rect -4461 8365 -4427 8399
rect -4393 8365 -4359 8399
rect -4325 8365 -4291 8399
rect -4257 8365 -4223 8399
rect -4189 8365 -4155 8399
rect -4121 8365 -4087 8399
rect -4053 8365 -4019 8399
rect -3985 8365 -3951 8399
rect -3917 8365 -3883 8399
rect -3849 8365 -3815 8399
rect -3781 8365 -3747 8399
rect -3713 8365 -3679 8399
rect -3645 8365 -3611 8399
rect -3577 8365 -3543 8399
rect -7749 7825 -7715 7859
rect -7681 7825 -7647 7859
rect -7613 7825 -7579 7859
rect -7545 7825 -7511 7859
rect -7477 7825 -7443 7859
rect -7409 7825 -7375 7859
rect -7341 7825 -7307 7859
rect -7273 7825 -7239 7859
rect -7205 7825 -7171 7859
rect -7137 7825 -7103 7859
rect -7069 7825 -7035 7859
rect -7001 7825 -6967 7859
rect -6933 7825 -6899 7859
rect -6865 7825 -6831 7859
rect -6797 7825 -6763 7859
rect -6729 7825 -6695 7859
rect -6661 7825 -6627 7859
rect -6593 7825 -6559 7859
rect -6525 7825 -6491 7859
rect -6457 7825 -6423 7859
rect -6389 7825 -6355 7859
rect -6321 7825 -6287 7859
rect -6253 7825 -6219 7859
rect -6185 7825 -6151 7859
rect -6117 7825 -6083 7859
rect -6049 7825 -6015 7859
rect -5981 7825 -5947 7859
rect -5913 7825 -5879 7859
rect -5845 7825 -5811 7859
rect -5777 7825 -5743 7859
rect -5709 7825 -5675 7859
rect -5641 7825 -5607 7859
rect -5573 7825 -5539 7859
rect -5505 7825 -5471 7859
rect -5437 7825 -5403 7859
rect -5369 7825 -5335 7859
rect -5301 7825 -5267 7859
rect -5233 7825 -5199 7859
rect -5165 7825 -5131 7859
rect -5097 7825 -5063 7859
rect -5029 7825 -4995 7859
rect -4961 7825 -4927 7859
rect -4893 7825 -4859 7859
rect -4825 7825 -4791 7859
rect -4757 7825 -4723 7859
rect -4689 7825 -4655 7859
rect -4621 7825 -4587 7859
rect -4553 7825 -4519 7859
rect -4485 7825 -4451 7859
rect -4417 7825 -4383 7859
rect -4349 7825 -4315 7859
rect -4281 7825 -4247 7859
rect -4213 7825 -4179 7859
rect -4145 7825 -4111 7859
rect -4077 7825 -4043 7859
rect -4009 7825 -3975 7859
rect -3941 7825 -3907 7859
rect -3873 7825 -3839 7859
rect -3805 7825 -3771 7859
rect -3737 7825 -3703 7859
rect -3669 7825 -3635 7859
rect -3601 7825 -3567 7859
rect -7968 7648 -7934 7682
rect -3456 7660 -3422 7694
rect -7968 7580 -7934 7614
rect -7968 7512 -7934 7546
rect -3456 7592 -3422 7626
rect -7968 7444 -7934 7478
rect -7968 7376 -7934 7410
rect -7968 7308 -7934 7342
rect -7968 7240 -7934 7274
rect -7968 7172 -7934 7206
rect -7968 7104 -7934 7138
rect -7968 7036 -7934 7070
rect -7968 6968 -7934 7002
rect -7968 6900 -7934 6934
rect -7968 6832 -7934 6866
rect -7968 6764 -7934 6798
rect -7968 6696 -7934 6730
rect -7968 6628 -7934 6662
rect -7968 6560 -7934 6594
rect -7968 6492 -7934 6526
rect -7968 6424 -7934 6458
rect -7968 6356 -7934 6390
rect -7968 6288 -7934 6322
rect -7968 6220 -7934 6254
rect -7968 6152 -7934 6186
rect -7968 6084 -7934 6118
rect -7968 6016 -7934 6050
rect -7968 5948 -7934 5982
rect -7968 5880 -7934 5914
rect -7968 5812 -7934 5846
rect -7968 5744 -7934 5778
rect -7968 5676 -7934 5710
rect -7968 5608 -7934 5642
rect -7968 5540 -7934 5574
rect -3456 7524 -3422 7558
rect -3456 7456 -3422 7490
rect -3456 7388 -3422 7422
rect -3456 7320 -3422 7354
rect -3456 7252 -3422 7286
rect -3456 7184 -3422 7218
rect -3456 7116 -3422 7150
rect 17419 7724 17453 7758
rect 17487 7724 17521 7758
rect 17555 7724 17589 7758
rect 17623 7724 17657 7758
rect 17691 7724 17725 7758
rect 17759 7724 17793 7758
rect 17827 7724 17861 7758
rect 17895 7724 17929 7758
rect 17963 7724 17997 7758
rect 18031 7724 18065 7758
rect 18099 7724 18133 7758
rect 18167 7724 18201 7758
rect 18235 7724 18269 7758
rect 18303 7724 18337 7758
rect 18371 7724 18405 7758
rect 18439 7724 18473 7758
rect 18507 7724 18541 7758
rect 17300 7595 17334 7629
rect 17300 7527 17334 7561
rect 18626 7595 18660 7629
rect 17300 7459 17334 7493
rect 17300 7391 17334 7425
rect 17300 7323 17334 7357
rect 17300 7255 17334 7289
rect -3456 7048 -3422 7082
rect -3456 6980 -3422 7014
rect -3456 6912 -3422 6946
rect -3456 6844 -3422 6878
rect -3456 6776 -3422 6810
rect -3456 6708 -3422 6742
rect -3456 6640 -3422 6674
rect -3456 6572 -3422 6606
rect -3456 6504 -3422 6538
rect -3456 6436 -3422 6470
rect -3456 6368 -3422 6402
rect -3456 6300 -3422 6334
rect -3456 6232 -3422 6266
rect -3456 6164 -3422 6198
rect -3456 6096 -3422 6130
rect -3456 6028 -3422 6062
rect -3456 5960 -3422 5994
rect -3456 5892 -3422 5926
rect -3456 5824 -3422 5858
rect -3456 5756 -3422 5790
rect -3456 5688 -3422 5722
rect -3456 5620 -3422 5654
rect -3456 5552 -3422 5586
rect -7968 5472 -7934 5506
rect -3456 5484 -3422 5518
rect -7968 5404 -7934 5438
rect -3456 5416 -3422 5450
rect -7773 5245 -7739 5279
rect -7705 5245 -7671 5279
rect -7637 5245 -7603 5279
rect -7569 5245 -7535 5279
rect -7501 5245 -7467 5279
rect -7433 5245 -7399 5279
rect -7365 5245 -7331 5279
rect -7297 5245 -7263 5279
rect -7229 5245 -7195 5279
rect -7161 5245 -7127 5279
rect -7093 5245 -7059 5279
rect -7025 5245 -6991 5279
rect -6957 5245 -6923 5279
rect -6889 5245 -6855 5279
rect -6821 5245 -6787 5279
rect -6753 5245 -6719 5279
rect -6685 5245 -6651 5279
rect -6617 5245 -6583 5279
rect -6549 5245 -6515 5279
rect -6481 5245 -6447 5279
rect -6413 5245 -6379 5279
rect -6345 5245 -6311 5279
rect -6277 5245 -6243 5279
rect -6209 5245 -6175 5279
rect -6141 5245 -6107 5279
rect -6073 5245 -6039 5279
rect -6005 5245 -5971 5279
rect -5937 5245 -5903 5279
rect -5869 5245 -5835 5279
rect -5801 5245 -5767 5279
rect -5733 5245 -5699 5279
rect -5665 5245 -5631 5279
rect -5597 5245 -5563 5279
rect -5529 5245 -5495 5279
rect -5461 5245 -5427 5279
rect -5393 5245 -5359 5279
rect -5325 5245 -5291 5279
rect -5257 5245 -5223 5279
rect -5189 5245 -5155 5279
rect -5121 5245 -5087 5279
rect -5053 5245 -5019 5279
rect -4985 5245 -4951 5279
rect -4917 5245 -4883 5279
rect -4849 5245 -4815 5279
rect -4781 5245 -4747 5279
rect -4713 5245 -4679 5279
rect -4645 5245 -4611 5279
rect -4577 5245 -4543 5279
rect -4509 5245 -4475 5279
rect -4441 5245 -4407 5279
rect -4373 5245 -4339 5279
rect -4305 5245 -4271 5279
rect -4237 5245 -4203 5279
rect -4169 5245 -4135 5279
rect -4101 5245 -4067 5279
rect -4033 5245 -3999 5279
rect -3965 5245 -3931 5279
rect -3897 5245 -3863 5279
rect -3829 5245 -3795 5279
rect -3761 5245 -3727 5279
rect -3693 5245 -3659 5279
rect -3625 5245 -3591 5279
rect 17300 7187 17334 7221
rect 17300 7119 17334 7153
rect 17300 7051 17334 7085
rect 17300 6983 17334 7017
rect 17300 6915 17334 6949
rect 17300 6847 17334 6881
rect 17300 6779 17334 6813
rect 17300 6711 17334 6745
rect 17300 6643 17334 6677
rect 17300 6575 17334 6609
rect 17300 6507 17334 6541
rect 17300 6439 17334 6473
rect 17300 6371 17334 6405
rect 17300 6303 17334 6337
rect 17300 6235 17334 6269
rect 17300 6167 17334 6201
rect 17300 6099 17334 6133
rect 17300 6031 17334 6065
rect 17300 5963 17334 5997
rect 17300 5895 17334 5929
rect 17300 5827 17334 5861
rect 17300 5759 17334 5793
rect 17300 5691 17334 5725
rect 17300 5623 17334 5657
rect 17300 5555 17334 5589
rect 17300 5487 17334 5521
rect 17300 5419 17334 5453
rect 17300 5351 17334 5385
rect 17300 5283 17334 5317
rect 17300 5215 17334 5249
rect 17300 5147 17334 5181
rect 17300 5079 17334 5113
rect 17300 5011 17334 5045
rect 17300 4943 17334 4977
rect 17300 4875 17334 4909
rect 17300 4807 17334 4841
rect 17300 4739 17334 4773
rect 17300 4671 17334 4705
rect 17300 4603 17334 4637
rect 17300 4535 17334 4569
rect 18626 7527 18660 7561
rect 18626 7459 18660 7493
rect 18626 7391 18660 7425
rect 18626 7323 18660 7357
rect 18626 7255 18660 7289
rect 18626 7187 18660 7221
rect 18626 7119 18660 7153
rect 18626 7051 18660 7085
rect 18626 6983 18660 7017
rect 18626 6915 18660 6949
rect 18626 6847 18660 6881
rect 18626 6779 18660 6813
rect 18626 6711 18660 6745
rect 18626 6643 18660 6677
rect 18626 6575 18660 6609
rect 18626 6507 18660 6541
rect 18626 6439 18660 6473
rect 18626 6371 18660 6405
rect 18626 6303 18660 6337
rect 18626 6235 18660 6269
rect 18626 6167 18660 6201
rect 18626 6099 18660 6133
rect 18626 6031 18660 6065
rect 18626 5963 18660 5997
rect 18626 5895 18660 5929
rect 18626 5827 18660 5861
rect 18626 5759 18660 5793
rect 18626 5691 18660 5725
rect 18626 5623 18660 5657
rect 18626 5555 18660 5589
rect 18626 5487 18660 5521
rect 18626 5419 18660 5453
rect 18626 5351 18660 5385
rect 18626 5283 18660 5317
rect 18626 5215 18660 5249
rect 18626 5147 18660 5181
rect 18626 5079 18660 5113
rect 18626 5011 18660 5045
rect 18626 4943 18660 4977
rect 18626 4875 18660 4909
rect 18626 4807 18660 4841
rect 18626 4739 18660 4773
rect 18626 4671 18660 4705
rect 18626 4603 18660 4637
rect 17300 4467 17334 4501
rect 18626 4535 18660 4569
rect 18626 4467 18660 4501
rect 17419 4338 17453 4372
rect 17487 4338 17521 4372
rect 17555 4338 17589 4372
rect 17623 4338 17657 4372
rect 17691 4338 17725 4372
rect 17759 4338 17793 4372
rect 17827 4338 17861 4372
rect 17895 4338 17929 4372
rect 17963 4338 17997 4372
rect 18031 4338 18065 4372
rect 18099 4338 18133 4372
rect 18167 4338 18201 4372
rect 18235 4338 18269 4372
rect 18303 4338 18337 4372
rect 18371 4338 18405 4372
rect 18439 4338 18473 4372
rect 18507 4338 18541 4372
rect 18869 7724 18903 7758
rect 18937 7724 18971 7758
rect 19005 7724 19039 7758
rect 19073 7724 19107 7758
rect 19141 7724 19175 7758
rect 19209 7724 19243 7758
rect 19277 7724 19311 7758
rect 19345 7724 19379 7758
rect 19413 7724 19447 7758
rect 19481 7724 19515 7758
rect 19549 7724 19583 7758
rect 19617 7724 19651 7758
rect 19685 7724 19719 7758
rect 19753 7724 19787 7758
rect 19821 7724 19855 7758
rect 19889 7724 19923 7758
rect 19957 7724 19991 7758
rect 18750 7595 18784 7629
rect 18750 7527 18784 7561
rect 20076 7595 20110 7629
rect 18750 7459 18784 7493
rect 18750 7391 18784 7425
rect 18750 7323 18784 7357
rect 18750 7255 18784 7289
rect 18750 7187 18784 7221
rect 18750 7119 18784 7153
rect 18750 7051 18784 7085
rect 18750 6983 18784 7017
rect 18750 6915 18784 6949
rect 18750 6847 18784 6881
rect 18750 6779 18784 6813
rect 18750 6711 18784 6745
rect 18750 6643 18784 6677
rect 18750 6575 18784 6609
rect 18750 6507 18784 6541
rect 18750 6439 18784 6473
rect 18750 6371 18784 6405
rect 18750 6303 18784 6337
rect 18750 6235 18784 6269
rect 18750 6167 18784 6201
rect 18750 6099 18784 6133
rect 18750 6031 18784 6065
rect 18750 5963 18784 5997
rect 18750 5895 18784 5929
rect 18750 5827 18784 5861
rect 18750 5759 18784 5793
rect 18750 5691 18784 5725
rect 18750 5623 18784 5657
rect 18750 5555 18784 5589
rect 18750 5487 18784 5521
rect 18750 5419 18784 5453
rect 18750 5351 18784 5385
rect 18750 5283 18784 5317
rect 18750 5215 18784 5249
rect 18750 5147 18784 5181
rect 18750 5079 18784 5113
rect 18750 5011 18784 5045
rect 18750 4943 18784 4977
rect 18750 4875 18784 4909
rect 18750 4807 18784 4841
rect 18750 4739 18784 4773
rect 18750 4671 18784 4705
rect 18750 4603 18784 4637
rect 18750 4535 18784 4569
rect 20076 7527 20110 7561
rect 20076 7459 20110 7493
rect 20076 7391 20110 7425
rect 20076 7323 20110 7357
rect 20076 7255 20110 7289
rect 20076 7187 20110 7221
rect 20076 7119 20110 7153
rect 20076 7051 20110 7085
rect 20076 6983 20110 7017
rect 20076 6915 20110 6949
rect 20076 6847 20110 6881
rect 20076 6779 20110 6813
rect 20076 6711 20110 6745
rect 20076 6643 20110 6677
rect 20076 6575 20110 6609
rect 20076 6507 20110 6541
rect 20076 6439 20110 6473
rect 20076 6371 20110 6405
rect 20076 6303 20110 6337
rect 20076 6235 20110 6269
rect 20076 6167 20110 6201
rect 20076 6099 20110 6133
rect 20076 6031 20110 6065
rect 20076 5963 20110 5997
rect 20076 5895 20110 5929
rect 20076 5827 20110 5861
rect 20076 5759 20110 5793
rect 20076 5691 20110 5725
rect 20076 5623 20110 5657
rect 20076 5555 20110 5589
rect 20076 5487 20110 5521
rect 20076 5419 20110 5453
rect 20076 5351 20110 5385
rect 20076 5283 20110 5317
rect 20076 5215 20110 5249
rect 20076 5147 20110 5181
rect 20076 5079 20110 5113
rect 20076 5011 20110 5045
rect 20076 4943 20110 4977
rect 20076 4875 20110 4909
rect 20076 4807 20110 4841
rect 20076 4739 20110 4773
rect 20076 4671 20110 4705
rect 20076 4603 20110 4637
rect 23035 11916 23069 11950
rect 23103 11916 23137 11950
rect 23171 11916 23205 11950
rect 23239 11916 23273 11950
rect 23307 11916 23341 11950
rect 23375 11916 23409 11950
rect 23443 11916 23477 11950
rect 23511 11916 23545 11950
rect 23579 11916 23613 11950
rect 23647 11916 23681 11950
rect 23715 11916 23749 11950
rect 23783 11916 23817 11950
rect 23851 11916 23885 11950
rect 23919 11916 23953 11950
rect 23987 11916 24021 11950
rect 24055 11916 24089 11950
rect 24123 11916 24157 11950
rect 24191 11916 24225 11950
rect 22920 11797 22954 11831
rect 24306 11797 24340 11831
rect 22920 11729 22954 11763
rect 22920 11661 22954 11695
rect 22920 11593 22954 11627
rect 22920 11525 22954 11559
rect 22920 11457 22954 11491
rect 22920 11389 22954 11423
rect 22920 11321 22954 11355
rect 22920 11253 22954 11287
rect 22920 11185 22954 11219
rect 22920 11117 22954 11151
rect 22920 11049 22954 11083
rect 22920 10981 22954 11015
rect 22920 10913 22954 10947
rect 22920 10845 22954 10879
rect 22920 10777 22954 10811
rect 24306 11729 24340 11763
rect 24306 11661 24340 11695
rect 24306 11593 24340 11627
rect 24306 11525 24340 11559
rect 24306 11457 24340 11491
rect 24306 11389 24340 11423
rect 24306 11321 24340 11355
rect 24306 11253 24340 11287
rect 24306 11185 24340 11219
rect 24306 11117 24340 11151
rect 24306 11049 24340 11083
rect 24306 10981 24340 11015
rect 24306 10913 24340 10947
rect 24306 10845 24340 10879
rect 24306 10777 24340 10811
rect 22920 10709 22954 10743
rect 24306 10709 24340 10743
rect 23035 10590 23069 10624
rect 23103 10590 23137 10624
rect 23171 10590 23205 10624
rect 23239 10590 23273 10624
rect 23307 10590 23341 10624
rect 23375 10590 23409 10624
rect 23443 10590 23477 10624
rect 23511 10590 23545 10624
rect 23579 10590 23613 10624
rect 23647 10590 23681 10624
rect 23715 10590 23749 10624
rect 23783 10590 23817 10624
rect 23851 10590 23885 10624
rect 23919 10590 23953 10624
rect 23987 10590 24021 10624
rect 24055 10590 24089 10624
rect 24123 10590 24157 10624
rect 24191 10590 24225 10624
rect 23515 7980 23549 8014
rect 23583 7980 23617 8014
rect 23651 7980 23685 8014
rect 23719 7980 23753 8014
rect 23787 7980 23821 8014
rect 23855 7980 23889 8014
rect 23923 7980 23957 8014
rect 23991 7980 24025 8014
rect 24059 7980 24093 8014
rect 24127 7980 24161 8014
rect 24195 7980 24229 8014
rect 24263 7980 24297 8014
rect 24331 7980 24365 8014
rect 24399 7980 24433 8014
rect 24467 7980 24501 8014
rect 24535 7980 24569 8014
rect 24603 7980 24637 8014
rect 24671 7980 24705 8014
rect 23400 7872 23434 7906
rect 23400 7804 23434 7838
rect 24786 7872 24820 7906
rect 23400 7736 23434 7770
rect 23400 7668 23434 7702
rect 23400 7600 23434 7634
rect 23400 7532 23434 7566
rect 23400 7464 23434 7498
rect 23400 7396 23434 7430
rect 23400 7328 23434 7362
rect 23400 7260 23434 7294
rect 23400 7192 23434 7226
rect 23400 7124 23434 7158
rect 23400 7056 23434 7090
rect 23400 6988 23434 7022
rect 23400 6920 23434 6954
rect 23400 6852 23434 6886
rect 24786 7804 24820 7838
rect 24786 7736 24820 7770
rect 24786 7668 24820 7702
rect 24786 7600 24820 7634
rect 24786 7532 24820 7566
rect 24786 7464 24820 7498
rect 24786 7396 24820 7430
rect 24786 7328 24820 7362
rect 24786 7260 24820 7294
rect 24786 7192 24820 7226
rect 24786 7124 24820 7158
rect 24786 7056 24820 7090
rect 24786 6988 24820 7022
rect 24786 6920 24820 6954
rect 24786 6852 24820 6886
rect 23400 6784 23434 6818
rect 24786 6784 24820 6818
rect 23400 6716 23434 6750
rect 23400 6648 23434 6682
rect 23400 6580 23434 6614
rect 23400 6512 23434 6546
rect 23400 6444 23434 6478
rect 23400 6376 23434 6410
rect 23400 6308 23434 6342
rect 23400 6240 23434 6274
rect 23400 6172 23434 6206
rect 23400 6104 23434 6138
rect 23400 6036 23434 6070
rect 23400 5968 23434 6002
rect 23400 5900 23434 5934
rect 23400 5832 23434 5866
rect 23400 5764 23434 5798
rect 24786 6716 24820 6750
rect 24786 6648 24820 6682
rect 24786 6580 24820 6614
rect 24786 6512 24820 6546
rect 24786 6444 24820 6478
rect 24786 6376 24820 6410
rect 24786 6308 24820 6342
rect 24786 6240 24820 6274
rect 24786 6172 24820 6206
rect 24786 6104 24820 6138
rect 24786 6036 24820 6070
rect 24786 5968 24820 6002
rect 24786 5900 24820 5934
rect 24786 5832 24820 5866
rect 23400 5696 23434 5730
rect 24786 5764 24820 5798
rect 23400 5628 23434 5662
rect 23400 5560 23434 5594
rect 23400 5492 23434 5526
rect 23400 5424 23434 5458
rect 23400 5356 23434 5390
rect 23400 5288 23434 5322
rect 23400 5220 23434 5254
rect 23400 5152 23434 5186
rect 23400 5084 23434 5118
rect 23400 5016 23434 5050
rect 23400 4948 23434 4982
rect 23400 4880 23434 4914
rect 23400 4812 23434 4846
rect 23400 4744 23434 4778
rect 24786 5696 24820 5730
rect 24786 5628 24820 5662
rect 24786 5560 24820 5594
rect 24786 5492 24820 5526
rect 24786 5424 24820 5458
rect 24786 5356 24820 5390
rect 24786 5288 24820 5322
rect 24786 5220 24820 5254
rect 24786 5152 24820 5186
rect 24786 5084 24820 5118
rect 24786 5016 24820 5050
rect 24786 4948 24820 4982
rect 24786 4880 24820 4914
rect 24786 4812 24820 4846
rect 24786 4744 24820 4778
rect 23400 4676 23434 4710
rect 24786 4676 24820 4710
rect 23400 4608 23434 4642
rect 18750 4467 18784 4501
rect 20076 4535 20110 4569
rect 20076 4467 20110 4501
rect 18869 4338 18903 4372
rect 18937 4338 18971 4372
rect 19005 4338 19039 4372
rect 19073 4338 19107 4372
rect 19141 4338 19175 4372
rect 19209 4338 19243 4372
rect 19277 4338 19311 4372
rect 19345 4338 19379 4372
rect 19413 4338 19447 4372
rect 19481 4338 19515 4372
rect 19549 4338 19583 4372
rect 19617 4338 19651 4372
rect 19685 4338 19719 4372
rect 19753 4338 19787 4372
rect 19821 4338 19855 4372
rect 19889 4338 19923 4372
rect 19957 4338 19991 4372
rect 23400 4540 23434 4574
rect 23400 4472 23434 4506
rect 23400 4404 23434 4438
rect 23400 4336 23434 4370
rect 23400 4268 23434 4302
rect 23400 4200 23434 4234
rect 23400 4132 23434 4166
rect 23400 4064 23434 4098
rect 23400 3996 23434 4030
rect 23400 3928 23434 3962
rect 23400 3860 23434 3894
rect 23400 3792 23434 3826
rect 23400 3724 23434 3758
rect 23400 3656 23434 3690
rect 24786 4608 24820 4642
rect 24786 4540 24820 4574
rect 24786 4472 24820 4506
rect 24786 4404 24820 4438
rect 24786 4336 24820 4370
rect 24786 4268 24820 4302
rect 24786 4200 24820 4234
rect 24786 4132 24820 4166
rect 24786 4064 24820 4098
rect 24786 3996 24820 4030
rect 24786 3928 24820 3962
rect 24786 3860 24820 3894
rect 24786 3792 24820 3826
rect 24786 3724 24820 3758
rect 23400 3588 23434 3622
rect 24786 3656 24820 3690
rect 24786 3588 24820 3622
rect 23515 3480 23549 3514
rect 23583 3480 23617 3514
rect 23651 3480 23685 3514
rect 23719 3480 23753 3514
rect 23787 3480 23821 3514
rect 23855 3480 23889 3514
rect 23923 3480 23957 3514
rect 23991 3480 24025 3514
rect 24059 3480 24093 3514
rect 24127 3480 24161 3514
rect 24195 3480 24229 3514
rect 24263 3480 24297 3514
rect 24331 3480 24365 3514
rect 24399 3480 24433 3514
rect 24467 3480 24501 3514
rect 24535 3480 24569 3514
rect 24603 3480 24637 3514
rect 24671 3480 24705 3514
rect 25015 7980 25049 8014
rect 25083 7980 25117 8014
rect 25151 7980 25185 8014
rect 25219 7980 25253 8014
rect 25287 7980 25321 8014
rect 25355 7980 25389 8014
rect 25423 7980 25457 8014
rect 25491 7980 25525 8014
rect 25559 7980 25593 8014
rect 25627 7980 25661 8014
rect 25695 7980 25729 8014
rect 25763 7980 25797 8014
rect 25831 7980 25865 8014
rect 25899 7980 25933 8014
rect 25967 7980 26001 8014
rect 26035 7980 26069 8014
rect 26103 7980 26137 8014
rect 26171 7980 26205 8014
rect 24900 7872 24934 7906
rect 24900 7804 24934 7838
rect 26286 7872 26320 7906
rect 24900 7736 24934 7770
rect 24900 7668 24934 7702
rect 24900 7600 24934 7634
rect 24900 7532 24934 7566
rect 24900 7464 24934 7498
rect 24900 7396 24934 7430
rect 24900 7328 24934 7362
rect 24900 7260 24934 7294
rect 24900 7192 24934 7226
rect 24900 7124 24934 7158
rect 24900 7056 24934 7090
rect 24900 6988 24934 7022
rect 24900 6920 24934 6954
rect 24900 6852 24934 6886
rect 26286 7804 26320 7838
rect 26286 7736 26320 7770
rect 26286 7668 26320 7702
rect 26286 7600 26320 7634
rect 26286 7532 26320 7566
rect 26286 7464 26320 7498
rect 26286 7396 26320 7430
rect 26286 7328 26320 7362
rect 26286 7260 26320 7294
rect 26286 7192 26320 7226
rect 26286 7124 26320 7158
rect 26286 7056 26320 7090
rect 26286 6988 26320 7022
rect 26286 6920 26320 6954
rect 26286 6852 26320 6886
rect 24900 6784 24934 6818
rect 26286 6784 26320 6818
rect 24900 6716 24934 6750
rect 24900 6648 24934 6682
rect 24900 6580 24934 6614
rect 24900 6512 24934 6546
rect 24900 6444 24934 6478
rect 24900 6376 24934 6410
rect 24900 6308 24934 6342
rect 24900 6240 24934 6274
rect 24900 6172 24934 6206
rect 24900 6104 24934 6138
rect 24900 6036 24934 6070
rect 24900 5968 24934 6002
rect 24900 5900 24934 5934
rect 24900 5832 24934 5866
rect 24900 5764 24934 5798
rect 26286 6716 26320 6750
rect 26286 6648 26320 6682
rect 26286 6580 26320 6614
rect 26286 6512 26320 6546
rect 26286 6444 26320 6478
rect 26286 6376 26320 6410
rect 26286 6308 26320 6342
rect 26286 6240 26320 6274
rect 26286 6172 26320 6206
rect 26286 6104 26320 6138
rect 26286 6036 26320 6070
rect 26286 5968 26320 6002
rect 26286 5900 26320 5934
rect 26286 5832 26320 5866
rect 24900 5696 24934 5730
rect 26286 5764 26320 5798
rect 24900 5628 24934 5662
rect 24900 5560 24934 5594
rect 24900 5492 24934 5526
rect 24900 5424 24934 5458
rect 24900 5356 24934 5390
rect 24900 5288 24934 5322
rect 24900 5220 24934 5254
rect 24900 5152 24934 5186
rect 24900 5084 24934 5118
rect 24900 5016 24934 5050
rect 24900 4948 24934 4982
rect 24900 4880 24934 4914
rect 24900 4812 24934 4846
rect 24900 4744 24934 4778
rect 26286 5696 26320 5730
rect 26286 5628 26320 5662
rect 26286 5560 26320 5594
rect 26286 5492 26320 5526
rect 26286 5424 26320 5458
rect 26286 5356 26320 5390
rect 26286 5288 26320 5322
rect 26286 5220 26320 5254
rect 26286 5152 26320 5186
rect 26286 5084 26320 5118
rect 26286 5016 26320 5050
rect 26286 4948 26320 4982
rect 26286 4880 26320 4914
rect 26286 4812 26320 4846
rect 26286 4744 26320 4778
rect 24900 4676 24934 4710
rect 26286 4676 26320 4710
rect 24900 4608 24934 4642
rect 24900 4540 24934 4574
rect 24900 4472 24934 4506
rect 24900 4404 24934 4438
rect 24900 4336 24934 4370
rect 24900 4268 24934 4302
rect 24900 4200 24934 4234
rect 24900 4132 24934 4166
rect 24900 4064 24934 4098
rect 24900 3996 24934 4030
rect 24900 3928 24934 3962
rect 24900 3860 24934 3894
rect 24900 3792 24934 3826
rect 24900 3724 24934 3758
rect 24900 3656 24934 3690
rect 26286 4608 26320 4642
rect 26286 4540 26320 4574
rect 26286 4472 26320 4506
rect 26286 4404 26320 4438
rect 26286 4336 26320 4370
rect 26286 4268 26320 4302
rect 26286 4200 26320 4234
rect 26286 4132 26320 4166
rect 26286 4064 26320 4098
rect 26286 3996 26320 4030
rect 26286 3928 26320 3962
rect 26286 3860 26320 3894
rect 26286 3792 26320 3826
rect 26286 3724 26320 3758
rect 24900 3588 24934 3622
rect 26286 3656 26320 3690
rect 26286 3588 26320 3622
rect 25015 3480 25049 3514
rect 25083 3480 25117 3514
rect 25151 3480 25185 3514
rect 25219 3480 25253 3514
rect 25287 3480 25321 3514
rect 25355 3480 25389 3514
rect 25423 3480 25457 3514
rect 25491 3480 25525 3514
rect 25559 3480 25593 3514
rect 25627 3480 25661 3514
rect 25695 3480 25729 3514
rect 25763 3480 25797 3514
rect 25831 3480 25865 3514
rect 25899 3480 25933 3514
rect 25967 3480 26001 3514
rect 26035 3480 26069 3514
rect 26103 3480 26137 3514
rect 26171 3480 26205 3514
rect 36760 12281 36794 12315
rect 36828 12281 36862 12315
rect 36896 12281 36930 12315
rect 36964 12281 36998 12315
rect 37032 12281 37066 12315
rect 37100 12281 37134 12315
rect 37168 12281 37202 12315
rect 37236 12281 37270 12315
rect 37304 12281 37338 12315
rect 37372 12281 37406 12315
rect 37440 12281 37474 12315
rect 37508 12281 37542 12315
rect 37576 12281 37610 12315
rect 37644 12281 37678 12315
rect 37712 12281 37746 12315
rect 37780 12281 37814 12315
rect 37848 12281 37882 12315
rect 37916 12281 37950 12315
rect 37984 12281 38018 12315
rect 38052 12281 38086 12315
rect 38120 12281 38154 12315
rect 38188 12281 38222 12315
rect 38256 12281 38290 12315
rect 38324 12281 38358 12315
rect 38392 12281 38426 12315
rect 38460 12281 38494 12315
rect 38528 12281 38562 12315
rect 38596 12281 38630 12315
rect 38664 12281 38698 12315
rect 38732 12281 38766 12315
rect 38800 12281 38834 12315
rect 38868 12281 38902 12315
rect 38936 12281 38970 12315
rect 39004 12281 39038 12315
rect 39072 12281 39106 12315
rect 39140 12281 39174 12315
rect 39208 12281 39242 12315
rect 39276 12281 39310 12315
rect 39344 12281 39378 12315
rect 39412 12281 39446 12315
rect 39480 12281 39514 12315
rect 39548 12281 39582 12315
rect 39616 12281 39650 12315
rect 39684 12281 39718 12315
rect 39752 12281 39786 12315
rect 39820 12281 39854 12315
rect 39888 12281 39922 12315
rect 39956 12281 39990 12315
rect 40024 12281 40058 12315
rect 40092 12281 40126 12315
rect 40160 12281 40194 12315
rect 40228 12281 40262 12315
rect 40296 12281 40330 12315
rect 40364 12281 40398 12315
rect 40432 12281 40466 12315
rect 40500 12281 40534 12315
rect 40568 12281 40602 12315
rect 40636 12281 40670 12315
rect 40704 12281 40738 12315
rect 40772 12281 40806 12315
rect 40840 12281 40874 12315
rect 40908 12281 40942 12315
rect 40976 12281 41010 12315
rect 41044 12281 41078 12315
rect 41112 12281 41146 12315
rect 41180 12281 41214 12315
rect 41248 12281 41282 12315
rect 41316 12281 41350 12315
rect 41384 12281 41418 12315
rect 41452 12281 41486 12315
rect 41520 12281 41554 12315
rect 41588 12281 41622 12315
rect 41656 12281 41690 12315
rect 41724 12281 41758 12315
rect 41792 12281 41826 12315
rect 41860 12281 41894 12315
rect 41928 12281 41962 12315
rect 41996 12281 42030 12315
rect 36511 12091 36545 12125
rect 36511 12023 36545 12057
rect 42237 12051 42271 12085
rect 36511 11955 36545 11989
rect 36511 11887 36545 11921
rect 42237 11983 42271 12017
rect 42237 11915 42271 11949
rect 36511 11819 36545 11853
rect 36511 11751 36545 11785
rect 36511 11683 36545 11717
rect 36511 11615 36545 11649
rect 36511 11547 36545 11581
rect 36511 11479 36545 11513
rect 36511 11411 36545 11445
rect 36511 11343 36545 11377
rect 36511 11275 36545 11309
rect 36511 11207 36545 11241
rect 36511 11139 36545 11173
rect 36511 11071 36545 11105
rect 36511 11003 36545 11037
rect 36511 10935 36545 10969
rect 42237 11847 42271 11881
rect 42237 11779 42271 11813
rect 42237 11711 42271 11745
rect 42237 11643 42271 11677
rect 42237 11575 42271 11609
rect 42237 11507 42271 11541
rect 42237 11439 42271 11473
rect 42237 11371 42271 11405
rect 42237 11303 42271 11337
rect 42237 11235 42271 11269
rect 42237 11167 42271 11201
rect 42237 11099 42271 11133
rect 42237 11031 42271 11065
rect 42237 10963 42271 10997
rect 36511 10867 36545 10901
rect 36511 10799 36545 10833
rect 42237 10895 42271 10929
rect 42237 10827 42271 10861
rect 36511 10731 36545 10765
rect 36511 10663 36545 10697
rect 42237 10759 42271 10793
rect 42237 10691 42271 10725
rect 36511 10595 36545 10629
rect 36511 10527 36545 10561
rect 42237 10623 42271 10657
rect 42237 10555 42271 10589
rect 36511 10459 36545 10493
rect 36511 10391 36545 10425
rect 36511 10323 36545 10357
rect 36511 10255 36545 10289
rect 36511 10187 36545 10221
rect 36511 10119 36545 10153
rect 36511 10051 36545 10085
rect 36511 9983 36545 10017
rect 36511 9915 36545 9949
rect 36511 9847 36545 9881
rect 36511 9779 36545 9813
rect 36511 9711 36545 9745
rect 36511 9643 36545 9677
rect 36511 9575 36545 9609
rect 42237 10487 42271 10521
rect 42237 10419 42271 10453
rect 42237 10351 42271 10385
rect 42237 10283 42271 10317
rect 42237 10215 42271 10249
rect 42237 10147 42271 10181
rect 42237 10079 42271 10113
rect 42237 10011 42271 10045
rect 42237 9943 42271 9977
rect 42237 9875 42271 9909
rect 42237 9807 42271 9841
rect 42237 9739 42271 9773
rect 42237 9671 42271 9705
rect 42237 9603 42271 9637
rect 36511 9507 36545 9541
rect 36511 9439 36545 9473
rect 42237 9535 42271 9569
rect 42237 9467 42271 9501
rect 36511 9371 36545 9405
rect 42237 9399 42271 9433
rect 42237 9331 42271 9365
rect 36779 9115 36813 9149
rect 36847 9115 36881 9149
rect 36915 9115 36949 9149
rect 36983 9115 37017 9149
rect 37051 9115 37085 9149
rect 37119 9115 37153 9149
rect 37187 9115 37221 9149
rect 37255 9115 37289 9149
rect 37323 9115 37357 9149
rect 37391 9115 37425 9149
rect 37459 9115 37493 9149
rect 37527 9115 37561 9149
rect 37595 9115 37629 9149
rect 37663 9115 37697 9149
rect 37731 9115 37765 9149
rect 37799 9115 37833 9149
rect 37867 9115 37901 9149
rect 37935 9115 37969 9149
rect 38003 9115 38037 9149
rect 38071 9115 38105 9149
rect 38139 9115 38173 9149
rect 38207 9115 38241 9149
rect 38275 9115 38309 9149
rect 38343 9115 38377 9149
rect 38411 9115 38445 9149
rect 38479 9115 38513 9149
rect 38547 9115 38581 9149
rect 38615 9115 38649 9149
rect 38683 9115 38717 9149
rect 38751 9115 38785 9149
rect 38819 9115 38853 9149
rect 38887 9115 38921 9149
rect 38955 9115 38989 9149
rect 39023 9115 39057 9149
rect 39091 9115 39125 9149
rect 39159 9115 39193 9149
rect 39227 9115 39261 9149
rect 39295 9115 39329 9149
rect 39363 9115 39397 9149
rect 39431 9115 39465 9149
rect 39499 9115 39533 9149
rect 39567 9115 39601 9149
rect 39635 9115 39669 9149
rect 39703 9115 39737 9149
rect 39771 9115 39805 9149
rect 39839 9115 39873 9149
rect 39907 9115 39941 9149
rect 39975 9115 40009 9149
rect 40043 9115 40077 9149
rect 40111 9115 40145 9149
rect 40179 9115 40213 9149
rect 40247 9115 40281 9149
rect 40315 9115 40349 9149
rect 40383 9115 40417 9149
rect 40451 9115 40485 9149
rect 40519 9115 40553 9149
rect 40587 9115 40621 9149
rect 40655 9115 40689 9149
rect 40723 9115 40757 9149
rect 40791 9115 40825 9149
rect 40859 9115 40893 9149
rect 40927 9115 40961 9149
rect 40995 9115 41029 9149
rect 41063 9115 41097 9149
rect 41131 9115 41165 9149
rect 41199 9115 41233 9149
rect 41267 9115 41301 9149
rect 41335 9115 41369 9149
rect 41403 9115 41437 9149
rect 41471 9115 41505 9149
rect 41539 9115 41573 9149
rect 41607 9115 41641 9149
rect 41675 9115 41709 9149
rect 41743 9115 41777 9149
rect 41811 9115 41845 9149
rect 41879 9115 41913 9149
rect 41947 9115 41981 9149
rect 42015 9115 42049 9149
rect 37843 8575 37877 8609
rect 37911 8575 37945 8609
rect 37979 8575 38013 8609
rect 38047 8575 38081 8609
rect 38115 8575 38149 8609
rect 38183 8575 38217 8609
rect 38251 8575 38285 8609
rect 38319 8575 38353 8609
rect 38387 8575 38421 8609
rect 38455 8575 38489 8609
rect 38523 8575 38557 8609
rect 38591 8575 38625 8609
rect 38659 8575 38693 8609
rect 38727 8575 38761 8609
rect 38795 8575 38829 8609
rect 38863 8575 38897 8609
rect 38931 8575 38965 8609
rect 38999 8575 39033 8609
rect 39067 8575 39101 8609
rect 39135 8575 39169 8609
rect 39203 8575 39237 8609
rect 39271 8575 39305 8609
rect 39339 8575 39373 8609
rect 39407 8575 39441 8609
rect 39475 8575 39509 8609
rect 39543 8575 39577 8609
rect 39611 8575 39645 8609
rect 39679 8575 39713 8609
rect 39747 8575 39781 8609
rect 39815 8575 39849 8609
rect 39883 8575 39917 8609
rect 39951 8575 39985 8609
rect 40019 8575 40053 8609
rect 40087 8575 40121 8609
rect 40155 8575 40189 8609
rect 40223 8575 40257 8609
rect 40291 8575 40325 8609
rect 40359 8575 40393 8609
rect 40427 8575 40461 8609
rect 40495 8575 40529 8609
rect 40563 8575 40597 8609
rect 40631 8575 40665 8609
rect 40699 8575 40733 8609
rect 40767 8575 40801 8609
rect 40835 8575 40869 8609
rect 40903 8575 40937 8609
rect 40971 8575 41005 8609
rect 41039 8575 41073 8609
rect 41107 8575 41141 8609
rect 41175 8575 41209 8609
rect 41243 8575 41277 8609
rect 41311 8575 41345 8609
rect 41379 8575 41413 8609
rect 41447 8575 41481 8609
rect 41515 8575 41549 8609
rect 41583 8575 41617 8609
rect 41651 8575 41685 8609
rect 41719 8575 41753 8609
rect 41787 8575 41821 8609
rect 41855 8575 41889 8609
rect 41923 8575 41957 8609
rect 41991 8575 42025 8609
rect 37624 8398 37658 8432
rect 42136 8410 42170 8444
rect 37624 8330 37658 8364
rect 37624 8262 37658 8296
rect 42136 8342 42170 8376
rect 37624 8194 37658 8228
rect 37624 8126 37658 8160
rect 37624 8058 37658 8092
rect 37624 7990 37658 8024
rect 37624 7922 37658 7956
rect 37624 7854 37658 7888
rect 37624 7786 37658 7820
rect 37624 7718 37658 7752
rect 37624 7650 37658 7684
rect 37624 7582 37658 7616
rect 37624 7514 37658 7548
rect 37624 7446 37658 7480
rect 37624 7378 37658 7412
rect 37624 7310 37658 7344
rect 37624 7242 37658 7276
rect 37624 7174 37658 7208
rect 37624 7106 37658 7140
rect 37624 7038 37658 7072
rect 37624 6970 37658 7004
rect 37624 6902 37658 6936
rect 37624 6834 37658 6868
rect 37624 6766 37658 6800
rect 37624 6698 37658 6732
rect 37624 6630 37658 6664
rect 37624 6562 37658 6596
rect 37624 6494 37658 6528
rect 37624 6426 37658 6460
rect 37624 6358 37658 6392
rect 37624 6290 37658 6324
rect 42136 8274 42170 8308
rect 42136 8206 42170 8240
rect 42136 8138 42170 8172
rect 42136 8070 42170 8104
rect 42136 8002 42170 8036
rect 42136 7934 42170 7968
rect 42136 7866 42170 7900
rect 42136 7798 42170 7832
rect 42136 7730 42170 7764
rect 42136 7662 42170 7696
rect 42136 7594 42170 7628
rect 42136 7526 42170 7560
rect 42136 7458 42170 7492
rect 42136 7390 42170 7424
rect 42136 7322 42170 7356
rect 42136 7254 42170 7288
rect 42136 7186 42170 7220
rect 42136 7118 42170 7152
rect 42136 7050 42170 7084
rect 42136 6982 42170 7016
rect 42136 6914 42170 6948
rect 42136 6846 42170 6880
rect 42136 6778 42170 6812
rect 42136 6710 42170 6744
rect 42136 6642 42170 6676
rect 42136 6574 42170 6608
rect 42136 6506 42170 6540
rect 42136 6438 42170 6472
rect 42136 6370 42170 6404
rect 42136 6302 42170 6336
rect 37624 6222 37658 6256
rect 42136 6234 42170 6268
rect 37624 6154 37658 6188
rect 42136 6166 42170 6200
rect 37819 5995 37853 6029
rect 37887 5995 37921 6029
rect 37955 5995 37989 6029
rect 38023 5995 38057 6029
rect 38091 5995 38125 6029
rect 38159 5995 38193 6029
rect 38227 5995 38261 6029
rect 38295 5995 38329 6029
rect 38363 5995 38397 6029
rect 38431 5995 38465 6029
rect 38499 5995 38533 6029
rect 38567 5995 38601 6029
rect 38635 5995 38669 6029
rect 38703 5995 38737 6029
rect 38771 5995 38805 6029
rect 38839 5995 38873 6029
rect 38907 5995 38941 6029
rect 38975 5995 39009 6029
rect 39043 5995 39077 6029
rect 39111 5995 39145 6029
rect 39179 5995 39213 6029
rect 39247 5995 39281 6029
rect 39315 5995 39349 6029
rect 39383 5995 39417 6029
rect 39451 5995 39485 6029
rect 39519 5995 39553 6029
rect 39587 5995 39621 6029
rect 39655 5995 39689 6029
rect 39723 5995 39757 6029
rect 39791 5995 39825 6029
rect 39859 5995 39893 6029
rect 39927 5995 39961 6029
rect 39995 5995 40029 6029
rect 40063 5995 40097 6029
rect 40131 5995 40165 6029
rect 40199 5995 40233 6029
rect 40267 5995 40301 6029
rect 40335 5995 40369 6029
rect 40403 5995 40437 6029
rect 40471 5995 40505 6029
rect 40539 5995 40573 6029
rect 40607 5995 40641 6029
rect 40675 5995 40709 6029
rect 40743 5995 40777 6029
rect 40811 5995 40845 6029
rect 40879 5995 40913 6029
rect 40947 5995 40981 6029
rect 41015 5995 41049 6029
rect 41083 5995 41117 6029
rect 41151 5995 41185 6029
rect 41219 5995 41253 6029
rect 41287 5995 41321 6029
rect 41355 5995 41389 6029
rect 41423 5995 41457 6029
rect 41491 5995 41525 6029
rect 41559 5995 41593 6029
rect 41627 5995 41661 6029
rect 41695 5995 41729 6029
rect 41763 5995 41797 6029
rect 41831 5995 41865 6029
rect 41899 5995 41933 6029
rect 41967 5995 42001 6029
<< mvnsubdiffcont >>
rect 42576 19028 42610 19062
rect 42644 19028 42678 19062
rect 42712 19028 42746 19062
rect 42780 19028 42814 19062
rect 42848 19028 42882 19062
rect 42916 19028 42950 19062
rect 42984 19028 43018 19062
rect 43052 19028 43086 19062
rect 43120 19028 43154 19062
rect 43188 19028 43222 19062
rect 43256 19028 43290 19062
rect 43324 19028 43358 19062
rect 43392 19028 43426 19062
rect 43460 19028 43494 19062
rect 43528 19028 43562 19062
rect 43596 19028 43630 19062
rect 43664 19028 43698 19062
rect 43732 19028 43766 19062
rect 43800 19028 43834 19062
rect 43868 19028 43902 19062
rect 43936 19028 43970 19062
rect 44004 19028 44038 19062
rect 44072 19028 44106 19062
rect 44140 19028 44174 19062
rect 44208 19028 44242 19062
rect 44276 19028 44310 19062
rect 44344 19028 44378 19062
rect 44412 19028 44446 19062
rect 44480 19028 44514 19062
rect 44548 19028 44582 19062
rect 44616 19028 44650 19062
rect 44684 19028 44718 19062
rect 44752 19028 44786 19062
rect 44820 19028 44854 19062
rect 44888 19028 44922 19062
rect 44956 19028 44990 19062
rect 45024 19028 45058 19062
rect 45092 19028 45126 19062
rect 45160 19028 45194 19062
rect 45228 19028 45262 19062
rect 23161 18932 23195 18966
rect 23229 18932 23263 18966
rect 23297 18932 23331 18966
rect 23365 18932 23399 18966
rect 23433 18932 23467 18966
rect 23501 18932 23535 18966
rect 23569 18932 23603 18966
rect 23637 18932 23671 18966
rect 23705 18932 23739 18966
rect 23773 18932 23807 18966
rect 23841 18932 23875 18966
rect 23909 18932 23943 18966
rect 23977 18932 24011 18966
rect 24045 18932 24079 18966
rect 24113 18932 24147 18966
rect 24181 18932 24215 18966
rect 24249 18932 24283 18966
rect 23042 18808 23076 18842
rect 23042 18740 23076 18774
rect 24368 18808 24402 18842
rect 23042 18672 23076 18706
rect 23042 18604 23076 18638
rect 23042 18536 23076 18570
rect 23042 18468 23076 18502
rect 23042 18400 23076 18434
rect 23042 18332 23076 18366
rect -3016 18278 -2982 18312
rect -2948 18278 -2914 18312
rect -2880 18278 -2846 18312
rect -2812 18278 -2778 18312
rect -2744 18278 -2710 18312
rect -2676 18278 -2642 18312
rect -2608 18278 -2574 18312
rect -2540 18278 -2506 18312
rect -2472 18278 -2438 18312
rect -2404 18278 -2370 18312
rect -2336 18278 -2302 18312
rect -2268 18278 -2234 18312
rect -2200 18278 -2166 18312
rect -2132 18278 -2098 18312
rect -2064 18278 -2030 18312
rect -1996 18278 -1962 18312
rect -1928 18278 -1894 18312
rect -1860 18278 -1826 18312
rect -1792 18278 -1758 18312
rect -1724 18278 -1690 18312
rect -1656 18278 -1622 18312
rect -1588 18278 -1554 18312
rect -1520 18278 -1486 18312
rect -1452 18278 -1418 18312
rect -1384 18278 -1350 18312
rect -1316 18278 -1282 18312
rect -1248 18278 -1214 18312
rect -1180 18278 -1146 18312
rect -1112 18278 -1078 18312
rect -1044 18278 -1010 18312
rect -976 18278 -942 18312
rect -908 18278 -874 18312
rect -840 18278 -806 18312
rect -772 18278 -738 18312
rect -704 18278 -670 18312
rect -636 18278 -602 18312
rect -568 18278 -534 18312
rect -500 18278 -466 18312
rect -432 18278 -398 18312
rect -364 18278 -330 18312
rect -3114 18164 -3080 18198
rect -3114 18096 -3080 18130
rect -266 18164 -232 18198
rect -266 18096 -232 18130
rect -3114 18028 -3080 18062
rect -3114 17960 -3080 17994
rect -3114 17892 -3080 17926
rect -3114 17824 -3080 17858
rect -3114 17756 -3080 17790
rect -3114 17688 -3080 17722
rect -3114 17620 -3080 17654
rect -6702 17502 -6668 17536
rect -6634 17502 -6600 17536
rect -6566 17502 -6532 17536
rect -6498 17502 -6464 17536
rect -6430 17502 -6396 17536
rect -6362 17502 -6328 17536
rect -6294 17502 -6260 17536
rect -6226 17502 -6192 17536
rect -6158 17502 -6124 17536
rect -6090 17502 -6056 17536
rect -6022 17502 -5988 17536
rect -5954 17502 -5920 17536
rect -5886 17502 -5852 17536
rect -5818 17502 -5784 17536
rect -5750 17502 -5716 17536
rect -5682 17502 -5648 17536
rect -5614 17502 -5580 17536
rect -6798 17407 -6764 17441
rect -6798 17339 -6764 17373
rect -5508 17427 -5474 17461
rect -5508 17359 -5474 17393
rect -6798 17271 -6764 17305
rect -6798 17203 -6764 17237
rect -5508 17291 -5474 17325
rect -6798 17135 -6764 17169
rect -6798 17067 -6764 17101
rect -6798 16999 -6764 17033
rect -6798 16931 -6764 16965
rect -6798 16863 -6764 16897
rect -6798 16795 -6764 16829
rect -6798 16727 -6764 16761
rect -6798 16659 -6764 16693
rect -6798 16591 -6764 16625
rect -6798 16523 -6764 16557
rect -6798 16455 -6764 16489
rect -6798 16387 -6764 16421
rect -6798 16319 -6764 16353
rect -6798 16251 -6764 16285
rect -5508 17223 -5474 17257
rect -5508 17155 -5474 17189
rect -5508 17087 -5474 17121
rect -5508 17019 -5474 17053
rect -5508 16951 -5474 16985
rect -5508 16883 -5474 16917
rect -5508 16815 -5474 16849
rect -5508 16747 -5474 16781
rect -5508 16679 -5474 16713
rect -5508 16611 -5474 16645
rect -5508 16543 -5474 16577
rect -5508 16475 -5474 16509
rect -5508 16407 -5474 16441
rect -5508 16339 -5474 16373
rect -5508 16271 -5474 16305
rect -6798 16183 -6764 16217
rect -6798 16115 -6764 16149
rect -5508 16203 -5474 16237
rect -5508 16135 -5474 16169
rect -6798 16047 -6764 16081
rect -5508 16067 -5474 16101
rect -6682 15962 -6648 15996
rect -6614 15962 -6580 15996
rect -6546 15962 -6512 15996
rect -6478 15962 -6444 15996
rect -6410 15962 -6376 15996
rect -6342 15962 -6308 15996
rect -6274 15962 -6240 15996
rect -6206 15962 -6172 15996
rect -6138 15962 -6104 15996
rect -6070 15962 -6036 15996
rect -6002 15962 -5968 15996
rect -5934 15962 -5900 15996
rect -5866 15962 -5832 15996
rect -5798 15962 -5764 15996
rect -5730 15962 -5696 15996
rect -5662 15962 -5628 15996
rect -5594 15962 -5560 15996
rect -3114 17552 -3080 17586
rect -3114 17484 -3080 17518
rect -3114 17416 -3080 17450
rect -3114 17348 -3080 17382
rect -3114 17280 -3080 17314
rect -3114 17212 -3080 17246
rect -3114 17144 -3080 17178
rect -3114 17076 -3080 17110
rect -3114 17008 -3080 17042
rect -3114 16940 -3080 16974
rect -3114 16872 -3080 16906
rect -3114 16804 -3080 16838
rect -3114 16736 -3080 16770
rect -3114 16668 -3080 16702
rect -3114 16600 -3080 16634
rect -3114 16532 -3080 16566
rect -3114 16464 -3080 16498
rect -3114 16396 -3080 16430
rect -3114 16328 -3080 16362
rect -3114 16260 -3080 16294
rect -3114 16192 -3080 16226
rect -3114 16124 -3080 16158
rect -266 18028 -232 18062
rect -266 17960 -232 17994
rect -266 17892 -232 17926
rect -266 17824 -232 17858
rect -266 17756 -232 17790
rect -266 17688 -232 17722
rect -266 17620 -232 17654
rect -266 17552 -232 17586
rect -266 17484 -232 17518
rect 23042 18264 23076 18298
rect 23042 18196 23076 18230
rect 23042 18128 23076 18162
rect 23042 18060 23076 18094
rect 23042 17992 23076 18026
rect 23042 17924 23076 17958
rect 23042 17856 23076 17890
rect 23042 17788 23076 17822
rect 23042 17720 23076 17754
rect 24368 18740 24402 18774
rect 24368 18672 24402 18706
rect 24368 18604 24402 18638
rect 24368 18536 24402 18570
rect 24368 18468 24402 18502
rect 24368 18400 24402 18434
rect 24368 18332 24402 18366
rect 24368 18264 24402 18298
rect 24368 18196 24402 18230
rect 24368 18128 24402 18162
rect 24368 18060 24402 18094
rect 24368 17992 24402 18026
rect 24368 17924 24402 17958
rect 24368 17856 24402 17890
rect 24368 17788 24402 17822
rect 23042 17652 23076 17686
rect 24368 17720 24402 17754
rect 24368 17652 24402 17686
rect 23161 17528 23195 17562
rect 23229 17528 23263 17562
rect 23297 17528 23331 17562
rect 23365 17528 23399 17562
rect 23433 17528 23467 17562
rect 23501 17528 23535 17562
rect 23569 17528 23603 17562
rect 23637 17528 23671 17562
rect 23705 17528 23739 17562
rect 23773 17528 23807 17562
rect 23841 17528 23875 17562
rect 23909 17528 23943 17562
rect 23977 17528 24011 17562
rect 24045 17528 24079 17562
rect 24113 17528 24147 17562
rect 24181 17528 24215 17562
rect 24249 17528 24283 17562
rect 24681 18932 24715 18966
rect 24749 18932 24783 18966
rect 24817 18932 24851 18966
rect 24885 18932 24919 18966
rect 24953 18932 24987 18966
rect 25021 18932 25055 18966
rect 25089 18932 25123 18966
rect 25157 18932 25191 18966
rect 25225 18932 25259 18966
rect 25293 18932 25327 18966
rect 25361 18932 25395 18966
rect 25429 18932 25463 18966
rect 25497 18932 25531 18966
rect 25565 18932 25599 18966
rect 25633 18932 25667 18966
rect 25701 18932 25735 18966
rect 25769 18932 25803 18966
rect 25837 18932 25871 18966
rect 25905 18932 25939 18966
rect 25973 18932 26007 18966
rect 26041 18932 26075 18966
rect 26109 18932 26143 18966
rect 26177 18932 26211 18966
rect 26245 18932 26279 18966
rect 26313 18932 26347 18966
rect 26381 18932 26415 18966
rect 26449 18932 26483 18966
rect 26517 18932 26551 18966
rect 26585 18932 26619 18966
rect 26653 18932 26687 18966
rect 26721 18932 26755 18966
rect 26789 18932 26823 18966
rect 26857 18932 26891 18966
rect 26925 18932 26959 18966
rect 26993 18932 27027 18966
rect 27061 18932 27095 18966
rect 27129 18932 27163 18966
rect 27197 18932 27231 18966
rect 27265 18932 27299 18966
rect 27333 18932 27367 18966
rect 27401 18932 27435 18966
rect 27469 18932 27503 18966
rect 27537 18932 27571 18966
rect 27605 18932 27639 18966
rect 27673 18932 27707 18966
rect 27741 18932 27775 18966
rect 27809 18932 27843 18966
rect 27877 18932 27911 18966
rect 24558 18814 24592 18848
rect 24558 18746 24592 18780
rect 28000 18814 28034 18848
rect 24558 18678 24592 18712
rect 24558 18610 24592 18644
rect 24558 18542 24592 18576
rect 24558 18474 24592 18508
rect 24558 18406 24592 18440
rect 24558 18338 24592 18372
rect 24558 18270 24592 18304
rect 24558 18202 24592 18236
rect 24558 18134 24592 18168
rect 24558 18066 24592 18100
rect 24558 17998 24592 18032
rect 24558 17930 24592 17964
rect 24558 17862 24592 17896
rect 24558 17794 24592 17828
rect 24558 17726 24592 17760
rect 24558 17658 24592 17692
rect 24558 17590 24592 17624
rect 24558 17522 24592 17556
rect -266 17416 -232 17450
rect -266 17348 -232 17382
rect 24558 17454 24592 17488
rect 24558 17386 24592 17420
rect -266 17280 -232 17314
rect -266 17212 -232 17246
rect -266 17144 -232 17178
rect -266 17076 -232 17110
rect -266 17008 -232 17042
rect -266 16940 -232 16974
rect -266 16872 -232 16906
rect -266 16804 -232 16838
rect -266 16736 -232 16770
rect -266 16668 -232 16702
rect -266 16600 -232 16634
rect -266 16532 -232 16566
rect -266 16464 -232 16498
rect -266 16396 -232 16430
rect -266 16328 -232 16362
rect -266 16260 -232 16294
rect -266 16192 -232 16226
rect -266 16124 -232 16158
rect -3114 16056 -3080 16090
rect -3114 15988 -3080 16022
rect -266 16056 -232 16090
rect -266 15988 -232 16022
rect 24558 17318 24592 17352
rect 24558 17250 24592 17284
rect 24558 17182 24592 17216
rect 24558 17114 24592 17148
rect 28000 18746 28034 18780
rect 28000 18678 28034 18712
rect 28000 18610 28034 18644
rect 28000 18542 28034 18576
rect 28000 18474 28034 18508
rect 28000 18406 28034 18440
rect 28000 18338 28034 18372
rect 42478 18914 42512 18948
rect 42478 18846 42512 18880
rect 45326 18914 45360 18948
rect 45326 18846 45360 18880
rect 42478 18778 42512 18812
rect 42478 18710 42512 18744
rect 42478 18642 42512 18676
rect 42478 18574 42512 18608
rect 42478 18506 42512 18540
rect 42478 18438 42512 18472
rect 42478 18370 42512 18404
rect 28000 18270 28034 18304
rect 28000 18202 28034 18236
rect 28000 18134 28034 18168
rect 28000 18066 28034 18100
rect 28000 17998 28034 18032
rect 28000 17930 28034 17964
rect 28000 17862 28034 17896
rect 28000 17794 28034 17828
rect 28000 17726 28034 17760
rect 28000 17658 28034 17692
rect 28000 17590 28034 17624
rect 28000 17522 28034 17556
rect 28000 17454 28034 17488
rect 28000 17386 28034 17420
rect 28000 17318 28034 17352
rect 28000 17250 28034 17284
rect 28000 17182 28034 17216
rect 24558 17046 24592 17080
rect 28000 17114 28034 17148
rect 28000 17046 28034 17080
rect 24681 16928 24715 16962
rect 24749 16928 24783 16962
rect 24817 16928 24851 16962
rect 24885 16928 24919 16962
rect 24953 16928 24987 16962
rect 25021 16928 25055 16962
rect 25089 16928 25123 16962
rect 25157 16928 25191 16962
rect 25225 16928 25259 16962
rect 25293 16928 25327 16962
rect 25361 16928 25395 16962
rect 25429 16928 25463 16962
rect 25497 16928 25531 16962
rect 25565 16928 25599 16962
rect 25633 16928 25667 16962
rect 25701 16928 25735 16962
rect 25769 16928 25803 16962
rect 25837 16928 25871 16962
rect 25905 16928 25939 16962
rect 25973 16928 26007 16962
rect 26041 16928 26075 16962
rect 26109 16928 26143 16962
rect 26177 16928 26211 16962
rect 26245 16928 26279 16962
rect 26313 16928 26347 16962
rect 26381 16928 26415 16962
rect 26449 16928 26483 16962
rect 26517 16928 26551 16962
rect 26585 16928 26619 16962
rect 26653 16928 26687 16962
rect 26721 16928 26755 16962
rect 26789 16928 26823 16962
rect 26857 16928 26891 16962
rect 26925 16928 26959 16962
rect 26993 16928 27027 16962
rect 27061 16928 27095 16962
rect 27129 16928 27163 16962
rect 27197 16928 27231 16962
rect 27265 16928 27299 16962
rect 27333 16928 27367 16962
rect 27401 16928 27435 16962
rect 27469 16928 27503 16962
rect 27537 16928 27571 16962
rect 27605 16928 27639 16962
rect 27673 16928 27707 16962
rect 27741 16928 27775 16962
rect 27809 16928 27843 16962
rect 27877 16928 27911 16962
rect 38890 18252 38924 18286
rect 38958 18252 38992 18286
rect 39026 18252 39060 18286
rect 39094 18252 39128 18286
rect 39162 18252 39196 18286
rect 39230 18252 39264 18286
rect 39298 18252 39332 18286
rect 39366 18252 39400 18286
rect 39434 18252 39468 18286
rect 39502 18252 39536 18286
rect 39570 18252 39604 18286
rect 39638 18252 39672 18286
rect 39706 18252 39740 18286
rect 39774 18252 39808 18286
rect 39842 18252 39876 18286
rect 39910 18252 39944 18286
rect 39978 18252 40012 18286
rect 38794 18157 38828 18191
rect 38794 18089 38828 18123
rect 40084 18177 40118 18211
rect 40084 18109 40118 18143
rect 38794 18021 38828 18055
rect 38794 17953 38828 17987
rect 40084 18041 40118 18075
rect 38794 17885 38828 17919
rect 38794 17817 38828 17851
rect 38794 17749 38828 17783
rect 38794 17681 38828 17715
rect 38794 17613 38828 17647
rect 38794 17545 38828 17579
rect 38794 17477 38828 17511
rect 38794 17409 38828 17443
rect 38794 17341 38828 17375
rect 38794 17273 38828 17307
rect 38794 17205 38828 17239
rect 38794 17137 38828 17171
rect 38794 17069 38828 17103
rect 38794 17001 38828 17035
rect 40084 17973 40118 18007
rect 40084 17905 40118 17939
rect 40084 17837 40118 17871
rect 40084 17769 40118 17803
rect 40084 17701 40118 17735
rect 40084 17633 40118 17667
rect 40084 17565 40118 17599
rect 40084 17497 40118 17531
rect 40084 17429 40118 17463
rect 40084 17361 40118 17395
rect 40084 17293 40118 17327
rect 40084 17225 40118 17259
rect 40084 17157 40118 17191
rect 40084 17089 40118 17123
rect 40084 17021 40118 17055
rect 38794 16933 38828 16967
rect 38794 16865 38828 16899
rect 40084 16953 40118 16987
rect 40084 16885 40118 16919
rect 38794 16797 38828 16831
rect 40084 16817 40118 16851
rect 38910 16712 38944 16746
rect 38978 16712 39012 16746
rect 39046 16712 39080 16746
rect 39114 16712 39148 16746
rect 39182 16712 39216 16746
rect 39250 16712 39284 16746
rect 39318 16712 39352 16746
rect 39386 16712 39420 16746
rect 39454 16712 39488 16746
rect 39522 16712 39556 16746
rect 39590 16712 39624 16746
rect 39658 16712 39692 16746
rect 39726 16712 39760 16746
rect 39794 16712 39828 16746
rect 39862 16712 39896 16746
rect 39930 16712 39964 16746
rect 39998 16712 40032 16746
rect 42478 18302 42512 18336
rect 42478 18234 42512 18268
rect 42478 18166 42512 18200
rect 42478 18098 42512 18132
rect 42478 18030 42512 18064
rect 42478 17962 42512 17996
rect 42478 17894 42512 17928
rect 42478 17826 42512 17860
rect 42478 17758 42512 17792
rect 42478 17690 42512 17724
rect 42478 17622 42512 17656
rect 42478 17554 42512 17588
rect 42478 17486 42512 17520
rect 42478 17418 42512 17452
rect 42478 17350 42512 17384
rect 42478 17282 42512 17316
rect 42478 17214 42512 17248
rect 42478 17146 42512 17180
rect 42478 17078 42512 17112
rect 42478 17010 42512 17044
rect 42478 16942 42512 16976
rect 42478 16874 42512 16908
rect 45326 18778 45360 18812
rect 45326 18710 45360 18744
rect 45326 18642 45360 18676
rect 45326 18574 45360 18608
rect 45326 18506 45360 18540
rect 45326 18438 45360 18472
rect 45326 18370 45360 18404
rect 45326 18302 45360 18336
rect 45326 18234 45360 18268
rect 45326 18166 45360 18200
rect 45326 18098 45360 18132
rect 45326 18030 45360 18064
rect 45326 17962 45360 17996
rect 45326 17894 45360 17928
rect 45326 17826 45360 17860
rect 45326 17758 45360 17792
rect 45326 17690 45360 17724
rect 45326 17622 45360 17656
rect 45326 17554 45360 17588
rect 45326 17486 45360 17520
rect 45326 17418 45360 17452
rect 45326 17350 45360 17384
rect 45326 17282 45360 17316
rect 45326 17214 45360 17248
rect 45326 17146 45360 17180
rect 45326 17078 45360 17112
rect 45326 17010 45360 17044
rect 45326 16942 45360 16976
rect 45326 16874 45360 16908
rect 42478 16806 42512 16840
rect 42478 16738 42512 16772
rect 45326 16806 45360 16840
rect 45326 16738 45360 16772
rect 42576 16624 42610 16658
rect 42644 16624 42678 16658
rect 42712 16624 42746 16658
rect 42780 16624 42814 16658
rect 42848 16624 42882 16658
rect 42916 16624 42950 16658
rect 42984 16624 43018 16658
rect 43052 16624 43086 16658
rect 43120 16624 43154 16658
rect 43188 16624 43222 16658
rect 43256 16624 43290 16658
rect 43324 16624 43358 16658
rect 43392 16624 43426 16658
rect 43460 16624 43494 16658
rect 43528 16624 43562 16658
rect 43596 16624 43630 16658
rect 43664 16624 43698 16658
rect 43732 16624 43766 16658
rect 43800 16624 43834 16658
rect 43868 16624 43902 16658
rect 43936 16624 43970 16658
rect 44004 16624 44038 16658
rect 44072 16624 44106 16658
rect 44140 16624 44174 16658
rect 44208 16624 44242 16658
rect 44276 16624 44310 16658
rect 44344 16624 44378 16658
rect 44412 16624 44446 16658
rect 44480 16624 44514 16658
rect 44548 16624 44582 16658
rect 44616 16624 44650 16658
rect 44684 16624 44718 16658
rect 44752 16624 44786 16658
rect 44820 16624 44854 16658
rect 44888 16624 44922 16658
rect 44956 16624 44990 16658
rect 45024 16624 45058 16658
rect 45092 16624 45126 16658
rect 45160 16624 45194 16658
rect 45228 16624 45262 16658
rect -3016 15874 -2982 15908
rect -2948 15874 -2914 15908
rect -2880 15874 -2846 15908
rect -2812 15874 -2778 15908
rect -2744 15874 -2710 15908
rect -2676 15874 -2642 15908
rect -2608 15874 -2574 15908
rect -2540 15874 -2506 15908
rect -2472 15874 -2438 15908
rect -2404 15874 -2370 15908
rect -2336 15874 -2302 15908
rect -2268 15874 -2234 15908
rect -2200 15874 -2166 15908
rect -2132 15874 -2098 15908
rect -2064 15874 -2030 15908
rect -1996 15874 -1962 15908
rect -1928 15874 -1894 15908
rect -1860 15874 -1826 15908
rect -1792 15874 -1758 15908
rect -1724 15874 -1690 15908
rect -1656 15874 -1622 15908
rect -1588 15874 -1554 15908
rect -1520 15874 -1486 15908
rect -1452 15874 -1418 15908
rect -1384 15874 -1350 15908
rect -1316 15874 -1282 15908
rect -1248 15874 -1214 15908
rect -1180 15874 -1146 15908
rect -1112 15874 -1078 15908
rect -1044 15874 -1010 15908
rect -976 15874 -942 15908
rect -908 15874 -874 15908
rect -840 15874 -806 15908
rect -772 15874 -738 15908
rect -704 15874 -670 15908
rect -636 15874 -602 15908
rect -568 15874 -534 15908
rect -500 15874 -466 15908
rect -432 15874 -398 15908
rect -364 15874 -330 15908
rect 12964 14952 12998 14986
rect 13032 14952 13066 14986
rect 13100 14952 13134 14986
rect 13168 14952 13202 14986
rect 13236 14952 13270 14986
rect 13304 14952 13338 14986
rect 13372 14952 13406 14986
rect 13440 14952 13474 14986
rect 13508 14952 13542 14986
rect 13576 14952 13610 14986
rect 13644 14952 13678 14986
rect 13712 14952 13746 14986
rect 13780 14952 13814 14986
rect 13848 14952 13882 14986
rect 13916 14952 13950 14986
rect 13984 14952 14018 14986
rect 14052 14952 14086 14986
rect 14120 14952 14154 14986
rect 14188 14952 14222 14986
rect 14256 14952 14290 14986
rect 14324 14952 14358 14986
rect 14392 14952 14426 14986
rect 14460 14952 14494 14986
rect 14528 14952 14562 14986
rect 14596 14952 14630 14986
rect 14664 14952 14698 14986
rect 14732 14952 14766 14986
rect 14800 14952 14834 14986
rect 14868 14952 14902 14986
rect 14936 14952 14970 14986
rect 15004 14952 15038 14986
rect 15072 14952 15106 14986
rect 15140 14952 15174 14986
rect 12860 14848 12894 14882
rect 12860 14780 12894 14814
rect 15244 14848 15278 14882
rect 15244 14780 15278 14814
rect 12860 14712 12894 14746
rect 12860 14644 12894 14678
rect 12860 14576 12894 14610
rect 12860 14508 12894 14542
rect 12860 14440 12894 14474
rect 12860 14372 12894 14406
rect 12860 14304 12894 14338
rect 12860 14236 12894 14270
rect 12860 14168 12894 14202
rect 12860 14100 12894 14134
rect 12860 14032 12894 14066
rect 12860 13964 12894 13998
rect 12860 13896 12894 13930
rect 12860 13828 12894 13862
rect 12860 13760 12894 13794
rect 12860 13692 12894 13726
rect 12860 13624 12894 13658
rect 12860 13556 12894 13590
rect 12860 13488 12894 13522
rect 12860 13420 12894 13454
rect 12860 13352 12894 13386
rect 12860 13284 12894 13318
rect 12860 13216 12894 13250
rect 12860 13148 12894 13182
rect 12860 13080 12894 13114
rect 12860 13012 12894 13046
rect 12860 12944 12894 12978
rect 12860 12876 12894 12910
rect 12860 12808 12894 12842
rect 12860 12740 12894 12774
rect 12860 12672 12894 12706
rect 12860 12604 12894 12638
rect 12860 12536 12894 12570
rect 12860 12468 12894 12502
rect 12860 12400 12894 12434
rect 12860 12332 12894 12366
rect 12860 12264 12894 12298
rect 12860 12196 12894 12230
rect 12860 12128 12894 12162
rect 12860 12060 12894 12094
rect 12860 11992 12894 12026
rect 12860 11924 12894 11958
rect 12860 11856 12894 11890
rect 12860 11788 12894 11822
rect 15244 14712 15278 14746
rect 15244 14644 15278 14678
rect 15244 14576 15278 14610
rect 15244 14508 15278 14542
rect 15244 14440 15278 14474
rect 15244 14372 15278 14406
rect 15244 14304 15278 14338
rect 15244 14236 15278 14270
rect 15244 14168 15278 14202
rect 15244 14100 15278 14134
rect 15244 14032 15278 14066
rect 15244 13964 15278 13998
rect 15244 13896 15278 13930
rect 15244 13828 15278 13862
rect 15244 13760 15278 13794
rect 15244 13692 15278 13726
rect 15244 13624 15278 13658
rect 15244 13556 15278 13590
rect 15244 13488 15278 13522
rect 15244 13420 15278 13454
rect 15244 13352 15278 13386
rect 15244 13284 15278 13318
rect 15244 13216 15278 13250
rect 15244 13148 15278 13182
rect 15244 13080 15278 13114
rect 15244 13012 15278 13046
rect 15244 12944 15278 12978
rect 15244 12876 15278 12910
rect 15244 12808 15278 12842
rect 15244 12740 15278 12774
rect 15244 12672 15278 12706
rect 15244 12604 15278 12638
rect 15244 12536 15278 12570
rect 15244 12468 15278 12502
rect 15244 12400 15278 12434
rect 15244 12332 15278 12366
rect 15244 12264 15278 12298
rect 15244 12196 15278 12230
rect 15244 12128 15278 12162
rect 15244 12060 15278 12094
rect 15244 11992 15278 12026
rect 15244 11924 15278 11958
rect 15244 11856 15278 11890
rect 15244 11788 15278 11822
rect 12860 11720 12894 11754
rect 12860 11652 12894 11686
rect 15244 11720 15278 11754
rect 15244 11652 15278 11686
rect 12964 11548 12998 11582
rect 13032 11548 13066 11582
rect 13100 11548 13134 11582
rect 13168 11548 13202 11582
rect 13236 11548 13270 11582
rect 13304 11548 13338 11582
rect 13372 11548 13406 11582
rect 13440 11548 13474 11582
rect 13508 11548 13542 11582
rect 13576 11548 13610 11582
rect 13644 11548 13678 11582
rect 13712 11548 13746 11582
rect 13780 11548 13814 11582
rect 13848 11548 13882 11582
rect 13916 11548 13950 11582
rect 13984 11548 14018 11582
rect 14052 11548 14086 11582
rect 14120 11548 14154 11582
rect 14188 11548 14222 11582
rect 14256 11548 14290 11582
rect 14324 11548 14358 11582
rect 14392 11548 14426 11582
rect 14460 11548 14494 11582
rect 14528 11548 14562 11582
rect 14596 11548 14630 11582
rect 14664 11548 14698 11582
rect 14732 11548 14766 11582
rect 14800 11548 14834 11582
rect 14868 11548 14902 11582
rect 14936 11548 14970 11582
rect 15004 11548 15038 11582
rect 15072 11548 15106 11582
rect 15140 11548 15174 11582
rect 15549 14952 15583 14986
rect 15617 14952 15651 14986
rect 15685 14952 15719 14986
rect 15753 14952 15787 14986
rect 15821 14952 15855 14986
rect 15889 14952 15923 14986
rect 15957 14952 15991 14986
rect 16025 14952 16059 14986
rect 16093 14952 16127 14986
rect 16161 14952 16195 14986
rect 16229 14952 16263 14986
rect 16297 14952 16331 14986
rect 16365 14952 16399 14986
rect 16433 14952 16467 14986
rect 16501 14952 16535 14986
rect 16569 14952 16603 14986
rect 16637 14952 16671 14986
rect 15430 14848 15464 14882
rect 15430 14780 15464 14814
rect 16756 14848 16790 14882
rect 16756 14780 16790 14814
rect 15430 14712 15464 14746
rect 15430 14644 15464 14678
rect 15430 14576 15464 14610
rect 15430 14508 15464 14542
rect 15430 14440 15464 14474
rect 15430 14372 15464 14406
rect 15430 14304 15464 14338
rect 15430 14236 15464 14270
rect 15430 14168 15464 14202
rect 15430 14100 15464 14134
rect 15430 14032 15464 14066
rect 15430 13964 15464 13998
rect 15430 13896 15464 13930
rect 15430 13828 15464 13862
rect 15430 13760 15464 13794
rect 15430 13692 15464 13726
rect 15430 13624 15464 13658
rect 15430 13556 15464 13590
rect 15430 13488 15464 13522
rect 15430 13420 15464 13454
rect 15430 13352 15464 13386
rect 15430 13284 15464 13318
rect 15430 13216 15464 13250
rect 15430 13148 15464 13182
rect 15430 13080 15464 13114
rect 15430 13012 15464 13046
rect 15430 12944 15464 12978
rect 15430 12876 15464 12910
rect 15430 12808 15464 12842
rect 15430 12740 15464 12774
rect 15430 12672 15464 12706
rect 15430 12604 15464 12638
rect 15430 12536 15464 12570
rect 15430 12468 15464 12502
rect 15430 12400 15464 12434
rect 15430 12332 15464 12366
rect 15430 12264 15464 12298
rect 15430 12196 15464 12230
rect 15430 12128 15464 12162
rect 15430 12060 15464 12094
rect 15430 11992 15464 12026
rect 15430 11924 15464 11958
rect 15430 11856 15464 11890
rect 15430 11788 15464 11822
rect 16756 14712 16790 14746
rect 16756 14644 16790 14678
rect 16756 14576 16790 14610
rect 16756 14508 16790 14542
rect 16756 14440 16790 14474
rect 16756 14372 16790 14406
rect 16756 14304 16790 14338
rect 16756 14236 16790 14270
rect 16756 14168 16790 14202
rect 16756 14100 16790 14134
rect 16756 14032 16790 14066
rect 16756 13964 16790 13998
rect 16756 13896 16790 13930
rect 16756 13828 16790 13862
rect 16756 13760 16790 13794
rect 16756 13692 16790 13726
rect 16756 13624 16790 13658
rect 16756 13556 16790 13590
rect 16756 13488 16790 13522
rect 16756 13420 16790 13454
rect 16756 13352 16790 13386
rect 16756 13284 16790 13318
rect 16756 13216 16790 13250
rect 16756 13148 16790 13182
rect 16756 13080 16790 13114
rect 16756 13012 16790 13046
rect 16756 12944 16790 12978
rect 16756 12876 16790 12910
rect 16756 12808 16790 12842
rect 16756 12740 16790 12774
rect 16756 12672 16790 12706
rect 16756 12604 16790 12638
rect 16756 12536 16790 12570
rect 16756 12468 16790 12502
rect 16756 12400 16790 12434
rect 16756 12332 16790 12366
rect 16756 12264 16790 12298
rect 16756 12196 16790 12230
rect 16756 12128 16790 12162
rect 16756 12060 16790 12094
rect 16756 11992 16790 12026
rect 16756 11924 16790 11958
rect 16756 11856 16790 11890
rect 16756 11788 16790 11822
rect 15430 11720 15464 11754
rect 15430 11652 15464 11686
rect 16756 11720 16790 11754
rect 16756 11652 16790 11686
rect 15549 11548 15583 11582
rect 15617 11548 15651 11582
rect 15685 11548 15719 11582
rect 15753 11548 15787 11582
rect 15821 11548 15855 11582
rect 15889 11548 15923 11582
rect 15957 11548 15991 11582
rect 16025 11548 16059 11582
rect 16093 11548 16127 11582
rect 16161 11548 16195 11582
rect 16229 11548 16263 11582
rect 16297 11548 16331 11582
rect 16365 11548 16399 11582
rect 16433 11548 16467 11582
rect 16501 11548 16535 11582
rect 16569 11548 16603 11582
rect 16637 11548 16671 11582
rect 17059 14962 17093 14996
rect 17127 14962 17161 14996
rect 17195 14962 17229 14996
rect 17263 14962 17297 14996
rect 17331 14962 17365 14996
rect 17399 14962 17433 14996
rect 17467 14962 17501 14996
rect 17535 14962 17569 14996
rect 17603 14962 17637 14996
rect 17671 14962 17705 14996
rect 17739 14962 17773 14996
rect 17807 14962 17841 14996
rect 17875 14962 17909 14996
rect 17943 14962 17977 14996
rect 18011 14962 18045 14996
rect 18079 14962 18113 14996
rect 18147 14962 18181 14996
rect 16940 14858 16974 14892
rect 16940 14790 16974 14824
rect 18266 14858 18300 14892
rect 18266 14790 18300 14824
rect 16940 14722 16974 14756
rect 16940 14654 16974 14688
rect 16940 14586 16974 14620
rect 16940 14518 16974 14552
rect 16940 14450 16974 14484
rect 16940 14382 16974 14416
rect 16940 14314 16974 14348
rect 16940 14246 16974 14280
rect 16940 14178 16974 14212
rect 16940 14110 16974 14144
rect 16940 14042 16974 14076
rect 16940 13974 16974 14008
rect 16940 13906 16974 13940
rect 16940 13838 16974 13872
rect 16940 13770 16974 13804
rect 16940 13702 16974 13736
rect 16940 13634 16974 13668
rect 16940 13566 16974 13600
rect 16940 13498 16974 13532
rect 16940 13430 16974 13464
rect 16940 13362 16974 13396
rect 16940 13294 16974 13328
rect 16940 13226 16974 13260
rect 16940 13158 16974 13192
rect 16940 13090 16974 13124
rect 16940 13022 16974 13056
rect 16940 12954 16974 12988
rect 16940 12886 16974 12920
rect 16940 12818 16974 12852
rect 16940 12750 16974 12784
rect 16940 12682 16974 12716
rect 16940 12614 16974 12648
rect 16940 12546 16974 12580
rect 16940 12478 16974 12512
rect 16940 12410 16974 12444
rect 16940 12342 16974 12376
rect 16940 12274 16974 12308
rect 16940 12206 16974 12240
rect 16940 12138 16974 12172
rect 16940 12070 16974 12104
rect 16940 12002 16974 12036
rect 16940 11934 16974 11968
rect 16940 11866 16974 11900
rect 16940 11798 16974 11832
rect 18266 14722 18300 14756
rect 18266 14654 18300 14688
rect 18266 14586 18300 14620
rect 18266 14518 18300 14552
rect 18266 14450 18300 14484
rect 18266 14382 18300 14416
rect 18266 14314 18300 14348
rect 18266 14246 18300 14280
rect 18266 14178 18300 14212
rect 18266 14110 18300 14144
rect 18266 14042 18300 14076
rect 18266 13974 18300 14008
rect 18266 13906 18300 13940
rect 18266 13838 18300 13872
rect 18266 13770 18300 13804
rect 18266 13702 18300 13736
rect 18266 13634 18300 13668
rect 18266 13566 18300 13600
rect 18266 13498 18300 13532
rect 18266 13430 18300 13464
rect 18266 13362 18300 13396
rect 18266 13294 18300 13328
rect 18266 13226 18300 13260
rect 18266 13158 18300 13192
rect 18266 13090 18300 13124
rect 18266 13022 18300 13056
rect 18266 12954 18300 12988
rect 18266 12886 18300 12920
rect 18266 12818 18300 12852
rect 18266 12750 18300 12784
rect 18266 12682 18300 12716
rect 18266 12614 18300 12648
rect 18266 12546 18300 12580
rect 18266 12478 18300 12512
rect 18266 12410 18300 12444
rect 18266 12342 18300 12376
rect 18266 12274 18300 12308
rect 18266 12206 18300 12240
rect 18266 12138 18300 12172
rect 18266 12070 18300 12104
rect 18266 12002 18300 12036
rect 18266 11934 18300 11968
rect 18266 11866 18300 11900
rect 18266 11798 18300 11832
rect 16940 11730 16974 11764
rect 16940 11662 16974 11696
rect 18266 11730 18300 11764
rect 18266 11662 18300 11696
rect 17059 11558 17093 11592
rect 17127 11558 17161 11592
rect 17195 11558 17229 11592
rect 17263 11558 17297 11592
rect 17331 11558 17365 11592
rect 17399 11558 17433 11592
rect 17467 11558 17501 11592
rect 17535 11558 17569 11592
rect 17603 11558 17637 11592
rect 17671 11558 17705 11592
rect 17739 11558 17773 11592
rect 17807 11558 17841 11592
rect 17875 11558 17909 11592
rect 17943 11558 17977 11592
rect 18011 11558 18045 11592
rect 18079 11558 18113 11592
rect 18147 11558 18181 11592
rect 18523 14946 18557 14980
rect 18591 14946 18625 14980
rect 18659 14946 18693 14980
rect 18727 14946 18761 14980
rect 18795 14946 18829 14980
rect 18863 14946 18897 14980
rect 18931 14946 18965 14980
rect 18999 14946 19033 14980
rect 19067 14946 19101 14980
rect 19135 14946 19169 14980
rect 19203 14946 19237 14980
rect 19271 14946 19305 14980
rect 19339 14946 19373 14980
rect 19407 14946 19441 14980
rect 19475 14946 19509 14980
rect 19543 14946 19577 14980
rect 19611 14946 19645 14980
rect 18404 14842 18438 14876
rect 18404 14774 18438 14808
rect 19730 14842 19764 14876
rect 19730 14774 19764 14808
rect 18404 14706 18438 14740
rect 18404 14638 18438 14672
rect 18404 14570 18438 14604
rect 18404 14502 18438 14536
rect 18404 14434 18438 14468
rect 18404 14366 18438 14400
rect 18404 14298 18438 14332
rect 18404 14230 18438 14264
rect 18404 14162 18438 14196
rect 18404 14094 18438 14128
rect 18404 14026 18438 14060
rect 18404 13958 18438 13992
rect 18404 13890 18438 13924
rect 18404 13822 18438 13856
rect 18404 13754 18438 13788
rect 18404 13686 18438 13720
rect 18404 13618 18438 13652
rect 18404 13550 18438 13584
rect 18404 13482 18438 13516
rect 18404 13414 18438 13448
rect 18404 13346 18438 13380
rect 18404 13278 18438 13312
rect 18404 13210 18438 13244
rect 18404 13142 18438 13176
rect 18404 13074 18438 13108
rect 18404 13006 18438 13040
rect 18404 12938 18438 12972
rect 18404 12870 18438 12904
rect 18404 12802 18438 12836
rect 18404 12734 18438 12768
rect 18404 12666 18438 12700
rect 18404 12598 18438 12632
rect 18404 12530 18438 12564
rect 18404 12462 18438 12496
rect 18404 12394 18438 12428
rect 18404 12326 18438 12360
rect 18404 12258 18438 12292
rect 18404 12190 18438 12224
rect 18404 12122 18438 12156
rect 18404 12054 18438 12088
rect 18404 11986 18438 12020
rect 18404 11918 18438 11952
rect 18404 11850 18438 11884
rect 18404 11782 18438 11816
rect 19730 14706 19764 14740
rect 19730 14638 19764 14672
rect 19730 14570 19764 14604
rect 19730 14502 19764 14536
rect 19730 14434 19764 14468
rect 19730 14366 19764 14400
rect 19730 14298 19764 14332
rect 19730 14230 19764 14264
rect 19730 14162 19764 14196
rect 19730 14094 19764 14128
rect 19730 14026 19764 14060
rect 19730 13958 19764 13992
rect 19730 13890 19764 13924
rect 19730 13822 19764 13856
rect 19730 13754 19764 13788
rect 19730 13686 19764 13720
rect 19730 13618 19764 13652
rect 19730 13550 19764 13584
rect 19730 13482 19764 13516
rect 19730 13414 19764 13448
rect 19730 13346 19764 13380
rect 19730 13278 19764 13312
rect 19730 13210 19764 13244
rect 19730 13142 19764 13176
rect 19730 13074 19764 13108
rect 19730 13006 19764 13040
rect 19730 12938 19764 12972
rect 19730 12870 19764 12904
rect 19730 12802 19764 12836
rect 19730 12734 19764 12768
rect 19730 12666 19764 12700
rect 19730 12598 19764 12632
rect 19730 12530 19764 12564
rect 19730 12462 19764 12496
rect 19730 12394 19764 12428
rect 19730 12326 19764 12360
rect 19730 12258 19764 12292
rect 19730 12190 19764 12224
rect 19730 12122 19764 12156
rect 19730 12054 19764 12088
rect 19730 11986 19764 12020
rect 19730 11918 19764 11952
rect 19730 11850 19764 11884
rect 19730 11782 19764 11816
rect 18404 11714 18438 11748
rect 18404 11646 18438 11680
rect 19730 11714 19764 11748
rect 19730 11646 19764 11680
rect 18523 11542 18557 11576
rect 18591 11542 18625 11576
rect 18659 11542 18693 11576
rect 18727 11542 18761 11576
rect 18795 11542 18829 11576
rect 18863 11542 18897 11576
rect 18931 11542 18965 11576
rect 18999 11542 19033 11576
rect 19067 11542 19101 11576
rect 19135 11542 19169 11576
rect 19203 11542 19237 11576
rect 19271 11542 19305 11576
rect 19339 11542 19373 11576
rect 19407 11542 19441 11576
rect 19475 11542 19509 11576
rect 19543 11542 19577 11576
rect 19611 11542 19645 11576
rect 14924 11432 14958 11466
rect 14992 11432 15026 11466
rect 15060 11432 15094 11466
rect 15128 11432 15162 11466
rect 15196 11432 15230 11466
rect 15264 11432 15298 11466
rect 15332 11432 15366 11466
rect 15400 11432 15434 11466
rect 15468 11432 15502 11466
rect 15536 11432 15570 11466
rect 15604 11432 15638 11466
rect 15672 11432 15706 11466
rect 15740 11432 15774 11466
rect 15808 11432 15842 11466
rect 15876 11432 15910 11466
rect 15944 11432 15978 11466
rect 16012 11432 16046 11466
rect 16080 11432 16114 11466
rect 16148 11432 16182 11466
rect 16216 11432 16250 11466
rect 16284 11432 16318 11466
rect 16352 11432 16386 11466
rect 16420 11432 16454 11466
rect 16488 11432 16522 11466
rect 16556 11432 16590 11466
rect 16624 11432 16658 11466
rect 16692 11432 16726 11466
rect 16760 11432 16794 11466
rect 16828 11432 16862 11466
rect 16896 11432 16930 11466
rect 16964 11432 16998 11466
rect 17032 11432 17066 11466
rect 17100 11432 17134 11466
rect 14820 11328 14854 11362
rect 14820 11260 14854 11294
rect 17204 11328 17238 11362
rect 17204 11260 17238 11294
rect 14820 11192 14854 11226
rect 14820 11124 14854 11158
rect 14820 11056 14854 11090
rect 14820 10988 14854 11022
rect 14820 10920 14854 10954
rect 14820 10852 14854 10886
rect 14820 10784 14854 10818
rect 14820 10716 14854 10750
rect 14820 10648 14854 10682
rect 14820 10580 14854 10614
rect 14820 10512 14854 10546
rect 14820 10444 14854 10478
rect 14820 10376 14854 10410
rect 14820 10308 14854 10342
rect 14820 10240 14854 10274
rect 14820 10172 14854 10206
rect 14820 10104 14854 10138
rect 14820 10036 14854 10070
rect 14820 9968 14854 10002
rect 14820 9900 14854 9934
rect 14820 9832 14854 9866
rect 14820 9764 14854 9798
rect 14820 9696 14854 9730
rect 14820 9628 14854 9662
rect 14820 9560 14854 9594
rect 14820 9492 14854 9526
rect 14820 9424 14854 9458
rect 14820 9356 14854 9390
rect 14820 9288 14854 9322
rect 14820 9220 14854 9254
rect 14820 9152 14854 9186
rect 14820 9084 14854 9118
rect 14820 9016 14854 9050
rect 14820 8948 14854 8982
rect 14820 8880 14854 8914
rect 14820 8812 14854 8846
rect 14820 8744 14854 8778
rect 14820 8676 14854 8710
rect 14820 8608 14854 8642
rect 14820 8540 14854 8574
rect 14820 8472 14854 8506
rect 14820 8404 14854 8438
rect 14820 8336 14854 8370
rect 14820 8268 14854 8302
rect 17204 11192 17238 11226
rect 17204 11124 17238 11158
rect 17204 11056 17238 11090
rect 17204 10988 17238 11022
rect 17204 10920 17238 10954
rect 17204 10852 17238 10886
rect 17204 10784 17238 10818
rect 17204 10716 17238 10750
rect 17204 10648 17238 10682
rect 17204 10580 17238 10614
rect 17204 10512 17238 10546
rect 17204 10444 17238 10478
rect 17204 10376 17238 10410
rect 17204 10308 17238 10342
rect 17204 10240 17238 10274
rect 17204 10172 17238 10206
rect 17204 10104 17238 10138
rect 17204 10036 17238 10070
rect 17204 9968 17238 10002
rect 17204 9900 17238 9934
rect 17204 9832 17238 9866
rect 17204 9764 17238 9798
rect 17204 9696 17238 9730
rect 17204 9628 17238 9662
rect 17204 9560 17238 9594
rect 17204 9492 17238 9526
rect 17204 9424 17238 9458
rect 17204 9356 17238 9390
rect 17204 9288 17238 9322
rect 17204 9220 17238 9254
rect 17204 9152 17238 9186
rect 17204 9084 17238 9118
rect 17204 9016 17238 9050
rect 17204 8948 17238 8982
rect 17204 8880 17238 8914
rect 17204 8812 17238 8846
rect 17204 8744 17238 8778
rect 17204 8676 17238 8710
rect 17204 8608 17238 8642
rect 17204 8540 17238 8574
rect 17204 8472 17238 8506
rect 17204 8404 17238 8438
rect 17204 8336 17238 8370
rect 17204 8268 17238 8302
rect 14820 8200 14854 8234
rect 14820 8132 14854 8166
rect 17204 8200 17238 8234
rect 17204 8132 17238 8166
rect 14924 8028 14958 8062
rect 14992 8028 15026 8062
rect 15060 8028 15094 8062
rect 15128 8028 15162 8062
rect 15196 8028 15230 8062
rect 15264 8028 15298 8062
rect 15332 8028 15366 8062
rect 15400 8028 15434 8062
rect 15468 8028 15502 8062
rect 15536 8028 15570 8062
rect 15604 8028 15638 8062
rect 15672 8028 15706 8062
rect 15740 8028 15774 8062
rect 15808 8028 15842 8062
rect 15876 8028 15910 8062
rect 15944 8028 15978 8062
rect 16012 8028 16046 8062
rect 16080 8028 16114 8062
rect 16148 8028 16182 8062
rect 16216 8028 16250 8062
rect 16284 8028 16318 8062
rect 16352 8028 16386 8062
rect 16420 8028 16454 8062
rect 16488 8028 16522 8062
rect 16556 8028 16590 8062
rect 16624 8028 16658 8062
rect 16692 8028 16726 8062
rect 16760 8028 16794 8062
rect 16828 8028 16862 8062
rect 16896 8028 16930 8062
rect 16964 8028 16998 8062
rect 17032 8028 17066 8062
rect 17100 8028 17134 8062
rect 17448 11406 17482 11440
rect 17516 11406 17550 11440
rect 17584 11406 17618 11440
rect 17652 11406 17686 11440
rect 17720 11406 17754 11440
rect 17788 11406 17822 11440
rect 17856 11406 17890 11440
rect 17924 11406 17958 11440
rect 17992 11406 18026 11440
rect 18060 11406 18094 11440
rect 18128 11406 18162 11440
rect 18196 11406 18230 11440
rect 18264 11406 18298 11440
rect 18332 11406 18366 11440
rect 18400 11406 18434 11440
rect 18468 11406 18502 11440
rect 18536 11406 18570 11440
rect 18604 11406 18638 11440
rect 18672 11406 18706 11440
rect 18740 11406 18774 11440
rect 18808 11406 18842 11440
rect 18876 11406 18910 11440
rect 18944 11406 18978 11440
rect 19012 11406 19046 11440
rect 19080 11406 19114 11440
rect 19148 11406 19182 11440
rect 19216 11406 19250 11440
rect 19284 11406 19318 11440
rect 19352 11406 19386 11440
rect 19420 11406 19454 11440
rect 19488 11406 19522 11440
rect 19556 11406 19590 11440
rect 19624 11406 19658 11440
rect 17344 11302 17378 11336
rect 17344 11234 17378 11268
rect 19728 11302 19762 11336
rect 19728 11234 19762 11268
rect 17344 11166 17378 11200
rect 17344 11098 17378 11132
rect 17344 11030 17378 11064
rect 17344 10962 17378 10996
rect 17344 10894 17378 10928
rect 17344 10826 17378 10860
rect 17344 10758 17378 10792
rect 17344 10690 17378 10724
rect 17344 10622 17378 10656
rect 17344 10554 17378 10588
rect 17344 10486 17378 10520
rect 17344 10418 17378 10452
rect 17344 10350 17378 10384
rect 17344 10282 17378 10316
rect 17344 10214 17378 10248
rect 17344 10146 17378 10180
rect 17344 10078 17378 10112
rect 17344 10010 17378 10044
rect 17344 9942 17378 9976
rect 17344 9874 17378 9908
rect 17344 9806 17378 9840
rect 17344 9738 17378 9772
rect 17344 9670 17378 9704
rect 17344 9602 17378 9636
rect 17344 9534 17378 9568
rect 17344 9466 17378 9500
rect 17344 9398 17378 9432
rect 17344 9330 17378 9364
rect 17344 9262 17378 9296
rect 17344 9194 17378 9228
rect 17344 9126 17378 9160
rect 17344 9058 17378 9092
rect 17344 8990 17378 9024
rect 17344 8922 17378 8956
rect 17344 8854 17378 8888
rect 17344 8786 17378 8820
rect 17344 8718 17378 8752
rect 17344 8650 17378 8684
rect 17344 8582 17378 8616
rect 17344 8514 17378 8548
rect 17344 8446 17378 8480
rect 17344 8378 17378 8412
rect 17344 8310 17378 8344
rect 17344 8242 17378 8276
rect 19728 11166 19762 11200
rect 19728 11098 19762 11132
rect 19728 11030 19762 11064
rect 19728 10962 19762 10996
rect 19728 10894 19762 10928
rect 19728 10826 19762 10860
rect 19728 10758 19762 10792
rect 19728 10690 19762 10724
rect 19728 10622 19762 10656
rect 19728 10554 19762 10588
rect 19728 10486 19762 10520
rect 19728 10418 19762 10452
rect 19728 10350 19762 10384
rect 19728 10282 19762 10316
rect 19728 10214 19762 10248
rect 19728 10146 19762 10180
rect 19728 10078 19762 10112
rect 19728 10010 19762 10044
rect 19728 9942 19762 9976
rect 19728 9874 19762 9908
rect 19728 9806 19762 9840
rect 19728 9738 19762 9772
rect 19728 9670 19762 9704
rect 19728 9602 19762 9636
rect 19728 9534 19762 9568
rect 19728 9466 19762 9500
rect 19728 9398 19762 9432
rect 19728 9330 19762 9364
rect 19728 9262 19762 9296
rect 19728 9194 19762 9228
rect 19728 9126 19762 9160
rect 19728 9058 19762 9092
rect 19728 8990 19762 9024
rect 19728 8922 19762 8956
rect 19728 8854 19762 8888
rect 19728 8786 19762 8820
rect 19728 8718 19762 8752
rect 19728 8650 19762 8684
rect 19728 8582 19762 8616
rect 19728 8514 19762 8548
rect 19728 8446 19762 8480
rect 19728 8378 19762 8412
rect 19728 8310 19762 8344
rect 19728 8242 19762 8276
rect 17344 8174 17378 8208
rect 17344 8106 17378 8140
rect 19728 8174 19762 8208
rect 19728 8106 19762 8140
rect 17448 8002 17482 8036
rect 17516 8002 17550 8036
rect 17584 8002 17618 8036
rect 17652 8002 17686 8036
rect 17720 8002 17754 8036
rect 17788 8002 17822 8036
rect 17856 8002 17890 8036
rect 17924 8002 17958 8036
rect 17992 8002 18026 8036
rect 18060 8002 18094 8036
rect 18128 8002 18162 8036
rect 18196 8002 18230 8036
rect 18264 8002 18298 8036
rect 18332 8002 18366 8036
rect 18400 8002 18434 8036
rect 18468 8002 18502 8036
rect 18536 8002 18570 8036
rect 18604 8002 18638 8036
rect 18672 8002 18706 8036
rect 18740 8002 18774 8036
rect 18808 8002 18842 8036
rect 18876 8002 18910 8036
rect 18944 8002 18978 8036
rect 19012 8002 19046 8036
rect 19080 8002 19114 8036
rect 19148 8002 19182 8036
rect 19216 8002 19250 8036
rect 19284 8002 19318 8036
rect 19352 8002 19386 8036
rect 19420 8002 19454 8036
rect 19488 8002 19522 8036
rect 19556 8002 19590 8036
rect 19624 8002 19658 8036
rect 23114 13456 23148 13490
rect 23182 13456 23216 13490
rect 23250 13456 23284 13490
rect 23318 13456 23352 13490
rect 23386 13456 23420 13490
rect 23454 13456 23488 13490
rect 23522 13456 23556 13490
rect 23590 13456 23624 13490
rect 23658 13456 23692 13490
rect 23726 13456 23760 13490
rect 23794 13456 23828 13490
rect 23862 13456 23896 13490
rect 23930 13456 23964 13490
rect 23998 13456 24032 13490
rect 24066 13456 24100 13490
rect 24134 13456 24168 13490
rect 24202 13456 24236 13490
rect 24270 13456 24304 13490
rect 22990 13337 23024 13371
rect 24394 13337 24428 13371
rect 22990 13269 23024 13303
rect 22990 13201 23024 13235
rect 22990 13133 23024 13167
rect 22990 13065 23024 13099
rect 22990 12997 23024 13031
rect 22990 12929 23024 12963
rect 22990 12861 23024 12895
rect 22990 12793 23024 12827
rect 22990 12725 23024 12759
rect 22990 12657 23024 12691
rect 22990 12589 23024 12623
rect 22990 12521 23024 12555
rect 22990 12453 23024 12487
rect 22990 12385 23024 12419
rect 22990 12317 23024 12351
rect 24394 13269 24428 13303
rect 24394 13201 24428 13235
rect 24394 13133 24428 13167
rect 24394 13065 24428 13099
rect 24394 12997 24428 13031
rect 24394 12929 24428 12963
rect 24394 12861 24428 12895
rect 24394 12793 24428 12827
rect 24394 12725 24428 12759
rect 24394 12657 24428 12691
rect 24394 12589 24428 12623
rect 24394 12521 24428 12555
rect 24394 12453 24428 12487
rect 24394 12385 24428 12419
rect 24394 12317 24428 12351
rect 22990 12249 23024 12283
rect 24394 12249 24428 12283
rect 23114 12130 23148 12164
rect 23182 12130 23216 12164
rect 23250 12130 23284 12164
rect 23318 12130 23352 12164
rect 23386 12130 23420 12164
rect 23454 12130 23488 12164
rect 23522 12130 23556 12164
rect 23590 12130 23624 12164
rect 23658 12130 23692 12164
rect 23726 12130 23760 12164
rect 23794 12130 23828 12164
rect 23862 12130 23896 12164
rect 23930 12130 23964 12164
rect 23998 12130 24032 12164
rect 24066 12130 24100 12164
rect 24134 12130 24168 12164
rect 24202 12130 24236 12164
rect 24270 12130 24304 12164
rect 24674 13450 24708 13484
rect 24742 13450 24776 13484
rect 24810 13450 24844 13484
rect 24878 13450 24912 13484
rect 24946 13450 24980 13484
rect 25014 13450 25048 13484
rect 25082 13450 25116 13484
rect 25150 13450 25184 13484
rect 25218 13450 25252 13484
rect 25286 13450 25320 13484
rect 25354 13450 25388 13484
rect 25422 13450 25456 13484
rect 25490 13450 25524 13484
rect 25558 13450 25592 13484
rect 25626 13450 25660 13484
rect 25694 13450 25728 13484
rect 25762 13450 25796 13484
rect 25830 13450 25864 13484
rect 24550 13342 24584 13376
rect 24550 13274 24584 13308
rect 25954 13342 25988 13376
rect 24550 13206 24584 13240
rect 24550 13138 24584 13172
rect 24550 13070 24584 13104
rect 24550 13002 24584 13036
rect 24550 12934 24584 12968
rect 24550 12866 24584 12900
rect 24550 12798 24584 12832
rect 24550 12730 24584 12764
rect 24550 12662 24584 12696
rect 24550 12594 24584 12628
rect 24550 12526 24584 12560
rect 24550 12458 24584 12492
rect 24550 12390 24584 12424
rect 24550 12322 24584 12356
rect 25954 13274 25988 13308
rect 25954 13206 25988 13240
rect 25954 13138 25988 13172
rect 25954 13070 25988 13104
rect 25954 13002 25988 13036
rect 25954 12934 25988 12968
rect 25954 12866 25988 12900
rect 25954 12798 25988 12832
rect 25954 12730 25988 12764
rect 25954 12662 25988 12696
rect 25954 12594 25988 12628
rect 25954 12526 25988 12560
rect 25954 12458 25988 12492
rect 25954 12390 25988 12424
rect 25954 12322 25988 12356
rect 24550 12254 24584 12288
rect 25954 12254 25988 12288
rect 24550 12186 24584 12220
rect 24550 12118 24584 12152
rect 24550 12050 24584 12084
rect 24550 11982 24584 12016
rect 24550 11914 24584 11948
rect 24550 11846 24584 11880
rect 24550 11778 24584 11812
rect 24550 11710 24584 11744
rect 24550 11642 24584 11676
rect 24550 11574 24584 11608
rect 24550 11506 24584 11540
rect 24550 11438 24584 11472
rect 24550 11370 24584 11404
rect 24550 11302 24584 11336
rect 24550 11234 24584 11268
rect 25954 12186 25988 12220
rect 25954 12118 25988 12152
rect 25954 12050 25988 12084
rect 25954 11982 25988 12016
rect 25954 11914 25988 11948
rect 25954 11846 25988 11880
rect 25954 11778 25988 11812
rect 25954 11710 25988 11744
rect 25954 11642 25988 11676
rect 25954 11574 25988 11608
rect 25954 11506 25988 11540
rect 25954 11438 25988 11472
rect 25954 11370 25988 11404
rect 25954 11302 25988 11336
rect 24550 11166 24584 11200
rect 25954 11234 25988 11268
rect 24550 11098 24584 11132
rect 24550 11030 24584 11064
rect 24550 10962 24584 10996
rect 24550 10894 24584 10928
rect 24550 10826 24584 10860
rect 24550 10758 24584 10792
rect 24550 10690 24584 10724
rect 24550 10622 24584 10656
rect 24550 10554 24584 10588
rect 24550 10486 24584 10520
rect 24550 10418 24584 10452
rect 24550 10350 24584 10384
rect 24550 10282 24584 10316
rect 24550 10214 24584 10248
rect 25954 11166 25988 11200
rect 25954 11098 25988 11132
rect 25954 11030 25988 11064
rect 25954 10962 25988 10996
rect 25954 10894 25988 10928
rect 25954 10826 25988 10860
rect 25954 10758 25988 10792
rect 25954 10690 25988 10724
rect 25954 10622 25988 10656
rect 25954 10554 25988 10588
rect 25954 10486 25988 10520
rect 25954 10418 25988 10452
rect 25954 10350 25988 10384
rect 25954 10282 25988 10316
rect 25954 10214 25988 10248
rect 24550 10146 24584 10180
rect 25954 10146 25988 10180
rect 24550 10078 24584 10112
rect 24550 10010 24584 10044
rect 24550 9942 24584 9976
rect 24550 9874 24584 9908
rect 24550 9806 24584 9840
rect 24550 9738 24584 9772
rect 24550 9670 24584 9704
rect 24550 9602 24584 9636
rect 24550 9534 24584 9568
rect 24550 9466 24584 9500
rect 24550 9398 24584 9432
rect 24550 9330 24584 9364
rect 24550 9262 24584 9296
rect 24550 9194 24584 9228
rect 24550 9126 24584 9160
rect 25954 10078 25988 10112
rect 25954 10010 25988 10044
rect 25954 9942 25988 9976
rect 25954 9874 25988 9908
rect 25954 9806 25988 9840
rect 25954 9738 25988 9772
rect 25954 9670 25988 9704
rect 25954 9602 25988 9636
rect 25954 9534 25988 9568
rect 25954 9466 25988 9500
rect 25954 9398 25988 9432
rect 25954 9330 25988 9364
rect 25954 9262 25988 9296
rect 25954 9194 25988 9228
rect 24550 9058 24584 9092
rect 25954 9126 25988 9160
rect 25954 9058 25988 9092
rect 24674 8950 24708 8984
rect 24742 8950 24776 8984
rect 24810 8950 24844 8984
rect 24878 8950 24912 8984
rect 24946 8950 24980 8984
rect 25014 8950 25048 8984
rect 25082 8950 25116 8984
rect 25150 8950 25184 8984
rect 25218 8950 25252 8984
rect 25286 8950 25320 8984
rect 25354 8950 25388 8984
rect 25422 8950 25456 8984
rect 25490 8950 25524 8984
rect 25558 8950 25592 8984
rect 25626 8950 25660 8984
rect 25694 8950 25728 8984
rect 25762 8950 25796 8984
rect 25830 8950 25864 8984
<< poly >>
rect 23222 18828 24222 18844
rect 23222 18794 23263 18828
rect 23297 18794 23331 18828
rect 23365 18794 23399 18828
rect 23433 18794 23467 18828
rect 23501 18794 23535 18828
rect 23569 18794 23603 18828
rect 23637 18794 23671 18828
rect 23705 18794 23739 18828
rect 23773 18794 23807 18828
rect 23841 18794 23875 18828
rect 23909 18794 23943 18828
rect 23977 18794 24011 18828
rect 24045 18794 24079 18828
rect 24113 18794 24147 18828
rect 24181 18794 24222 18828
rect 23222 18747 24222 18794
rect -2934 18174 -2734 18190
rect -2934 18140 -2885 18174
rect -2851 18140 -2817 18174
rect -2783 18140 -2734 18174
rect -2934 18093 -2734 18140
rect -2676 18174 -2476 18190
rect -2676 18140 -2627 18174
rect -2593 18140 -2559 18174
rect -2525 18140 -2476 18174
rect -2676 18093 -2476 18140
rect -2418 18174 -2218 18190
rect -2418 18140 -2369 18174
rect -2335 18140 -2301 18174
rect -2267 18140 -2218 18174
rect -2418 18093 -2218 18140
rect -2160 18174 -1960 18190
rect -2160 18140 -2111 18174
rect -2077 18140 -2043 18174
rect -2009 18140 -1960 18174
rect -2160 18093 -1960 18140
rect -1902 18174 -1702 18190
rect -1902 18140 -1853 18174
rect -1819 18140 -1785 18174
rect -1751 18140 -1702 18174
rect -1902 18093 -1702 18140
rect -1644 18174 -1444 18190
rect -1644 18140 -1595 18174
rect -1561 18140 -1527 18174
rect -1493 18140 -1444 18174
rect -1644 18093 -1444 18140
rect -1386 18174 -1186 18190
rect -1386 18140 -1337 18174
rect -1303 18140 -1269 18174
rect -1235 18140 -1186 18174
rect -1386 18093 -1186 18140
rect -1128 18174 -928 18190
rect -1128 18140 -1079 18174
rect -1045 18140 -1011 18174
rect -977 18140 -928 18174
rect -1128 18093 -928 18140
rect -870 18174 -670 18190
rect -870 18140 -821 18174
rect -787 18140 -753 18174
rect -719 18140 -670 18174
rect -870 18093 -670 18140
rect -612 18174 -412 18190
rect -612 18140 -563 18174
rect -529 18140 -495 18174
rect -461 18140 -412 18174
rect -612 18093 -412 18140
rect -6402 17305 -6202 17321
rect -6402 17271 -6353 17305
rect -6319 17271 -6285 17305
rect -6251 17271 -6202 17305
rect -6402 17224 -6202 17271
rect -6144 17305 -5944 17321
rect -6144 17271 -6095 17305
rect -6061 17271 -6027 17305
rect -5993 17271 -5944 17305
rect -6144 17224 -5944 17271
rect -6402 16177 -6202 16224
rect -6402 16143 -6353 16177
rect -6319 16143 -6285 16177
rect -6251 16143 -6202 16177
rect -6402 16127 -6202 16143
rect -6144 16177 -5944 16224
rect -6144 16143 -6095 16177
rect -6061 16143 -6027 16177
rect -5993 16143 -5944 16177
rect -6144 16127 -5944 16143
rect 23222 17700 24222 17747
rect 23222 17666 23263 17700
rect 23297 17666 23331 17700
rect 23365 17666 23399 17700
rect 23433 17666 23467 17700
rect 23501 17666 23535 17700
rect 23569 17666 23603 17700
rect 23637 17666 23671 17700
rect 23705 17666 23739 17700
rect 23773 17666 23807 17700
rect 23841 17666 23875 17700
rect 23909 17666 23943 17700
rect 23977 17666 24011 17700
rect 24045 17666 24079 17700
rect 24113 17666 24147 17700
rect 24181 17666 24222 17700
rect 23222 17650 24222 17666
rect 24738 18828 25738 18844
rect 24738 18794 24779 18828
rect 24813 18794 24847 18828
rect 24881 18794 24915 18828
rect 24949 18794 24983 18828
rect 25017 18794 25051 18828
rect 25085 18794 25119 18828
rect 25153 18794 25187 18828
rect 25221 18794 25255 18828
rect 25289 18794 25323 18828
rect 25357 18794 25391 18828
rect 25425 18794 25459 18828
rect 25493 18794 25527 18828
rect 25561 18794 25595 18828
rect 25629 18794 25663 18828
rect 25697 18794 25738 18828
rect 24738 18747 25738 18794
rect 25796 18828 26796 18844
rect 25796 18794 25837 18828
rect 25871 18794 25905 18828
rect 25939 18794 25973 18828
rect 26007 18794 26041 18828
rect 26075 18794 26109 18828
rect 26143 18794 26177 18828
rect 26211 18794 26245 18828
rect 26279 18794 26313 18828
rect 26347 18794 26381 18828
rect 26415 18794 26449 18828
rect 26483 18794 26517 18828
rect 26551 18794 26585 18828
rect 26619 18794 26653 18828
rect 26687 18794 26721 18828
rect 26755 18794 26796 18828
rect 25796 18747 26796 18794
rect 26854 18828 27854 18844
rect 26854 18794 26895 18828
rect 26929 18794 26963 18828
rect 26997 18794 27031 18828
rect 27065 18794 27099 18828
rect 27133 18794 27167 18828
rect 27201 18794 27235 18828
rect 27269 18794 27303 18828
rect 27337 18794 27371 18828
rect 27405 18794 27439 18828
rect 27473 18794 27507 18828
rect 27541 18794 27575 18828
rect 27609 18794 27643 18828
rect 27677 18794 27711 18828
rect 27745 18794 27779 18828
rect 27813 18794 27854 18828
rect 26854 18747 27854 18794
rect -2934 16046 -2734 16093
rect -2934 16012 -2885 16046
rect -2851 16012 -2817 16046
rect -2783 16012 -2734 16046
rect -2934 15996 -2734 16012
rect -2676 16046 -2476 16093
rect -2676 16012 -2627 16046
rect -2593 16012 -2559 16046
rect -2525 16012 -2476 16046
rect -2676 15996 -2476 16012
rect -2418 16046 -2218 16093
rect -2418 16012 -2369 16046
rect -2335 16012 -2301 16046
rect -2267 16012 -2218 16046
rect -2418 15996 -2218 16012
rect -2160 16046 -1960 16093
rect -2160 16012 -2111 16046
rect -2077 16012 -2043 16046
rect -2009 16012 -1960 16046
rect -2160 15996 -1960 16012
rect -1902 16046 -1702 16093
rect -1902 16012 -1853 16046
rect -1819 16012 -1785 16046
rect -1751 16012 -1702 16046
rect -1902 15996 -1702 16012
rect -1644 16046 -1444 16093
rect -1644 16012 -1595 16046
rect -1561 16012 -1527 16046
rect -1493 16012 -1444 16046
rect -1644 15996 -1444 16012
rect -1386 16046 -1186 16093
rect -1386 16012 -1337 16046
rect -1303 16012 -1269 16046
rect -1235 16012 -1186 16046
rect -1386 15996 -1186 16012
rect -1128 16046 -928 16093
rect -1128 16012 -1079 16046
rect -1045 16012 -1011 16046
rect -977 16012 -928 16046
rect -1128 15996 -928 16012
rect -870 16046 -670 16093
rect -870 16012 -821 16046
rect -787 16012 -753 16046
rect -719 16012 -670 16046
rect -870 15996 -670 16012
rect -612 16046 -412 16093
rect -612 16012 -563 16046
rect -529 16012 -495 16046
rect -461 16012 -412 16046
rect -612 15996 -412 16012
rect 23196 17208 24196 17224
rect 23196 17174 23237 17208
rect 23271 17174 23305 17208
rect 23339 17174 23373 17208
rect 23407 17174 23441 17208
rect 23475 17174 23509 17208
rect 23543 17174 23577 17208
rect 23611 17174 23645 17208
rect 23679 17174 23713 17208
rect 23747 17174 23781 17208
rect 23815 17174 23849 17208
rect 23883 17174 23917 17208
rect 23951 17174 23985 17208
rect 24019 17174 24053 17208
rect 24087 17174 24121 17208
rect 24155 17174 24196 17208
rect 23196 17136 24196 17174
rect 42658 18924 42858 18940
rect 42658 18890 42707 18924
rect 42741 18890 42775 18924
rect 42809 18890 42858 18924
rect 42658 18843 42858 18890
rect 42916 18924 43116 18940
rect 42916 18890 42965 18924
rect 42999 18890 43033 18924
rect 43067 18890 43116 18924
rect 42916 18843 43116 18890
rect 43174 18924 43374 18940
rect 43174 18890 43223 18924
rect 43257 18890 43291 18924
rect 43325 18890 43374 18924
rect 43174 18843 43374 18890
rect 43432 18924 43632 18940
rect 43432 18890 43481 18924
rect 43515 18890 43549 18924
rect 43583 18890 43632 18924
rect 43432 18843 43632 18890
rect 43690 18924 43890 18940
rect 43690 18890 43739 18924
rect 43773 18890 43807 18924
rect 43841 18890 43890 18924
rect 43690 18843 43890 18890
rect 43948 18924 44148 18940
rect 43948 18890 43997 18924
rect 44031 18890 44065 18924
rect 44099 18890 44148 18924
rect 43948 18843 44148 18890
rect 44206 18924 44406 18940
rect 44206 18890 44255 18924
rect 44289 18890 44323 18924
rect 44357 18890 44406 18924
rect 44206 18843 44406 18890
rect 44464 18924 44664 18940
rect 44464 18890 44513 18924
rect 44547 18890 44581 18924
rect 44615 18890 44664 18924
rect 44464 18843 44664 18890
rect 44722 18924 44922 18940
rect 44722 18890 44771 18924
rect 44805 18890 44839 18924
rect 44873 18890 44922 18924
rect 44722 18843 44922 18890
rect 44980 18924 45180 18940
rect 44980 18890 45029 18924
rect 45063 18890 45097 18924
rect 45131 18890 45180 18924
rect 44980 18843 45180 18890
rect 24738 17100 25738 17147
rect 24738 17066 24779 17100
rect 24813 17066 24847 17100
rect 24881 17066 24915 17100
rect 24949 17066 24983 17100
rect 25017 17066 25051 17100
rect 25085 17066 25119 17100
rect 25153 17066 25187 17100
rect 25221 17066 25255 17100
rect 25289 17066 25323 17100
rect 25357 17066 25391 17100
rect 25425 17066 25459 17100
rect 25493 17066 25527 17100
rect 25561 17066 25595 17100
rect 25629 17066 25663 17100
rect 25697 17066 25738 17100
rect 24738 17050 25738 17066
rect 25796 17100 26796 17147
rect 25796 17066 25837 17100
rect 25871 17066 25905 17100
rect 25939 17066 25973 17100
rect 26007 17066 26041 17100
rect 26075 17066 26109 17100
rect 26143 17066 26177 17100
rect 26211 17066 26245 17100
rect 26279 17066 26313 17100
rect 26347 17066 26381 17100
rect 26415 17066 26449 17100
rect 26483 17066 26517 17100
rect 26551 17066 26585 17100
rect 26619 17066 26653 17100
rect 26687 17066 26721 17100
rect 26755 17066 26796 17100
rect 25796 17050 26796 17066
rect 26854 17100 27854 17147
rect 26854 17066 26895 17100
rect 26929 17066 26963 17100
rect 26997 17066 27031 17100
rect 27065 17066 27099 17100
rect 27133 17066 27167 17100
rect 27201 17066 27235 17100
rect 27269 17066 27303 17100
rect 27337 17066 27371 17100
rect 27405 17066 27439 17100
rect 27473 17066 27507 17100
rect 27541 17066 27575 17100
rect 27609 17066 27643 17100
rect 27677 17066 27711 17100
rect 27745 17066 27779 17100
rect 27813 17066 27854 17100
rect 26854 17050 27854 17066
rect 39190 18055 39390 18071
rect 39190 18021 39239 18055
rect 39273 18021 39307 18055
rect 39341 18021 39390 18055
rect 39190 17974 39390 18021
rect 39448 18055 39648 18071
rect 39448 18021 39497 18055
rect 39531 18021 39565 18055
rect 39599 18021 39648 18055
rect 39448 17974 39648 18021
rect 39190 16927 39390 16974
rect 39190 16893 39239 16927
rect 39273 16893 39307 16927
rect 39341 16893 39390 16927
rect 39190 16877 39390 16893
rect 39448 16927 39648 16974
rect 39448 16893 39497 16927
rect 39531 16893 39565 16927
rect 39599 16893 39648 16927
rect 39448 16877 39648 16893
rect 23196 16098 24196 16136
rect 23196 16064 23237 16098
rect 23271 16064 23305 16098
rect 23339 16064 23373 16098
rect 23407 16064 23441 16098
rect 23475 16064 23509 16098
rect 23543 16064 23577 16098
rect 23611 16064 23645 16098
rect 23679 16064 23713 16098
rect 23747 16064 23781 16098
rect 23815 16064 23849 16098
rect 23883 16064 23917 16098
rect 23951 16064 23985 16098
rect 24019 16064 24053 16098
rect 24087 16064 24121 16098
rect 24155 16064 24196 16098
rect 23196 16048 24196 16064
rect 42658 16796 42858 16843
rect 42658 16762 42707 16796
rect 42741 16762 42775 16796
rect 42809 16762 42858 16796
rect 42658 16746 42858 16762
rect 42916 16796 43116 16843
rect 42916 16762 42965 16796
rect 42999 16762 43033 16796
rect 43067 16762 43116 16796
rect 42916 16746 43116 16762
rect 43174 16796 43374 16843
rect 43174 16762 43223 16796
rect 43257 16762 43291 16796
rect 43325 16762 43374 16796
rect 43174 16746 43374 16762
rect 43432 16796 43632 16843
rect 43432 16762 43481 16796
rect 43515 16762 43549 16796
rect 43583 16762 43632 16796
rect 43432 16746 43632 16762
rect 43690 16796 43890 16843
rect 43690 16762 43739 16796
rect 43773 16762 43807 16796
rect 43841 16762 43890 16796
rect 43690 16746 43890 16762
rect 43948 16796 44148 16843
rect 43948 16762 43997 16796
rect 44031 16762 44065 16796
rect 44099 16762 44148 16796
rect 43948 16746 44148 16762
rect 44206 16796 44406 16843
rect 44206 16762 44255 16796
rect 44289 16762 44323 16796
rect 44357 16762 44406 16796
rect 44206 16746 44406 16762
rect 44464 16796 44664 16843
rect 44464 16762 44513 16796
rect 44547 16762 44581 16796
rect 44615 16762 44664 16796
rect 44464 16746 44664 16762
rect 44722 16796 44922 16843
rect 44722 16762 44771 16796
rect 44805 16762 44839 16796
rect 44873 16762 44922 16796
rect 44722 16746 44922 16762
rect 44980 16796 45180 16843
rect 44980 16762 45029 16796
rect 45063 16762 45097 16796
rect 45131 16762 45180 16796
rect 44980 16746 45180 16762
rect -7136 14968 -6973 14998
rect -7136 14934 -7080 14968
rect -7046 14934 -6973 14968
rect -7136 14861 -6973 14934
rect -6878 14968 -6715 14996
rect -6878 14934 -6820 14968
rect -6786 14934 -6715 14968
rect -6878 14861 -6715 14934
rect -6097 14957 -5944 14982
rect -6097 14923 -6028 14957
rect -5994 14923 -5944 14957
rect -6097 14861 -5944 14923
rect -5844 14944 -5691 14982
rect -5844 14910 -5778 14944
rect -5744 14910 -5691 14944
rect -5844 14861 -5691 14910
rect -5060 14948 -4921 14982
rect -5060 14914 -5007 14948
rect -4973 14914 -4921 14948
rect -5060 14861 -4921 14914
rect -7413 14835 -7213 14861
rect -7155 14835 -6955 14861
rect -6897 14835 -6697 14861
rect -6639 14835 -6439 14861
rect -6381 14835 -6181 14861
rect -6123 14835 -5923 14861
rect -5865 14835 -5665 14861
rect -5607 14835 -5407 14861
rect -5349 14835 -5149 14861
rect -5091 14835 -4891 14861
rect -7413 12809 -7213 12835
rect -7155 12809 -6955 12835
rect -6897 12809 -6697 12835
rect -6639 12809 -6439 12835
rect -6381 12809 -6181 12835
rect -6123 12809 -5923 12835
rect -5865 12809 -5665 12835
rect -5607 12809 -5407 12835
rect -5349 12809 -5149 12835
rect -5091 12809 -4891 12835
rect -7392 12721 -7246 12809
rect -7392 12687 -7343 12721
rect -7309 12687 -7246 12721
rect -7392 12674 -7246 12687
rect -6617 12729 -6457 12809
rect -6617 12695 -6547 12729
rect -6513 12695 -6457 12729
rect -7392 12640 -7232 12674
rect -6617 12649 -6457 12695
rect -6359 12724 -6199 12809
rect -6359 12690 -6310 12724
rect -6276 12690 -6199 12724
rect -6359 12645 -6199 12690
rect -5586 12726 -5426 12809
rect -5586 12692 -5516 12726
rect -5482 12692 -5426 12726
rect -5586 12646 -5426 12692
rect -5328 12726 -5168 12809
rect -5328 12692 -5261 12726
rect -5227 12692 -5168 12726
rect -5328 12646 -5168 12692
rect 13040 14848 14040 14864
rect 13040 14814 13081 14848
rect 13115 14814 13149 14848
rect 13183 14814 13217 14848
rect 13251 14814 13285 14848
rect 13319 14814 13353 14848
rect 13387 14814 13421 14848
rect 13455 14814 13489 14848
rect 13523 14814 13557 14848
rect 13591 14814 13625 14848
rect 13659 14814 13693 14848
rect 13727 14814 13761 14848
rect 13795 14814 13829 14848
rect 13863 14814 13897 14848
rect 13931 14814 13965 14848
rect 13999 14814 14040 14848
rect 13040 14767 14040 14814
rect 14098 14848 15098 14864
rect 14098 14814 14139 14848
rect 14173 14814 14207 14848
rect 14241 14814 14275 14848
rect 14309 14814 14343 14848
rect 14377 14814 14411 14848
rect 14445 14814 14479 14848
rect 14513 14814 14547 14848
rect 14581 14814 14615 14848
rect 14649 14814 14683 14848
rect 14717 14814 14751 14848
rect 14785 14814 14819 14848
rect 14853 14814 14887 14848
rect 14921 14814 14955 14848
rect 14989 14814 15023 14848
rect 15057 14814 15098 14848
rect 14098 14767 15098 14814
rect 13040 11720 14040 11767
rect 13040 11686 13081 11720
rect 13115 11686 13149 11720
rect 13183 11686 13217 11720
rect 13251 11686 13285 11720
rect 13319 11686 13353 11720
rect 13387 11686 13421 11720
rect 13455 11686 13489 11720
rect 13523 11686 13557 11720
rect 13591 11686 13625 11720
rect 13659 11686 13693 11720
rect 13727 11686 13761 11720
rect 13795 11686 13829 11720
rect 13863 11686 13897 11720
rect 13931 11686 13965 11720
rect 13999 11686 14040 11720
rect 13040 11670 14040 11686
rect 14098 11720 15098 11767
rect 14098 11686 14139 11720
rect 14173 11686 14207 11720
rect 14241 11686 14275 11720
rect 14309 11686 14343 11720
rect 14377 11686 14411 11720
rect 14445 11686 14479 11720
rect 14513 11686 14547 11720
rect 14581 11686 14615 11720
rect 14649 11686 14683 11720
rect 14717 11686 14751 11720
rect 14785 11686 14819 11720
rect 14853 11686 14887 11720
rect 14921 11686 14955 11720
rect 14989 11686 15023 11720
rect 15057 11686 15098 11720
rect 14098 11670 15098 11686
rect 15610 14848 16610 14864
rect 15610 14814 15651 14848
rect 15685 14814 15719 14848
rect 15753 14814 15787 14848
rect 15821 14814 15855 14848
rect 15889 14814 15923 14848
rect 15957 14814 15991 14848
rect 16025 14814 16059 14848
rect 16093 14814 16127 14848
rect 16161 14814 16195 14848
rect 16229 14814 16263 14848
rect 16297 14814 16331 14848
rect 16365 14814 16399 14848
rect 16433 14814 16467 14848
rect 16501 14814 16535 14848
rect 16569 14814 16610 14848
rect 15610 14767 16610 14814
rect 15610 11720 16610 11767
rect 15610 11686 15651 11720
rect 15685 11686 15719 11720
rect 15753 11686 15787 11720
rect 15821 11686 15855 11720
rect 15889 11686 15923 11720
rect 15957 11686 15991 11720
rect 16025 11686 16059 11720
rect 16093 11686 16127 11720
rect 16161 11686 16195 11720
rect 16229 11686 16263 11720
rect 16297 11686 16331 11720
rect 16365 11686 16399 11720
rect 16433 11686 16467 11720
rect 16501 11686 16535 11720
rect 16569 11686 16610 11720
rect 15610 11670 16610 11686
rect 17120 14858 18120 14874
rect 17120 14824 17161 14858
rect 17195 14824 17229 14858
rect 17263 14824 17297 14858
rect 17331 14824 17365 14858
rect 17399 14824 17433 14858
rect 17467 14824 17501 14858
rect 17535 14824 17569 14858
rect 17603 14824 17637 14858
rect 17671 14824 17705 14858
rect 17739 14824 17773 14858
rect 17807 14824 17841 14858
rect 17875 14824 17909 14858
rect 17943 14824 17977 14858
rect 18011 14824 18045 14858
rect 18079 14824 18120 14858
rect 17120 14777 18120 14824
rect 17120 11730 18120 11777
rect 17120 11696 17161 11730
rect 17195 11696 17229 11730
rect 17263 11696 17297 11730
rect 17331 11696 17365 11730
rect 17399 11696 17433 11730
rect 17467 11696 17501 11730
rect 17535 11696 17569 11730
rect 17603 11696 17637 11730
rect 17671 11696 17705 11730
rect 17739 11696 17773 11730
rect 17807 11696 17841 11730
rect 17875 11696 17909 11730
rect 17943 11696 17977 11730
rect 18011 11696 18045 11730
rect 18079 11696 18120 11730
rect 17120 11680 18120 11696
rect 18584 14842 19584 14858
rect 18584 14808 18625 14842
rect 18659 14808 18693 14842
rect 18727 14808 18761 14842
rect 18795 14808 18829 14842
rect 18863 14808 18897 14842
rect 18931 14808 18965 14842
rect 18999 14808 19033 14842
rect 19067 14808 19101 14842
rect 19135 14808 19169 14842
rect 19203 14808 19237 14842
rect 19271 14808 19305 14842
rect 19339 14808 19373 14842
rect 19407 14808 19441 14842
rect 19475 14808 19509 14842
rect 19543 14808 19584 14842
rect 18584 14761 19584 14808
rect 38456 15718 38619 15748
rect 38456 15684 38512 15718
rect 38546 15684 38619 15718
rect 38456 15611 38619 15684
rect 38714 15718 38877 15746
rect 38714 15684 38772 15718
rect 38806 15684 38877 15718
rect 38714 15611 38877 15684
rect 39495 15707 39648 15732
rect 39495 15673 39564 15707
rect 39598 15673 39648 15707
rect 39495 15611 39648 15673
rect 39748 15694 39901 15732
rect 39748 15660 39814 15694
rect 39848 15660 39901 15694
rect 39748 15611 39901 15660
rect 40532 15698 40671 15732
rect 40532 15664 40585 15698
rect 40619 15664 40671 15698
rect 40532 15611 40671 15664
rect 38179 15585 38379 15611
rect 38437 15585 38637 15611
rect 38695 15585 38895 15611
rect 38953 15585 39153 15611
rect 39211 15585 39411 15611
rect 39469 15585 39669 15611
rect 39727 15585 39927 15611
rect 39985 15585 40185 15611
rect 40243 15585 40443 15611
rect 40501 15585 40701 15611
rect 18584 11714 19584 11761
rect 18584 11680 18625 11714
rect 18659 11680 18693 11714
rect 18727 11680 18761 11714
rect 18795 11680 18829 11714
rect 18863 11680 18897 11714
rect 18931 11680 18965 11714
rect 18999 11680 19033 11714
rect 19067 11680 19101 11714
rect 19135 11680 19169 11714
rect 19203 11680 19237 11714
rect 19271 11680 19305 11714
rect 19339 11680 19373 11714
rect 19407 11680 19441 11714
rect 19475 11680 19509 11714
rect 19543 11680 19584 11714
rect 18584 11664 19584 11680
rect -8769 11236 -8569 11252
rect -8769 11202 -8720 11236
rect -8686 11202 -8652 11236
rect -8618 11202 -8569 11236
rect -8769 11164 -8569 11202
rect -8511 11236 -8311 11252
rect -8511 11202 -8462 11236
rect -8428 11202 -8394 11236
rect -8360 11202 -8311 11236
rect -8511 11164 -8311 11202
rect -8253 11236 -8053 11252
rect -8253 11202 -8204 11236
rect -8170 11202 -8136 11236
rect -8102 11202 -8053 11236
rect -8253 11164 -8053 11202
rect -7995 11236 -7795 11252
rect -7995 11202 -7946 11236
rect -7912 11202 -7878 11236
rect -7844 11202 -7795 11236
rect -7995 11164 -7795 11202
rect -7737 11236 -7537 11252
rect -7737 11202 -7688 11236
rect -7654 11202 -7620 11236
rect -7586 11202 -7537 11236
rect -7737 11164 -7537 11202
rect -7479 11236 -7279 11252
rect -7479 11202 -7430 11236
rect -7396 11202 -7362 11236
rect -7328 11202 -7279 11236
rect -7479 11164 -7279 11202
rect -7221 11236 -7021 11252
rect -7221 11202 -7172 11236
rect -7138 11202 -7104 11236
rect -7070 11202 -7021 11236
rect -7221 11164 -7021 11202
rect -6963 11236 -6763 11252
rect -6963 11202 -6914 11236
rect -6880 11202 -6846 11236
rect -6812 11202 -6763 11236
rect -6963 11164 -6763 11202
rect -6705 11236 -6505 11252
rect -6705 11202 -6656 11236
rect -6622 11202 -6588 11236
rect -6554 11202 -6505 11236
rect -6705 11164 -6505 11202
rect -6447 11236 -6247 11252
rect -6447 11202 -6398 11236
rect -6364 11202 -6330 11236
rect -6296 11202 -6247 11236
rect -6447 11164 -6247 11202
rect -6189 11236 -5989 11252
rect -6189 11202 -6140 11236
rect -6106 11202 -6072 11236
rect -6038 11202 -5989 11236
rect -6189 11164 -5989 11202
rect -5931 11236 -5731 11252
rect -5931 11202 -5882 11236
rect -5848 11202 -5814 11236
rect -5780 11202 -5731 11236
rect -5931 11164 -5731 11202
rect -5673 11236 -5473 11252
rect -5673 11202 -5624 11236
rect -5590 11202 -5556 11236
rect -5522 11202 -5473 11236
rect -5673 11164 -5473 11202
rect -5415 11236 -5215 11252
rect -5415 11202 -5366 11236
rect -5332 11202 -5298 11236
rect -5264 11202 -5215 11236
rect -5415 11164 -5215 11202
rect -5157 11236 -4957 11252
rect -5157 11202 -5108 11236
rect -5074 11202 -5040 11236
rect -5006 11202 -4957 11236
rect -5157 11164 -4957 11202
rect -4899 11236 -4699 11252
rect -4899 11202 -4850 11236
rect -4816 11202 -4782 11236
rect -4748 11202 -4699 11236
rect -4899 11164 -4699 11202
rect -4641 11236 -4441 11252
rect -4641 11202 -4592 11236
rect -4558 11202 -4524 11236
rect -4490 11202 -4441 11236
rect -4641 11164 -4441 11202
rect -4383 11236 -4183 11252
rect -4383 11202 -4334 11236
rect -4300 11202 -4266 11236
rect -4232 11202 -4183 11236
rect -4383 11164 -4183 11202
rect -4125 11236 -3925 11252
rect -4125 11202 -4076 11236
rect -4042 11202 -4008 11236
rect -3974 11202 -3925 11236
rect -4125 11164 -3925 11202
rect -3867 11236 -3667 11252
rect -3867 11202 -3818 11236
rect -3784 11202 -3750 11236
rect -3716 11202 -3667 11236
rect -3867 11164 -3667 11202
rect -8769 10126 -8569 10164
rect -8769 10092 -8720 10126
rect -8686 10092 -8652 10126
rect -8618 10092 -8569 10126
rect -8769 10076 -8569 10092
rect -8511 10126 -8311 10164
rect -8511 10092 -8462 10126
rect -8428 10092 -8394 10126
rect -8360 10092 -8311 10126
rect -8511 10076 -8311 10092
rect -8253 10126 -8053 10164
rect -8253 10092 -8204 10126
rect -8170 10092 -8136 10126
rect -8102 10092 -8053 10126
rect -8253 10076 -8053 10092
rect -7995 10126 -7795 10164
rect -7995 10092 -7946 10126
rect -7912 10092 -7878 10126
rect -7844 10092 -7795 10126
rect -7995 10076 -7795 10092
rect -7737 10126 -7537 10164
rect -7737 10092 -7688 10126
rect -7654 10092 -7620 10126
rect -7586 10092 -7537 10126
rect -7737 10076 -7537 10092
rect -7479 10126 -7279 10164
rect -7479 10092 -7430 10126
rect -7396 10092 -7362 10126
rect -7328 10092 -7279 10126
rect -7479 10076 -7279 10092
rect -7221 10126 -7021 10164
rect -7221 10092 -7172 10126
rect -7138 10092 -7104 10126
rect -7070 10092 -7021 10126
rect -7221 10076 -7021 10092
rect -6963 10126 -6763 10164
rect -6963 10092 -6914 10126
rect -6880 10092 -6846 10126
rect -6812 10092 -6763 10126
rect -6963 10076 -6763 10092
rect -6705 10126 -6505 10164
rect -6705 10092 -6656 10126
rect -6622 10092 -6588 10126
rect -6554 10092 -6505 10126
rect -6705 10076 -6505 10092
rect -6447 10126 -6247 10164
rect -6447 10092 -6398 10126
rect -6364 10092 -6330 10126
rect -6296 10092 -6247 10126
rect -6447 10076 -6247 10092
rect -6189 10126 -5989 10164
rect -6189 10092 -6140 10126
rect -6106 10092 -6072 10126
rect -6038 10092 -5989 10126
rect -6189 10076 -5989 10092
rect -5931 10126 -5731 10164
rect -5931 10092 -5882 10126
rect -5848 10092 -5814 10126
rect -5780 10092 -5731 10126
rect -5931 10076 -5731 10092
rect -5673 10126 -5473 10164
rect -5673 10092 -5624 10126
rect -5590 10092 -5556 10126
rect -5522 10092 -5473 10126
rect -5673 10076 -5473 10092
rect -5415 10126 -5215 10164
rect -5415 10092 -5366 10126
rect -5332 10092 -5298 10126
rect -5264 10092 -5215 10126
rect -5415 10076 -5215 10092
rect -5157 10126 -4957 10164
rect -5157 10092 -5108 10126
rect -5074 10092 -5040 10126
rect -5006 10092 -4957 10126
rect -5157 10076 -4957 10092
rect -4899 10126 -4699 10164
rect -4899 10092 -4850 10126
rect -4816 10092 -4782 10126
rect -4748 10092 -4699 10126
rect -4899 10076 -4699 10092
rect -4641 10126 -4441 10164
rect -4641 10092 -4592 10126
rect -4558 10092 -4524 10126
rect -4490 10092 -4441 10126
rect -4641 10076 -4441 10092
rect -4383 10126 -4183 10164
rect -4383 10092 -4334 10126
rect -4300 10092 -4266 10126
rect -4232 10092 -4183 10126
rect -4383 10076 -4183 10092
rect -4125 10126 -3925 10164
rect -4125 10092 -4076 10126
rect -4042 10092 -4008 10126
rect -3974 10092 -3925 10126
rect -4125 10076 -3925 10092
rect -3867 10126 -3667 10164
rect -3867 10092 -3818 10126
rect -3784 10092 -3750 10126
rect -3716 10092 -3667 10126
rect -3867 10076 -3667 10092
rect 15000 11328 16000 11344
rect 15000 11294 15041 11328
rect 15075 11294 15109 11328
rect 15143 11294 15177 11328
rect 15211 11294 15245 11328
rect 15279 11294 15313 11328
rect 15347 11294 15381 11328
rect 15415 11294 15449 11328
rect 15483 11294 15517 11328
rect 15551 11294 15585 11328
rect 15619 11294 15653 11328
rect 15687 11294 15721 11328
rect 15755 11294 15789 11328
rect 15823 11294 15857 11328
rect 15891 11294 15925 11328
rect 15959 11294 16000 11328
rect 15000 11247 16000 11294
rect 16058 11328 17058 11344
rect 16058 11294 16099 11328
rect 16133 11294 16167 11328
rect 16201 11294 16235 11328
rect 16269 11294 16303 11328
rect 16337 11294 16371 11328
rect 16405 11294 16439 11328
rect 16473 11294 16507 11328
rect 16541 11294 16575 11328
rect 16609 11294 16643 11328
rect 16677 11294 16711 11328
rect 16745 11294 16779 11328
rect 16813 11294 16847 11328
rect 16881 11294 16915 11328
rect 16949 11294 16983 11328
rect 17017 11294 17058 11328
rect 16058 11247 17058 11294
rect -7734 9871 -7534 9887
rect -7734 9837 -7685 9871
rect -7651 9837 -7617 9871
rect -7583 9837 -7534 9871
rect -7734 9799 -7534 9837
rect -7268 9871 -7068 9887
rect -7268 9837 -7219 9871
rect -7185 9837 -7151 9871
rect -7117 9837 -7068 9871
rect -7268 9799 -7068 9837
rect -7010 9871 -6810 9887
rect -7010 9837 -6961 9871
rect -6927 9837 -6893 9871
rect -6859 9837 -6810 9871
rect -7010 9799 -6810 9837
rect -6752 9871 -6552 9887
rect -6752 9837 -6703 9871
rect -6669 9837 -6635 9871
rect -6601 9837 -6552 9871
rect -6752 9799 -6552 9837
rect -6494 9871 -6294 9887
rect -6494 9837 -6445 9871
rect -6411 9837 -6377 9871
rect -6343 9837 -6294 9871
rect -6494 9799 -6294 9837
rect -6236 9871 -6036 9887
rect -6236 9837 -6187 9871
rect -6153 9837 -6119 9871
rect -6085 9837 -6036 9871
rect -6236 9799 -6036 9837
rect -5978 9871 -5778 9887
rect -5978 9837 -5929 9871
rect -5895 9837 -5861 9871
rect -5827 9837 -5778 9871
rect -5978 9799 -5778 9837
rect -5720 9871 -5520 9887
rect -5720 9837 -5671 9871
rect -5637 9837 -5603 9871
rect -5569 9837 -5520 9871
rect -5720 9799 -5520 9837
rect -5462 9871 -5262 9887
rect -5462 9837 -5413 9871
rect -5379 9837 -5345 9871
rect -5311 9837 -5262 9871
rect -5462 9799 -5262 9837
rect -5204 9871 -5004 9887
rect -5204 9837 -5155 9871
rect -5121 9837 -5087 9871
rect -5053 9837 -5004 9871
rect -5204 9799 -5004 9837
rect -4946 9871 -4746 9887
rect -4946 9837 -4897 9871
rect -4863 9837 -4829 9871
rect -4795 9837 -4746 9871
rect -4946 9799 -4746 9837
rect -7734 8761 -7534 8799
rect -7734 8727 -7685 8761
rect -7651 8727 -7617 8761
rect -7583 8727 -7534 8761
rect -7734 8711 -7534 8727
rect -7268 8761 -7068 8799
rect -7268 8727 -7219 8761
rect -7185 8727 -7151 8761
rect -7117 8727 -7068 8761
rect -7268 8711 -7068 8727
rect -7010 8761 -6810 8799
rect -7010 8727 -6961 8761
rect -6927 8727 -6893 8761
rect -6859 8727 -6810 8761
rect -7010 8711 -6810 8727
rect -6752 8761 -6552 8799
rect -6752 8727 -6703 8761
rect -6669 8727 -6635 8761
rect -6601 8727 -6552 8761
rect -6752 8711 -6552 8727
rect -6494 8761 -6294 8799
rect -6494 8727 -6445 8761
rect -6411 8727 -6377 8761
rect -6343 8727 -6294 8761
rect -6494 8711 -6294 8727
rect -6236 8761 -6036 8799
rect -6236 8727 -6187 8761
rect -6153 8727 -6119 8761
rect -6085 8727 -6036 8761
rect -6236 8711 -6036 8727
rect -5978 8761 -5778 8799
rect -5978 8727 -5929 8761
rect -5895 8727 -5861 8761
rect -5827 8727 -5778 8761
rect -5978 8711 -5778 8727
rect -5720 8761 -5520 8799
rect -5720 8727 -5671 8761
rect -5637 8727 -5603 8761
rect -5569 8727 -5520 8761
rect -5720 8711 -5520 8727
rect -5462 8761 -5262 8799
rect -5462 8727 -5413 8761
rect -5379 8727 -5345 8761
rect -5311 8727 -5262 8761
rect -5462 8711 -5262 8727
rect -5204 8761 -5004 8799
rect -5204 8727 -5155 8761
rect -5121 8727 -5087 8761
rect -5053 8727 -5004 8761
rect -5204 8711 -5004 8727
rect -4946 8761 -4746 8799
rect -4946 8727 -4897 8761
rect -4863 8727 -4829 8761
rect -4795 8727 -4746 8761
rect -4946 8711 -4746 8727
rect -7734 7610 -7534 7626
rect -7734 7576 -7685 7610
rect -7651 7576 -7617 7610
rect -7583 7576 -7534 7610
rect -7734 7538 -7534 7576
rect -7476 7610 -7276 7626
rect -7476 7576 -7427 7610
rect -7393 7576 -7359 7610
rect -7325 7576 -7276 7610
rect -7476 7538 -7276 7576
rect -7218 7610 -7018 7626
rect -7218 7576 -7169 7610
rect -7135 7576 -7101 7610
rect -7067 7576 -7018 7610
rect -7218 7538 -7018 7576
rect -6960 7610 -6760 7626
rect -6960 7576 -6911 7610
rect -6877 7576 -6843 7610
rect -6809 7576 -6760 7610
rect -6960 7538 -6760 7576
rect -6702 7610 -6502 7626
rect -6702 7576 -6653 7610
rect -6619 7576 -6585 7610
rect -6551 7576 -6502 7610
rect -6702 7538 -6502 7576
rect -6444 7610 -6244 7626
rect -6444 7576 -6395 7610
rect -6361 7576 -6327 7610
rect -6293 7576 -6244 7610
rect -6444 7538 -6244 7576
rect -6186 7610 -5986 7626
rect -6186 7576 -6137 7610
rect -6103 7576 -6069 7610
rect -6035 7576 -5986 7610
rect -6186 7538 -5986 7576
rect -5928 7610 -5728 7626
rect -5928 7576 -5879 7610
rect -5845 7576 -5811 7610
rect -5777 7576 -5728 7610
rect -5928 7538 -5728 7576
rect -5670 7610 -5470 7626
rect -5670 7576 -5621 7610
rect -5587 7576 -5553 7610
rect -5519 7576 -5470 7610
rect -5670 7538 -5470 7576
rect -5412 7610 -5212 7626
rect -5412 7576 -5363 7610
rect -5329 7576 -5295 7610
rect -5261 7576 -5212 7610
rect -5412 7538 -5212 7576
rect -5154 7610 -4954 7626
rect -5154 7576 -5105 7610
rect -5071 7576 -5037 7610
rect -5003 7576 -4954 7610
rect -5154 7538 -4954 7576
rect -4896 7610 -4696 7626
rect -4896 7576 -4847 7610
rect -4813 7576 -4779 7610
rect -4745 7576 -4696 7610
rect -4896 7538 -4696 7576
rect -4638 7610 -4438 7626
rect -4638 7576 -4589 7610
rect -4555 7576 -4521 7610
rect -4487 7576 -4438 7610
rect -4638 7538 -4438 7576
rect -4380 7610 -4180 7626
rect -4380 7576 -4331 7610
rect -4297 7576 -4263 7610
rect -4229 7576 -4180 7610
rect -4380 7538 -4180 7576
rect -4122 7610 -3922 7626
rect -4122 7576 -4073 7610
rect -4039 7576 -4005 7610
rect -3971 7576 -3922 7610
rect -4122 7538 -3922 7576
rect -3864 7610 -3664 7626
rect -3864 7576 -3815 7610
rect -3781 7576 -3747 7610
rect -3713 7576 -3664 7610
rect -3864 7538 -3664 7576
rect 15000 8200 16000 8247
rect 15000 8166 15041 8200
rect 15075 8166 15109 8200
rect 15143 8166 15177 8200
rect 15211 8166 15245 8200
rect 15279 8166 15313 8200
rect 15347 8166 15381 8200
rect 15415 8166 15449 8200
rect 15483 8166 15517 8200
rect 15551 8166 15585 8200
rect 15619 8166 15653 8200
rect 15687 8166 15721 8200
rect 15755 8166 15789 8200
rect 15823 8166 15857 8200
rect 15891 8166 15925 8200
rect 15959 8166 16000 8200
rect 15000 8150 16000 8166
rect 16058 8200 17058 8247
rect 16058 8166 16099 8200
rect 16133 8166 16167 8200
rect 16201 8166 16235 8200
rect 16269 8166 16303 8200
rect 16337 8166 16371 8200
rect 16405 8166 16439 8200
rect 16473 8166 16507 8200
rect 16541 8166 16575 8200
rect 16609 8166 16643 8200
rect 16677 8166 16711 8200
rect 16745 8166 16779 8200
rect 16813 8166 16847 8200
rect 16881 8166 16915 8200
rect 16949 8166 16983 8200
rect 17017 8166 17058 8200
rect 16058 8150 17058 8166
rect 17524 11302 18524 11318
rect 17524 11268 17565 11302
rect 17599 11268 17633 11302
rect 17667 11268 17701 11302
rect 17735 11268 17769 11302
rect 17803 11268 17837 11302
rect 17871 11268 17905 11302
rect 17939 11268 17973 11302
rect 18007 11268 18041 11302
rect 18075 11268 18109 11302
rect 18143 11268 18177 11302
rect 18211 11268 18245 11302
rect 18279 11268 18313 11302
rect 18347 11268 18381 11302
rect 18415 11268 18449 11302
rect 18483 11268 18524 11302
rect 17524 11221 18524 11268
rect 18582 11302 19582 11318
rect 18582 11268 18623 11302
rect 18657 11268 18691 11302
rect 18725 11268 18759 11302
rect 18793 11268 18827 11302
rect 18861 11268 18895 11302
rect 18929 11268 18963 11302
rect 18997 11268 19031 11302
rect 19065 11268 19099 11302
rect 19133 11268 19167 11302
rect 19201 11268 19235 11302
rect 19269 11268 19303 11302
rect 19337 11268 19371 11302
rect 19405 11268 19439 11302
rect 19473 11268 19507 11302
rect 19541 11268 19582 11302
rect 18582 11221 19582 11268
rect 17524 8174 18524 8221
rect 17524 8140 17565 8174
rect 17599 8140 17633 8174
rect 17667 8140 17701 8174
rect 17735 8140 17769 8174
rect 17803 8140 17837 8174
rect 17871 8140 17905 8174
rect 17939 8140 17973 8174
rect 18007 8140 18041 8174
rect 18075 8140 18109 8174
rect 18143 8140 18177 8174
rect 18211 8140 18245 8174
rect 18279 8140 18313 8174
rect 18347 8140 18381 8174
rect 18415 8140 18449 8174
rect 18483 8140 18524 8174
rect 17524 8124 18524 8140
rect 18582 8174 19582 8221
rect 18582 8140 18623 8174
rect 18657 8140 18691 8174
rect 18725 8140 18759 8174
rect 18793 8140 18827 8174
rect 18861 8140 18895 8174
rect 18929 8140 18963 8174
rect 18997 8140 19031 8174
rect 19065 8140 19099 8174
rect 19133 8140 19167 8174
rect 19201 8140 19235 8174
rect 19269 8140 19303 8174
rect 19337 8140 19371 8174
rect 19405 8140 19439 8174
rect 19473 8140 19507 8174
rect 19541 8140 19582 8174
rect 18582 8124 19582 8140
rect 17480 7620 18480 7636
rect 17480 7586 17521 7620
rect 17555 7586 17589 7620
rect 17623 7586 17657 7620
rect 17691 7586 17725 7620
rect 17759 7586 17793 7620
rect 17827 7586 17861 7620
rect 17895 7586 17929 7620
rect 17963 7586 17997 7620
rect 18031 7586 18065 7620
rect 18099 7586 18133 7620
rect 18167 7586 18201 7620
rect 18235 7586 18269 7620
rect 18303 7586 18337 7620
rect 18371 7586 18405 7620
rect 18439 7586 18480 7620
rect 17480 7548 18480 7586
rect -7734 5500 -7534 5538
rect -7734 5466 -7685 5500
rect -7651 5466 -7617 5500
rect -7583 5466 -7534 5500
rect -7734 5450 -7534 5466
rect -7476 5500 -7276 5538
rect -7476 5466 -7427 5500
rect -7393 5466 -7359 5500
rect -7325 5466 -7276 5500
rect -7476 5450 -7276 5466
rect -7218 5500 -7018 5538
rect -7218 5466 -7169 5500
rect -7135 5466 -7101 5500
rect -7067 5466 -7018 5500
rect -7218 5450 -7018 5466
rect -6960 5500 -6760 5538
rect -6960 5466 -6911 5500
rect -6877 5466 -6843 5500
rect -6809 5466 -6760 5500
rect -6960 5450 -6760 5466
rect -6702 5500 -6502 5538
rect -6702 5466 -6653 5500
rect -6619 5466 -6585 5500
rect -6551 5466 -6502 5500
rect -6702 5450 -6502 5466
rect -6444 5500 -6244 5538
rect -6444 5466 -6395 5500
rect -6361 5466 -6327 5500
rect -6293 5466 -6244 5500
rect -6444 5450 -6244 5466
rect -6186 5500 -5986 5538
rect -6186 5466 -6137 5500
rect -6103 5466 -6069 5500
rect -6035 5466 -5986 5500
rect -6186 5450 -5986 5466
rect -5928 5500 -5728 5538
rect -5928 5466 -5879 5500
rect -5845 5466 -5811 5500
rect -5777 5466 -5728 5500
rect -5928 5450 -5728 5466
rect -5670 5500 -5470 5538
rect -5670 5466 -5621 5500
rect -5587 5466 -5553 5500
rect -5519 5466 -5470 5500
rect -5670 5450 -5470 5466
rect -5412 5500 -5212 5538
rect -5412 5466 -5363 5500
rect -5329 5466 -5295 5500
rect -5261 5466 -5212 5500
rect -5412 5450 -5212 5466
rect -5154 5500 -4954 5538
rect -5154 5466 -5105 5500
rect -5071 5466 -5037 5500
rect -5003 5466 -4954 5500
rect -5154 5450 -4954 5466
rect -4896 5500 -4696 5538
rect -4896 5466 -4847 5500
rect -4813 5466 -4779 5500
rect -4745 5466 -4696 5500
rect -4896 5450 -4696 5466
rect -4638 5500 -4438 5538
rect -4638 5466 -4589 5500
rect -4555 5466 -4521 5500
rect -4487 5466 -4438 5500
rect -4638 5450 -4438 5466
rect -4380 5500 -4180 5538
rect -4380 5466 -4331 5500
rect -4297 5466 -4263 5500
rect -4229 5466 -4180 5500
rect -4380 5450 -4180 5466
rect -4122 5500 -3922 5538
rect -4122 5466 -4073 5500
rect -4039 5466 -4005 5500
rect -3971 5466 -3922 5500
rect -4122 5450 -3922 5466
rect -3864 5500 -3664 5538
rect -3864 5466 -3815 5500
rect -3781 5466 -3747 5500
rect -3713 5466 -3664 5500
rect -3864 5450 -3664 5466
rect 17480 4510 18480 4548
rect 17480 4476 17521 4510
rect 17555 4476 17589 4510
rect 17623 4476 17657 4510
rect 17691 4476 17725 4510
rect 17759 4476 17793 4510
rect 17827 4476 17861 4510
rect 17895 4476 17929 4510
rect 17963 4476 17997 4510
rect 18031 4476 18065 4510
rect 18099 4476 18133 4510
rect 18167 4476 18201 4510
rect 18235 4476 18269 4510
rect 18303 4476 18337 4510
rect 18371 4476 18405 4510
rect 18439 4476 18480 4510
rect 17480 4460 18480 4476
rect 18930 7620 19930 7636
rect 18930 7586 18971 7620
rect 19005 7586 19039 7620
rect 19073 7586 19107 7620
rect 19141 7586 19175 7620
rect 19209 7586 19243 7620
rect 19277 7586 19311 7620
rect 19345 7586 19379 7620
rect 19413 7586 19447 7620
rect 19481 7586 19515 7620
rect 19549 7586 19583 7620
rect 19617 7586 19651 7620
rect 19685 7586 19719 7620
rect 19753 7586 19787 7620
rect 19821 7586 19855 7620
rect 19889 7586 19930 7620
rect 18930 7548 19930 7586
rect 38179 13559 38379 13585
rect 38437 13559 38637 13585
rect 38695 13559 38895 13585
rect 38953 13559 39153 13585
rect 39211 13559 39411 13585
rect 39469 13559 39669 13585
rect 39727 13559 39927 13585
rect 39985 13559 40185 13585
rect 40243 13559 40443 13585
rect 40501 13559 40701 13585
rect 23112 13269 23209 13310
rect 23112 13235 23128 13269
rect 23162 13235 23209 13269
rect 23112 13201 23209 13235
rect 23112 13167 23128 13201
rect 23162 13167 23209 13201
rect 23112 13133 23209 13167
rect 23112 13099 23128 13133
rect 23162 13099 23209 13133
rect 23112 13065 23209 13099
rect 23112 13031 23128 13065
rect 23162 13031 23209 13065
rect 23112 12997 23209 13031
rect 23112 12963 23128 12997
rect 23162 12963 23209 12997
rect 23112 12929 23209 12963
rect 23112 12895 23128 12929
rect 23162 12895 23209 12929
rect 23112 12861 23209 12895
rect 23112 12827 23128 12861
rect 23162 12827 23209 12861
rect 23112 12793 23209 12827
rect 23112 12759 23128 12793
rect 23162 12759 23209 12793
rect 23112 12725 23209 12759
rect 23112 12691 23128 12725
rect 23162 12691 23209 12725
rect 23112 12657 23209 12691
rect 23112 12623 23128 12657
rect 23162 12623 23209 12657
rect 23112 12589 23209 12623
rect 23112 12555 23128 12589
rect 23162 12555 23209 12589
rect 23112 12521 23209 12555
rect 23112 12487 23128 12521
rect 23162 12487 23209 12521
rect 23112 12453 23209 12487
rect 23112 12419 23128 12453
rect 23162 12419 23209 12453
rect 23112 12385 23209 12419
rect 23112 12351 23128 12385
rect 23162 12351 23209 12385
rect 23112 12310 23209 12351
rect 24209 13269 24306 13310
rect 24209 13235 24256 13269
rect 24290 13235 24306 13269
rect 24209 13201 24306 13235
rect 24209 13167 24256 13201
rect 24290 13167 24306 13201
rect 24209 13133 24306 13167
rect 24209 13099 24256 13133
rect 24290 13099 24306 13133
rect 24209 13065 24306 13099
rect 24209 13031 24256 13065
rect 24290 13031 24306 13065
rect 24209 12997 24306 13031
rect 24209 12963 24256 12997
rect 24290 12963 24306 12997
rect 24209 12929 24306 12963
rect 24209 12895 24256 12929
rect 24290 12895 24306 12929
rect 24209 12861 24306 12895
rect 24209 12827 24256 12861
rect 24290 12827 24306 12861
rect 24209 12793 24306 12827
rect 24209 12759 24256 12793
rect 24290 12759 24306 12793
rect 24209 12725 24306 12759
rect 24209 12691 24256 12725
rect 24290 12691 24306 12725
rect 24209 12657 24306 12691
rect 24209 12623 24256 12657
rect 24290 12623 24306 12657
rect 24209 12589 24306 12623
rect 24209 12555 24256 12589
rect 24290 12555 24306 12589
rect 24209 12521 24306 12555
rect 24209 12487 24256 12521
rect 24290 12487 24306 12521
rect 24209 12453 24306 12487
rect 24209 12419 24256 12453
rect 24290 12419 24306 12453
rect 24209 12385 24306 12419
rect 24209 12351 24256 12385
rect 24290 12351 24306 12385
rect 24209 12310 24306 12351
rect 24672 13263 24769 13304
rect 24672 13229 24688 13263
rect 24722 13229 24769 13263
rect 24672 13195 24769 13229
rect 24672 13161 24688 13195
rect 24722 13161 24769 13195
rect 24672 13127 24769 13161
rect 24672 13093 24688 13127
rect 24722 13093 24769 13127
rect 24672 13059 24769 13093
rect 24672 13025 24688 13059
rect 24722 13025 24769 13059
rect 24672 12991 24769 13025
rect 24672 12957 24688 12991
rect 24722 12957 24769 12991
rect 24672 12923 24769 12957
rect 24672 12889 24688 12923
rect 24722 12889 24769 12923
rect 24672 12855 24769 12889
rect 24672 12821 24688 12855
rect 24722 12821 24769 12855
rect 24672 12787 24769 12821
rect 24672 12753 24688 12787
rect 24722 12753 24769 12787
rect 24672 12719 24769 12753
rect 24672 12685 24688 12719
rect 24722 12685 24769 12719
rect 24672 12651 24769 12685
rect 24672 12617 24688 12651
rect 24722 12617 24769 12651
rect 24672 12583 24769 12617
rect 24672 12549 24688 12583
rect 24722 12549 24769 12583
rect 24672 12515 24769 12549
rect 24672 12481 24688 12515
rect 24722 12481 24769 12515
rect 24672 12447 24769 12481
rect 24672 12413 24688 12447
rect 24722 12413 24769 12447
rect 24672 12379 24769 12413
rect 24672 12345 24688 12379
rect 24722 12345 24769 12379
rect 24672 12304 24769 12345
rect 25769 13263 25866 13304
rect 25769 13229 25816 13263
rect 25850 13229 25866 13263
rect 25769 13195 25866 13229
rect 25769 13161 25816 13195
rect 25850 13161 25866 13195
rect 25769 13127 25866 13161
rect 25769 13093 25816 13127
rect 25850 13093 25866 13127
rect 25769 13059 25866 13093
rect 25769 13025 25816 13059
rect 25850 13025 25866 13059
rect 25769 12991 25866 13025
rect 25769 12957 25816 12991
rect 25850 12957 25866 12991
rect 25769 12923 25866 12957
rect 25769 12889 25816 12923
rect 25850 12889 25866 12923
rect 25769 12855 25866 12889
rect 25769 12821 25816 12855
rect 25850 12821 25866 12855
rect 25769 12787 25866 12821
rect 25769 12753 25816 12787
rect 25850 12753 25866 12787
rect 25769 12719 25866 12753
rect 25769 12685 25816 12719
rect 25850 12685 25866 12719
rect 25769 12651 25866 12685
rect 25769 12617 25816 12651
rect 25850 12617 25866 12651
rect 25769 12583 25866 12617
rect 25769 12549 25816 12583
rect 25850 12549 25866 12583
rect 25769 12515 25866 12549
rect 25769 12481 25816 12515
rect 25850 12481 25866 12515
rect 25769 12447 25866 12481
rect 25769 12413 25816 12447
rect 25850 12413 25866 12447
rect 25769 12379 25866 12413
rect 25769 12345 25816 12379
rect 25850 12345 25866 12379
rect 25769 12304 25866 12345
rect 23042 11729 23130 11770
rect 23042 11695 23058 11729
rect 23092 11695 23130 11729
rect 23042 11661 23130 11695
rect 23042 11627 23058 11661
rect 23092 11627 23130 11661
rect 23042 11593 23130 11627
rect 23042 11559 23058 11593
rect 23092 11559 23130 11593
rect 23042 11525 23130 11559
rect 23042 11491 23058 11525
rect 23092 11491 23130 11525
rect 23042 11457 23130 11491
rect 23042 11423 23058 11457
rect 23092 11423 23130 11457
rect 23042 11389 23130 11423
rect 23042 11355 23058 11389
rect 23092 11355 23130 11389
rect 23042 11321 23130 11355
rect 23042 11287 23058 11321
rect 23092 11287 23130 11321
rect 23042 11253 23130 11287
rect 23042 11219 23058 11253
rect 23092 11219 23130 11253
rect 23042 11185 23130 11219
rect 23042 11151 23058 11185
rect 23092 11151 23130 11185
rect 23042 11117 23130 11151
rect 23042 11083 23058 11117
rect 23092 11083 23130 11117
rect 23042 11049 23130 11083
rect 23042 11015 23058 11049
rect 23092 11015 23130 11049
rect 23042 10981 23130 11015
rect 23042 10947 23058 10981
rect 23092 10947 23130 10981
rect 23042 10913 23130 10947
rect 23042 10879 23058 10913
rect 23092 10879 23130 10913
rect 23042 10845 23130 10879
rect 23042 10811 23058 10845
rect 23092 10811 23130 10845
rect 23042 10770 23130 10811
rect 24130 11729 24218 11770
rect 24130 11695 24168 11729
rect 24202 11695 24218 11729
rect 24130 11661 24218 11695
rect 24130 11627 24168 11661
rect 24202 11627 24218 11661
rect 24130 11593 24218 11627
rect 24130 11559 24168 11593
rect 24202 11559 24218 11593
rect 24130 11525 24218 11559
rect 24130 11491 24168 11525
rect 24202 11491 24218 11525
rect 24130 11457 24218 11491
rect 24130 11423 24168 11457
rect 24202 11423 24218 11457
rect 24130 11389 24218 11423
rect 24130 11355 24168 11389
rect 24202 11355 24218 11389
rect 24130 11321 24218 11355
rect 24130 11287 24168 11321
rect 24202 11287 24218 11321
rect 24130 11253 24218 11287
rect 24130 11219 24168 11253
rect 24202 11219 24218 11253
rect 24130 11185 24218 11219
rect 24130 11151 24168 11185
rect 24202 11151 24218 11185
rect 24130 11117 24218 11151
rect 24130 11083 24168 11117
rect 24202 11083 24218 11117
rect 24130 11049 24218 11083
rect 24130 11015 24168 11049
rect 24202 11015 24218 11049
rect 24130 10981 24218 11015
rect 24130 10947 24168 10981
rect 24202 10947 24218 10981
rect 24130 10913 24218 10947
rect 24130 10879 24168 10913
rect 24202 10879 24218 10913
rect 24130 10845 24218 10879
rect 24130 10811 24168 10845
rect 24202 10811 24218 10845
rect 24130 10770 24218 10811
rect 24672 12205 24769 12246
rect 24672 12171 24688 12205
rect 24722 12171 24769 12205
rect 24672 12137 24769 12171
rect 24672 12103 24688 12137
rect 24722 12103 24769 12137
rect 24672 12069 24769 12103
rect 24672 12035 24688 12069
rect 24722 12035 24769 12069
rect 24672 12001 24769 12035
rect 24672 11967 24688 12001
rect 24722 11967 24769 12001
rect 24672 11933 24769 11967
rect 24672 11899 24688 11933
rect 24722 11899 24769 11933
rect 24672 11865 24769 11899
rect 24672 11831 24688 11865
rect 24722 11831 24769 11865
rect 24672 11797 24769 11831
rect 24672 11763 24688 11797
rect 24722 11763 24769 11797
rect 24672 11729 24769 11763
rect 24672 11695 24688 11729
rect 24722 11695 24769 11729
rect 24672 11661 24769 11695
rect 24672 11627 24688 11661
rect 24722 11627 24769 11661
rect 24672 11593 24769 11627
rect 24672 11559 24688 11593
rect 24722 11559 24769 11593
rect 24672 11525 24769 11559
rect 24672 11491 24688 11525
rect 24722 11491 24769 11525
rect 24672 11457 24769 11491
rect 24672 11423 24688 11457
rect 24722 11423 24769 11457
rect 24672 11389 24769 11423
rect 24672 11355 24688 11389
rect 24722 11355 24769 11389
rect 24672 11321 24769 11355
rect 24672 11287 24688 11321
rect 24722 11287 24769 11321
rect 24672 11246 24769 11287
rect 25769 12205 25866 12246
rect 25769 12171 25816 12205
rect 25850 12171 25866 12205
rect 25769 12137 25866 12171
rect 25769 12103 25816 12137
rect 25850 12103 25866 12137
rect 25769 12069 25866 12103
rect 25769 12035 25816 12069
rect 25850 12035 25866 12069
rect 25769 12001 25866 12035
rect 25769 11967 25816 12001
rect 25850 11967 25866 12001
rect 25769 11933 25866 11967
rect 25769 11899 25816 11933
rect 25850 11899 25866 11933
rect 25769 11865 25866 11899
rect 25769 11831 25816 11865
rect 25850 11831 25866 11865
rect 25769 11797 25866 11831
rect 25769 11763 25816 11797
rect 25850 11763 25866 11797
rect 25769 11729 25866 11763
rect 25769 11695 25816 11729
rect 25850 11695 25866 11729
rect 25769 11661 25866 11695
rect 25769 11627 25816 11661
rect 25850 11627 25866 11661
rect 25769 11593 25866 11627
rect 25769 11559 25816 11593
rect 25850 11559 25866 11593
rect 25769 11525 25866 11559
rect 25769 11491 25816 11525
rect 25850 11491 25866 11525
rect 25769 11457 25866 11491
rect 25769 11423 25816 11457
rect 25850 11423 25866 11457
rect 25769 11389 25866 11423
rect 25769 11355 25816 11389
rect 25850 11355 25866 11389
rect 25769 11321 25866 11355
rect 25769 11287 25816 11321
rect 25850 11287 25866 11321
rect 25769 11246 25866 11287
rect 24672 11147 24769 11188
rect 24672 11113 24688 11147
rect 24722 11113 24769 11147
rect 24672 11079 24769 11113
rect 24672 11045 24688 11079
rect 24722 11045 24769 11079
rect 24672 11011 24769 11045
rect 24672 10977 24688 11011
rect 24722 10977 24769 11011
rect 24672 10943 24769 10977
rect 24672 10909 24688 10943
rect 24722 10909 24769 10943
rect 24672 10875 24769 10909
rect 24672 10841 24688 10875
rect 24722 10841 24769 10875
rect 24672 10807 24769 10841
rect 24672 10773 24688 10807
rect 24722 10773 24769 10807
rect 24672 10739 24769 10773
rect 24672 10705 24688 10739
rect 24722 10705 24769 10739
rect 24672 10671 24769 10705
rect 24672 10637 24688 10671
rect 24722 10637 24769 10671
rect 24672 10603 24769 10637
rect 24672 10569 24688 10603
rect 24722 10569 24769 10603
rect 24672 10535 24769 10569
rect 24672 10501 24688 10535
rect 24722 10501 24769 10535
rect 24672 10467 24769 10501
rect 24672 10433 24688 10467
rect 24722 10433 24769 10467
rect 24672 10399 24769 10433
rect 24672 10365 24688 10399
rect 24722 10365 24769 10399
rect 24672 10331 24769 10365
rect 24672 10297 24688 10331
rect 24722 10297 24769 10331
rect 24672 10263 24769 10297
rect 24672 10229 24688 10263
rect 24722 10229 24769 10263
rect 24672 10188 24769 10229
rect 25769 11147 25866 11188
rect 25769 11113 25816 11147
rect 25850 11113 25866 11147
rect 25769 11079 25866 11113
rect 25769 11045 25816 11079
rect 25850 11045 25866 11079
rect 25769 11011 25866 11045
rect 25769 10977 25816 11011
rect 25850 10977 25866 11011
rect 25769 10943 25866 10977
rect 25769 10909 25816 10943
rect 25850 10909 25866 10943
rect 25769 10875 25866 10909
rect 25769 10841 25816 10875
rect 25850 10841 25866 10875
rect 25769 10807 25866 10841
rect 25769 10773 25816 10807
rect 25850 10773 25866 10807
rect 25769 10739 25866 10773
rect 25769 10705 25816 10739
rect 25850 10705 25866 10739
rect 25769 10671 25866 10705
rect 25769 10637 25816 10671
rect 25850 10637 25866 10671
rect 25769 10603 25866 10637
rect 25769 10569 25816 10603
rect 25850 10569 25866 10603
rect 25769 10535 25866 10569
rect 25769 10501 25816 10535
rect 25850 10501 25866 10535
rect 25769 10467 25866 10501
rect 25769 10433 25816 10467
rect 25850 10433 25866 10467
rect 25769 10399 25866 10433
rect 25769 10365 25816 10399
rect 25850 10365 25866 10399
rect 25769 10331 25866 10365
rect 25769 10297 25816 10331
rect 25850 10297 25866 10331
rect 25769 10263 25866 10297
rect 25769 10229 25816 10263
rect 25850 10229 25866 10263
rect 25769 10188 25866 10229
rect 24672 10089 24769 10130
rect 24672 10055 24688 10089
rect 24722 10055 24769 10089
rect 24672 10021 24769 10055
rect 24672 9987 24688 10021
rect 24722 9987 24769 10021
rect 24672 9953 24769 9987
rect 24672 9919 24688 9953
rect 24722 9919 24769 9953
rect 24672 9885 24769 9919
rect 24672 9851 24688 9885
rect 24722 9851 24769 9885
rect 24672 9817 24769 9851
rect 24672 9783 24688 9817
rect 24722 9783 24769 9817
rect 24672 9749 24769 9783
rect 24672 9715 24688 9749
rect 24722 9715 24769 9749
rect 24672 9681 24769 9715
rect 24672 9647 24688 9681
rect 24722 9647 24769 9681
rect 24672 9613 24769 9647
rect 24672 9579 24688 9613
rect 24722 9579 24769 9613
rect 24672 9545 24769 9579
rect 24672 9511 24688 9545
rect 24722 9511 24769 9545
rect 24672 9477 24769 9511
rect 24672 9443 24688 9477
rect 24722 9443 24769 9477
rect 24672 9409 24769 9443
rect 24672 9375 24688 9409
rect 24722 9375 24769 9409
rect 24672 9341 24769 9375
rect 24672 9307 24688 9341
rect 24722 9307 24769 9341
rect 24672 9273 24769 9307
rect 24672 9239 24688 9273
rect 24722 9239 24769 9273
rect 24672 9205 24769 9239
rect 24672 9171 24688 9205
rect 24722 9171 24769 9205
rect 24672 9130 24769 9171
rect 25769 10089 25866 10130
rect 25769 10055 25816 10089
rect 25850 10055 25866 10089
rect 25769 10021 25866 10055
rect 25769 9987 25816 10021
rect 25850 9987 25866 10021
rect 25769 9953 25866 9987
rect 25769 9919 25816 9953
rect 25850 9919 25866 9953
rect 25769 9885 25866 9919
rect 25769 9851 25816 9885
rect 25850 9851 25866 9885
rect 25769 9817 25866 9851
rect 25769 9783 25816 9817
rect 25850 9783 25866 9817
rect 25769 9749 25866 9783
rect 25769 9715 25816 9749
rect 25850 9715 25866 9749
rect 25769 9681 25866 9715
rect 25769 9647 25816 9681
rect 25850 9647 25866 9681
rect 25769 9613 25866 9647
rect 25769 9579 25816 9613
rect 25850 9579 25866 9613
rect 25769 9545 25866 9579
rect 25769 9511 25816 9545
rect 25850 9511 25866 9545
rect 25769 9477 25866 9511
rect 25769 9443 25816 9477
rect 25850 9443 25866 9477
rect 25769 9409 25866 9443
rect 25769 9375 25816 9409
rect 25850 9375 25866 9409
rect 25769 9341 25866 9375
rect 25769 9307 25816 9341
rect 25850 9307 25866 9341
rect 25769 9273 25866 9307
rect 25769 9239 25816 9273
rect 25850 9239 25866 9273
rect 25769 9205 25866 9239
rect 25769 9171 25816 9205
rect 25850 9171 25866 9205
rect 25769 9130 25866 9171
rect 23522 7793 23610 7834
rect 23522 7759 23538 7793
rect 23572 7759 23610 7793
rect 23522 7725 23610 7759
rect 23522 7691 23538 7725
rect 23572 7691 23610 7725
rect 23522 7657 23610 7691
rect 23522 7623 23538 7657
rect 23572 7623 23610 7657
rect 23522 7589 23610 7623
rect 23522 7555 23538 7589
rect 23572 7555 23610 7589
rect 23522 7521 23610 7555
rect 23522 7487 23538 7521
rect 23572 7487 23610 7521
rect 23522 7453 23610 7487
rect 23522 7419 23538 7453
rect 23572 7419 23610 7453
rect 23522 7385 23610 7419
rect 23522 7351 23538 7385
rect 23572 7351 23610 7385
rect 23522 7317 23610 7351
rect 23522 7283 23538 7317
rect 23572 7283 23610 7317
rect 23522 7249 23610 7283
rect 23522 7215 23538 7249
rect 23572 7215 23610 7249
rect 23522 7181 23610 7215
rect 23522 7147 23538 7181
rect 23572 7147 23610 7181
rect 23522 7113 23610 7147
rect 23522 7079 23538 7113
rect 23572 7079 23610 7113
rect 23522 7045 23610 7079
rect 23522 7011 23538 7045
rect 23572 7011 23610 7045
rect 23522 6977 23610 7011
rect 23522 6943 23538 6977
rect 23572 6943 23610 6977
rect 23522 6909 23610 6943
rect 23522 6875 23538 6909
rect 23572 6875 23610 6909
rect 23522 6834 23610 6875
rect 24610 7793 24698 7834
rect 24610 7759 24648 7793
rect 24682 7759 24698 7793
rect 24610 7725 24698 7759
rect 24610 7691 24648 7725
rect 24682 7691 24698 7725
rect 24610 7657 24698 7691
rect 24610 7623 24648 7657
rect 24682 7623 24698 7657
rect 24610 7589 24698 7623
rect 24610 7555 24648 7589
rect 24682 7555 24698 7589
rect 24610 7521 24698 7555
rect 24610 7487 24648 7521
rect 24682 7487 24698 7521
rect 24610 7453 24698 7487
rect 24610 7419 24648 7453
rect 24682 7419 24698 7453
rect 24610 7385 24698 7419
rect 24610 7351 24648 7385
rect 24682 7351 24698 7385
rect 24610 7317 24698 7351
rect 24610 7283 24648 7317
rect 24682 7283 24698 7317
rect 24610 7249 24698 7283
rect 24610 7215 24648 7249
rect 24682 7215 24698 7249
rect 24610 7181 24698 7215
rect 24610 7147 24648 7181
rect 24682 7147 24698 7181
rect 24610 7113 24698 7147
rect 24610 7079 24648 7113
rect 24682 7079 24698 7113
rect 24610 7045 24698 7079
rect 24610 7011 24648 7045
rect 24682 7011 24698 7045
rect 24610 6977 24698 7011
rect 24610 6943 24648 6977
rect 24682 6943 24698 6977
rect 24610 6909 24698 6943
rect 24610 6875 24648 6909
rect 24682 6875 24698 6909
rect 24610 6834 24698 6875
rect 23522 6735 23610 6776
rect 23522 6701 23538 6735
rect 23572 6701 23610 6735
rect 23522 6667 23610 6701
rect 23522 6633 23538 6667
rect 23572 6633 23610 6667
rect 23522 6599 23610 6633
rect 23522 6565 23538 6599
rect 23572 6565 23610 6599
rect 23522 6531 23610 6565
rect 23522 6497 23538 6531
rect 23572 6497 23610 6531
rect 23522 6463 23610 6497
rect 23522 6429 23538 6463
rect 23572 6429 23610 6463
rect 23522 6395 23610 6429
rect 23522 6361 23538 6395
rect 23572 6361 23610 6395
rect 23522 6327 23610 6361
rect 23522 6293 23538 6327
rect 23572 6293 23610 6327
rect 23522 6259 23610 6293
rect 23522 6225 23538 6259
rect 23572 6225 23610 6259
rect 23522 6191 23610 6225
rect 23522 6157 23538 6191
rect 23572 6157 23610 6191
rect 23522 6123 23610 6157
rect 23522 6089 23538 6123
rect 23572 6089 23610 6123
rect 23522 6055 23610 6089
rect 23522 6021 23538 6055
rect 23572 6021 23610 6055
rect 23522 5987 23610 6021
rect 23522 5953 23538 5987
rect 23572 5953 23610 5987
rect 23522 5919 23610 5953
rect 23522 5885 23538 5919
rect 23572 5885 23610 5919
rect 23522 5851 23610 5885
rect 23522 5817 23538 5851
rect 23572 5817 23610 5851
rect 23522 5776 23610 5817
rect 24610 6735 24698 6776
rect 24610 6701 24648 6735
rect 24682 6701 24698 6735
rect 24610 6667 24698 6701
rect 24610 6633 24648 6667
rect 24682 6633 24698 6667
rect 24610 6599 24698 6633
rect 24610 6565 24648 6599
rect 24682 6565 24698 6599
rect 24610 6531 24698 6565
rect 24610 6497 24648 6531
rect 24682 6497 24698 6531
rect 24610 6463 24698 6497
rect 24610 6429 24648 6463
rect 24682 6429 24698 6463
rect 24610 6395 24698 6429
rect 24610 6361 24648 6395
rect 24682 6361 24698 6395
rect 24610 6327 24698 6361
rect 24610 6293 24648 6327
rect 24682 6293 24698 6327
rect 24610 6259 24698 6293
rect 24610 6225 24648 6259
rect 24682 6225 24698 6259
rect 24610 6191 24698 6225
rect 24610 6157 24648 6191
rect 24682 6157 24698 6191
rect 24610 6123 24698 6157
rect 24610 6089 24648 6123
rect 24682 6089 24698 6123
rect 24610 6055 24698 6089
rect 24610 6021 24648 6055
rect 24682 6021 24698 6055
rect 24610 5987 24698 6021
rect 24610 5953 24648 5987
rect 24682 5953 24698 5987
rect 24610 5919 24698 5953
rect 24610 5885 24648 5919
rect 24682 5885 24698 5919
rect 24610 5851 24698 5885
rect 24610 5817 24648 5851
rect 24682 5817 24698 5851
rect 24610 5776 24698 5817
rect 23522 5677 23610 5718
rect 23522 5643 23538 5677
rect 23572 5643 23610 5677
rect 23522 5609 23610 5643
rect 23522 5575 23538 5609
rect 23572 5575 23610 5609
rect 23522 5541 23610 5575
rect 23522 5507 23538 5541
rect 23572 5507 23610 5541
rect 23522 5473 23610 5507
rect 23522 5439 23538 5473
rect 23572 5439 23610 5473
rect 23522 5405 23610 5439
rect 23522 5371 23538 5405
rect 23572 5371 23610 5405
rect 23522 5337 23610 5371
rect 23522 5303 23538 5337
rect 23572 5303 23610 5337
rect 23522 5269 23610 5303
rect 23522 5235 23538 5269
rect 23572 5235 23610 5269
rect 23522 5201 23610 5235
rect 23522 5167 23538 5201
rect 23572 5167 23610 5201
rect 23522 5133 23610 5167
rect 23522 5099 23538 5133
rect 23572 5099 23610 5133
rect 23522 5065 23610 5099
rect 23522 5031 23538 5065
rect 23572 5031 23610 5065
rect 23522 4997 23610 5031
rect 23522 4963 23538 4997
rect 23572 4963 23610 4997
rect 23522 4929 23610 4963
rect 23522 4895 23538 4929
rect 23572 4895 23610 4929
rect 23522 4861 23610 4895
rect 23522 4827 23538 4861
rect 23572 4827 23610 4861
rect 23522 4793 23610 4827
rect 23522 4759 23538 4793
rect 23572 4759 23610 4793
rect 23522 4718 23610 4759
rect 24610 5677 24698 5718
rect 24610 5643 24648 5677
rect 24682 5643 24698 5677
rect 24610 5609 24698 5643
rect 24610 5575 24648 5609
rect 24682 5575 24698 5609
rect 24610 5541 24698 5575
rect 24610 5507 24648 5541
rect 24682 5507 24698 5541
rect 24610 5473 24698 5507
rect 24610 5439 24648 5473
rect 24682 5439 24698 5473
rect 24610 5405 24698 5439
rect 24610 5371 24648 5405
rect 24682 5371 24698 5405
rect 24610 5337 24698 5371
rect 24610 5303 24648 5337
rect 24682 5303 24698 5337
rect 24610 5269 24698 5303
rect 24610 5235 24648 5269
rect 24682 5235 24698 5269
rect 24610 5201 24698 5235
rect 24610 5167 24648 5201
rect 24682 5167 24698 5201
rect 24610 5133 24698 5167
rect 24610 5099 24648 5133
rect 24682 5099 24698 5133
rect 24610 5065 24698 5099
rect 24610 5031 24648 5065
rect 24682 5031 24698 5065
rect 24610 4997 24698 5031
rect 24610 4963 24648 4997
rect 24682 4963 24698 4997
rect 24610 4929 24698 4963
rect 24610 4895 24648 4929
rect 24682 4895 24698 4929
rect 24610 4861 24698 4895
rect 24610 4827 24648 4861
rect 24682 4827 24698 4861
rect 24610 4793 24698 4827
rect 24610 4759 24648 4793
rect 24682 4759 24698 4793
rect 24610 4718 24698 4759
rect 18930 4510 19930 4548
rect 18930 4476 18971 4510
rect 19005 4476 19039 4510
rect 19073 4476 19107 4510
rect 19141 4476 19175 4510
rect 19209 4476 19243 4510
rect 19277 4476 19311 4510
rect 19345 4476 19379 4510
rect 19413 4476 19447 4510
rect 19481 4476 19515 4510
rect 19549 4476 19583 4510
rect 19617 4476 19651 4510
rect 19685 4476 19719 4510
rect 19753 4476 19787 4510
rect 19821 4476 19855 4510
rect 19889 4476 19930 4510
rect 18930 4460 19930 4476
rect 23522 4619 23610 4660
rect 23522 4585 23538 4619
rect 23572 4585 23610 4619
rect 23522 4551 23610 4585
rect 23522 4517 23538 4551
rect 23572 4517 23610 4551
rect 23522 4483 23610 4517
rect 23522 4449 23538 4483
rect 23572 4449 23610 4483
rect 23522 4415 23610 4449
rect 23522 4381 23538 4415
rect 23572 4381 23610 4415
rect 23522 4347 23610 4381
rect 23522 4313 23538 4347
rect 23572 4313 23610 4347
rect 23522 4279 23610 4313
rect 23522 4245 23538 4279
rect 23572 4245 23610 4279
rect 23522 4211 23610 4245
rect 23522 4177 23538 4211
rect 23572 4177 23610 4211
rect 23522 4143 23610 4177
rect 23522 4109 23538 4143
rect 23572 4109 23610 4143
rect 23522 4075 23610 4109
rect 23522 4041 23538 4075
rect 23572 4041 23610 4075
rect 23522 4007 23610 4041
rect 23522 3973 23538 4007
rect 23572 3973 23610 4007
rect 23522 3939 23610 3973
rect 23522 3905 23538 3939
rect 23572 3905 23610 3939
rect 23522 3871 23610 3905
rect 23522 3837 23538 3871
rect 23572 3837 23610 3871
rect 23522 3803 23610 3837
rect 23522 3769 23538 3803
rect 23572 3769 23610 3803
rect 23522 3735 23610 3769
rect 23522 3701 23538 3735
rect 23572 3701 23610 3735
rect 23522 3660 23610 3701
rect 24610 4619 24698 4660
rect 24610 4585 24648 4619
rect 24682 4585 24698 4619
rect 24610 4551 24698 4585
rect 24610 4517 24648 4551
rect 24682 4517 24698 4551
rect 24610 4483 24698 4517
rect 24610 4449 24648 4483
rect 24682 4449 24698 4483
rect 24610 4415 24698 4449
rect 24610 4381 24648 4415
rect 24682 4381 24698 4415
rect 24610 4347 24698 4381
rect 24610 4313 24648 4347
rect 24682 4313 24698 4347
rect 24610 4279 24698 4313
rect 24610 4245 24648 4279
rect 24682 4245 24698 4279
rect 24610 4211 24698 4245
rect 24610 4177 24648 4211
rect 24682 4177 24698 4211
rect 24610 4143 24698 4177
rect 24610 4109 24648 4143
rect 24682 4109 24698 4143
rect 24610 4075 24698 4109
rect 24610 4041 24648 4075
rect 24682 4041 24698 4075
rect 24610 4007 24698 4041
rect 24610 3973 24648 4007
rect 24682 3973 24698 4007
rect 24610 3939 24698 3973
rect 24610 3905 24648 3939
rect 24682 3905 24698 3939
rect 24610 3871 24698 3905
rect 24610 3837 24648 3871
rect 24682 3837 24698 3871
rect 24610 3803 24698 3837
rect 24610 3769 24648 3803
rect 24682 3769 24698 3803
rect 24610 3735 24698 3769
rect 24610 3701 24648 3735
rect 24682 3701 24698 3735
rect 24610 3660 24698 3701
rect 25022 7793 25110 7834
rect 25022 7759 25038 7793
rect 25072 7759 25110 7793
rect 25022 7725 25110 7759
rect 25022 7691 25038 7725
rect 25072 7691 25110 7725
rect 25022 7657 25110 7691
rect 25022 7623 25038 7657
rect 25072 7623 25110 7657
rect 25022 7589 25110 7623
rect 25022 7555 25038 7589
rect 25072 7555 25110 7589
rect 25022 7521 25110 7555
rect 25022 7487 25038 7521
rect 25072 7487 25110 7521
rect 25022 7453 25110 7487
rect 25022 7419 25038 7453
rect 25072 7419 25110 7453
rect 25022 7385 25110 7419
rect 25022 7351 25038 7385
rect 25072 7351 25110 7385
rect 25022 7317 25110 7351
rect 25022 7283 25038 7317
rect 25072 7283 25110 7317
rect 25022 7249 25110 7283
rect 25022 7215 25038 7249
rect 25072 7215 25110 7249
rect 25022 7181 25110 7215
rect 25022 7147 25038 7181
rect 25072 7147 25110 7181
rect 25022 7113 25110 7147
rect 25022 7079 25038 7113
rect 25072 7079 25110 7113
rect 25022 7045 25110 7079
rect 25022 7011 25038 7045
rect 25072 7011 25110 7045
rect 25022 6977 25110 7011
rect 25022 6943 25038 6977
rect 25072 6943 25110 6977
rect 25022 6909 25110 6943
rect 25022 6875 25038 6909
rect 25072 6875 25110 6909
rect 25022 6834 25110 6875
rect 26110 7793 26198 7834
rect 26110 7759 26148 7793
rect 26182 7759 26198 7793
rect 26110 7725 26198 7759
rect 26110 7691 26148 7725
rect 26182 7691 26198 7725
rect 26110 7657 26198 7691
rect 26110 7623 26148 7657
rect 26182 7623 26198 7657
rect 26110 7589 26198 7623
rect 26110 7555 26148 7589
rect 26182 7555 26198 7589
rect 26110 7521 26198 7555
rect 26110 7487 26148 7521
rect 26182 7487 26198 7521
rect 26110 7453 26198 7487
rect 26110 7419 26148 7453
rect 26182 7419 26198 7453
rect 26110 7385 26198 7419
rect 26110 7351 26148 7385
rect 26182 7351 26198 7385
rect 26110 7317 26198 7351
rect 26110 7283 26148 7317
rect 26182 7283 26198 7317
rect 26110 7249 26198 7283
rect 26110 7215 26148 7249
rect 26182 7215 26198 7249
rect 26110 7181 26198 7215
rect 26110 7147 26148 7181
rect 26182 7147 26198 7181
rect 26110 7113 26198 7147
rect 26110 7079 26148 7113
rect 26182 7079 26198 7113
rect 26110 7045 26198 7079
rect 26110 7011 26148 7045
rect 26182 7011 26198 7045
rect 26110 6977 26198 7011
rect 26110 6943 26148 6977
rect 26182 6943 26198 6977
rect 26110 6909 26198 6943
rect 26110 6875 26148 6909
rect 26182 6875 26198 6909
rect 26110 6834 26198 6875
rect 25022 6735 25110 6776
rect 25022 6701 25038 6735
rect 25072 6701 25110 6735
rect 25022 6667 25110 6701
rect 25022 6633 25038 6667
rect 25072 6633 25110 6667
rect 25022 6599 25110 6633
rect 25022 6565 25038 6599
rect 25072 6565 25110 6599
rect 25022 6531 25110 6565
rect 25022 6497 25038 6531
rect 25072 6497 25110 6531
rect 25022 6463 25110 6497
rect 25022 6429 25038 6463
rect 25072 6429 25110 6463
rect 25022 6395 25110 6429
rect 25022 6361 25038 6395
rect 25072 6361 25110 6395
rect 25022 6327 25110 6361
rect 25022 6293 25038 6327
rect 25072 6293 25110 6327
rect 25022 6259 25110 6293
rect 25022 6225 25038 6259
rect 25072 6225 25110 6259
rect 25022 6191 25110 6225
rect 25022 6157 25038 6191
rect 25072 6157 25110 6191
rect 25022 6123 25110 6157
rect 25022 6089 25038 6123
rect 25072 6089 25110 6123
rect 25022 6055 25110 6089
rect 25022 6021 25038 6055
rect 25072 6021 25110 6055
rect 25022 5987 25110 6021
rect 25022 5953 25038 5987
rect 25072 5953 25110 5987
rect 25022 5919 25110 5953
rect 25022 5885 25038 5919
rect 25072 5885 25110 5919
rect 25022 5851 25110 5885
rect 25022 5817 25038 5851
rect 25072 5817 25110 5851
rect 25022 5776 25110 5817
rect 26110 6735 26198 6776
rect 26110 6701 26148 6735
rect 26182 6701 26198 6735
rect 26110 6667 26198 6701
rect 26110 6633 26148 6667
rect 26182 6633 26198 6667
rect 26110 6599 26198 6633
rect 26110 6565 26148 6599
rect 26182 6565 26198 6599
rect 26110 6531 26198 6565
rect 26110 6497 26148 6531
rect 26182 6497 26198 6531
rect 26110 6463 26198 6497
rect 26110 6429 26148 6463
rect 26182 6429 26198 6463
rect 26110 6395 26198 6429
rect 26110 6361 26148 6395
rect 26182 6361 26198 6395
rect 26110 6327 26198 6361
rect 26110 6293 26148 6327
rect 26182 6293 26198 6327
rect 26110 6259 26198 6293
rect 26110 6225 26148 6259
rect 26182 6225 26198 6259
rect 26110 6191 26198 6225
rect 26110 6157 26148 6191
rect 26182 6157 26198 6191
rect 26110 6123 26198 6157
rect 26110 6089 26148 6123
rect 26182 6089 26198 6123
rect 26110 6055 26198 6089
rect 26110 6021 26148 6055
rect 26182 6021 26198 6055
rect 26110 5987 26198 6021
rect 26110 5953 26148 5987
rect 26182 5953 26198 5987
rect 26110 5919 26198 5953
rect 26110 5885 26148 5919
rect 26182 5885 26198 5919
rect 26110 5851 26198 5885
rect 26110 5817 26148 5851
rect 26182 5817 26198 5851
rect 26110 5776 26198 5817
rect 25022 5677 25110 5718
rect 25022 5643 25038 5677
rect 25072 5643 25110 5677
rect 25022 5609 25110 5643
rect 25022 5575 25038 5609
rect 25072 5575 25110 5609
rect 25022 5541 25110 5575
rect 25022 5507 25038 5541
rect 25072 5507 25110 5541
rect 25022 5473 25110 5507
rect 25022 5439 25038 5473
rect 25072 5439 25110 5473
rect 25022 5405 25110 5439
rect 25022 5371 25038 5405
rect 25072 5371 25110 5405
rect 25022 5337 25110 5371
rect 25022 5303 25038 5337
rect 25072 5303 25110 5337
rect 25022 5269 25110 5303
rect 25022 5235 25038 5269
rect 25072 5235 25110 5269
rect 25022 5201 25110 5235
rect 25022 5167 25038 5201
rect 25072 5167 25110 5201
rect 25022 5133 25110 5167
rect 25022 5099 25038 5133
rect 25072 5099 25110 5133
rect 25022 5065 25110 5099
rect 25022 5031 25038 5065
rect 25072 5031 25110 5065
rect 25022 4997 25110 5031
rect 25022 4963 25038 4997
rect 25072 4963 25110 4997
rect 25022 4929 25110 4963
rect 25022 4895 25038 4929
rect 25072 4895 25110 4929
rect 25022 4861 25110 4895
rect 25022 4827 25038 4861
rect 25072 4827 25110 4861
rect 25022 4793 25110 4827
rect 25022 4759 25038 4793
rect 25072 4759 25110 4793
rect 25022 4718 25110 4759
rect 26110 5677 26198 5718
rect 26110 5643 26148 5677
rect 26182 5643 26198 5677
rect 26110 5609 26198 5643
rect 26110 5575 26148 5609
rect 26182 5575 26198 5609
rect 26110 5541 26198 5575
rect 26110 5507 26148 5541
rect 26182 5507 26198 5541
rect 26110 5473 26198 5507
rect 26110 5439 26148 5473
rect 26182 5439 26198 5473
rect 26110 5405 26198 5439
rect 26110 5371 26148 5405
rect 26182 5371 26198 5405
rect 26110 5337 26198 5371
rect 26110 5303 26148 5337
rect 26182 5303 26198 5337
rect 26110 5269 26198 5303
rect 26110 5235 26148 5269
rect 26182 5235 26198 5269
rect 26110 5201 26198 5235
rect 26110 5167 26148 5201
rect 26182 5167 26198 5201
rect 26110 5133 26198 5167
rect 26110 5099 26148 5133
rect 26182 5099 26198 5133
rect 26110 5065 26198 5099
rect 26110 5031 26148 5065
rect 26182 5031 26198 5065
rect 26110 4997 26198 5031
rect 26110 4963 26148 4997
rect 26182 4963 26198 4997
rect 26110 4929 26198 4963
rect 26110 4895 26148 4929
rect 26182 4895 26198 4929
rect 26110 4861 26198 4895
rect 26110 4827 26148 4861
rect 26182 4827 26198 4861
rect 26110 4793 26198 4827
rect 26110 4759 26148 4793
rect 26182 4759 26198 4793
rect 26110 4718 26198 4759
rect 25022 4619 25110 4660
rect 25022 4585 25038 4619
rect 25072 4585 25110 4619
rect 25022 4551 25110 4585
rect 25022 4517 25038 4551
rect 25072 4517 25110 4551
rect 25022 4483 25110 4517
rect 25022 4449 25038 4483
rect 25072 4449 25110 4483
rect 25022 4415 25110 4449
rect 25022 4381 25038 4415
rect 25072 4381 25110 4415
rect 25022 4347 25110 4381
rect 25022 4313 25038 4347
rect 25072 4313 25110 4347
rect 25022 4279 25110 4313
rect 25022 4245 25038 4279
rect 25072 4245 25110 4279
rect 25022 4211 25110 4245
rect 25022 4177 25038 4211
rect 25072 4177 25110 4211
rect 25022 4143 25110 4177
rect 25022 4109 25038 4143
rect 25072 4109 25110 4143
rect 25022 4075 25110 4109
rect 25022 4041 25038 4075
rect 25072 4041 25110 4075
rect 25022 4007 25110 4041
rect 25022 3973 25038 4007
rect 25072 3973 25110 4007
rect 25022 3939 25110 3973
rect 25022 3905 25038 3939
rect 25072 3905 25110 3939
rect 25022 3871 25110 3905
rect 25022 3837 25038 3871
rect 25072 3837 25110 3871
rect 25022 3803 25110 3837
rect 25022 3769 25038 3803
rect 25072 3769 25110 3803
rect 25022 3735 25110 3769
rect 25022 3701 25038 3735
rect 25072 3701 25110 3735
rect 25022 3660 25110 3701
rect 26110 4619 26198 4660
rect 26110 4585 26148 4619
rect 26182 4585 26198 4619
rect 26110 4551 26198 4585
rect 26110 4517 26148 4551
rect 26182 4517 26198 4551
rect 26110 4483 26198 4517
rect 26110 4449 26148 4483
rect 26182 4449 26198 4483
rect 26110 4415 26198 4449
rect 26110 4381 26148 4415
rect 26182 4381 26198 4415
rect 26110 4347 26198 4381
rect 26110 4313 26148 4347
rect 26182 4313 26198 4347
rect 26110 4279 26198 4313
rect 26110 4245 26148 4279
rect 26182 4245 26198 4279
rect 26110 4211 26198 4245
rect 26110 4177 26148 4211
rect 26182 4177 26198 4211
rect 26110 4143 26198 4177
rect 26110 4109 26148 4143
rect 26182 4109 26198 4143
rect 26110 4075 26198 4109
rect 26110 4041 26148 4075
rect 26182 4041 26198 4075
rect 26110 4007 26198 4041
rect 26110 3973 26148 4007
rect 26182 3973 26198 4007
rect 26110 3939 26198 3973
rect 26110 3905 26148 3939
rect 26182 3905 26198 3939
rect 26110 3871 26198 3905
rect 26110 3837 26148 3871
rect 26182 3837 26198 3871
rect 26110 3803 26198 3837
rect 26110 3769 26148 3803
rect 26182 3769 26198 3803
rect 26110 3735 26198 3769
rect 26110 3701 26148 3735
rect 26182 3701 26198 3735
rect 26110 3660 26198 3701
rect 38200 13471 38346 13559
rect 38200 13437 38249 13471
rect 38283 13437 38346 13471
rect 38200 13424 38346 13437
rect 38975 13479 39135 13559
rect 38975 13445 39045 13479
rect 39079 13445 39135 13479
rect 38200 13390 38360 13424
rect 38975 13399 39135 13445
rect 39233 13474 39393 13559
rect 39233 13440 39282 13474
rect 39316 13440 39393 13474
rect 39233 13395 39393 13440
rect 40006 13476 40166 13559
rect 40006 13442 40076 13476
rect 40110 13442 40166 13476
rect 40006 13396 40166 13442
rect 40264 13476 40424 13559
rect 40264 13442 40331 13476
rect 40365 13442 40424 13476
rect 40264 13396 40424 13442
rect 36823 11986 37023 12002
rect 36823 11952 36872 11986
rect 36906 11952 36940 11986
rect 36974 11952 37023 11986
rect 36823 11914 37023 11952
rect 37081 11986 37281 12002
rect 37081 11952 37130 11986
rect 37164 11952 37198 11986
rect 37232 11952 37281 11986
rect 37081 11914 37281 11952
rect 37339 11986 37539 12002
rect 37339 11952 37388 11986
rect 37422 11952 37456 11986
rect 37490 11952 37539 11986
rect 37339 11914 37539 11952
rect 37597 11986 37797 12002
rect 37597 11952 37646 11986
rect 37680 11952 37714 11986
rect 37748 11952 37797 11986
rect 37597 11914 37797 11952
rect 37855 11986 38055 12002
rect 37855 11952 37904 11986
rect 37938 11952 37972 11986
rect 38006 11952 38055 11986
rect 37855 11914 38055 11952
rect 38113 11986 38313 12002
rect 38113 11952 38162 11986
rect 38196 11952 38230 11986
rect 38264 11952 38313 11986
rect 38113 11914 38313 11952
rect 38371 11986 38571 12002
rect 38371 11952 38420 11986
rect 38454 11952 38488 11986
rect 38522 11952 38571 11986
rect 38371 11914 38571 11952
rect 38629 11986 38829 12002
rect 38629 11952 38678 11986
rect 38712 11952 38746 11986
rect 38780 11952 38829 11986
rect 38629 11914 38829 11952
rect 38887 11986 39087 12002
rect 38887 11952 38936 11986
rect 38970 11952 39004 11986
rect 39038 11952 39087 11986
rect 38887 11914 39087 11952
rect 39145 11986 39345 12002
rect 39145 11952 39194 11986
rect 39228 11952 39262 11986
rect 39296 11952 39345 11986
rect 39145 11914 39345 11952
rect 39403 11986 39603 12002
rect 39403 11952 39452 11986
rect 39486 11952 39520 11986
rect 39554 11952 39603 11986
rect 39403 11914 39603 11952
rect 39661 11986 39861 12002
rect 39661 11952 39710 11986
rect 39744 11952 39778 11986
rect 39812 11952 39861 11986
rect 39661 11914 39861 11952
rect 39919 11986 40119 12002
rect 39919 11952 39968 11986
rect 40002 11952 40036 11986
rect 40070 11952 40119 11986
rect 39919 11914 40119 11952
rect 40177 11986 40377 12002
rect 40177 11952 40226 11986
rect 40260 11952 40294 11986
rect 40328 11952 40377 11986
rect 40177 11914 40377 11952
rect 40435 11986 40635 12002
rect 40435 11952 40484 11986
rect 40518 11952 40552 11986
rect 40586 11952 40635 11986
rect 40435 11914 40635 11952
rect 40693 11986 40893 12002
rect 40693 11952 40742 11986
rect 40776 11952 40810 11986
rect 40844 11952 40893 11986
rect 40693 11914 40893 11952
rect 40951 11986 41151 12002
rect 40951 11952 41000 11986
rect 41034 11952 41068 11986
rect 41102 11952 41151 11986
rect 40951 11914 41151 11952
rect 41209 11986 41409 12002
rect 41209 11952 41258 11986
rect 41292 11952 41326 11986
rect 41360 11952 41409 11986
rect 41209 11914 41409 11952
rect 41467 11986 41667 12002
rect 41467 11952 41516 11986
rect 41550 11952 41584 11986
rect 41618 11952 41667 11986
rect 41467 11914 41667 11952
rect 41725 11986 41925 12002
rect 41725 11952 41774 11986
rect 41808 11952 41842 11986
rect 41876 11952 41925 11986
rect 41725 11914 41925 11952
rect 36823 10876 37023 10914
rect 36823 10842 36872 10876
rect 36906 10842 36940 10876
rect 36974 10842 37023 10876
rect 36823 10826 37023 10842
rect 37081 10876 37281 10914
rect 37081 10842 37130 10876
rect 37164 10842 37198 10876
rect 37232 10842 37281 10876
rect 37081 10826 37281 10842
rect 37339 10876 37539 10914
rect 37339 10842 37388 10876
rect 37422 10842 37456 10876
rect 37490 10842 37539 10876
rect 37339 10826 37539 10842
rect 37597 10876 37797 10914
rect 37597 10842 37646 10876
rect 37680 10842 37714 10876
rect 37748 10842 37797 10876
rect 37597 10826 37797 10842
rect 37855 10876 38055 10914
rect 37855 10842 37904 10876
rect 37938 10842 37972 10876
rect 38006 10842 38055 10876
rect 37855 10826 38055 10842
rect 38113 10876 38313 10914
rect 38113 10842 38162 10876
rect 38196 10842 38230 10876
rect 38264 10842 38313 10876
rect 38113 10826 38313 10842
rect 38371 10876 38571 10914
rect 38371 10842 38420 10876
rect 38454 10842 38488 10876
rect 38522 10842 38571 10876
rect 38371 10826 38571 10842
rect 38629 10876 38829 10914
rect 38629 10842 38678 10876
rect 38712 10842 38746 10876
rect 38780 10842 38829 10876
rect 38629 10826 38829 10842
rect 38887 10876 39087 10914
rect 38887 10842 38936 10876
rect 38970 10842 39004 10876
rect 39038 10842 39087 10876
rect 38887 10826 39087 10842
rect 39145 10876 39345 10914
rect 39145 10842 39194 10876
rect 39228 10842 39262 10876
rect 39296 10842 39345 10876
rect 39145 10826 39345 10842
rect 39403 10876 39603 10914
rect 39403 10842 39452 10876
rect 39486 10842 39520 10876
rect 39554 10842 39603 10876
rect 39403 10826 39603 10842
rect 39661 10876 39861 10914
rect 39661 10842 39710 10876
rect 39744 10842 39778 10876
rect 39812 10842 39861 10876
rect 39661 10826 39861 10842
rect 39919 10876 40119 10914
rect 39919 10842 39968 10876
rect 40002 10842 40036 10876
rect 40070 10842 40119 10876
rect 39919 10826 40119 10842
rect 40177 10876 40377 10914
rect 40177 10842 40226 10876
rect 40260 10842 40294 10876
rect 40328 10842 40377 10876
rect 40177 10826 40377 10842
rect 40435 10876 40635 10914
rect 40435 10842 40484 10876
rect 40518 10842 40552 10876
rect 40586 10842 40635 10876
rect 40435 10826 40635 10842
rect 40693 10876 40893 10914
rect 40693 10842 40742 10876
rect 40776 10842 40810 10876
rect 40844 10842 40893 10876
rect 40693 10826 40893 10842
rect 40951 10876 41151 10914
rect 40951 10842 41000 10876
rect 41034 10842 41068 10876
rect 41102 10842 41151 10876
rect 40951 10826 41151 10842
rect 41209 10876 41409 10914
rect 41209 10842 41258 10876
rect 41292 10842 41326 10876
rect 41360 10842 41409 10876
rect 41209 10826 41409 10842
rect 41467 10876 41667 10914
rect 41467 10842 41516 10876
rect 41550 10842 41584 10876
rect 41618 10842 41667 10876
rect 41467 10826 41667 10842
rect 41725 10876 41925 10914
rect 41725 10842 41774 10876
rect 41808 10842 41842 10876
rect 41876 10842 41925 10876
rect 41725 10826 41925 10842
rect 37858 10621 38058 10637
rect 37858 10587 37907 10621
rect 37941 10587 37975 10621
rect 38009 10587 38058 10621
rect 37858 10549 38058 10587
rect 38324 10621 38524 10637
rect 38324 10587 38373 10621
rect 38407 10587 38441 10621
rect 38475 10587 38524 10621
rect 38324 10549 38524 10587
rect 38582 10621 38782 10637
rect 38582 10587 38631 10621
rect 38665 10587 38699 10621
rect 38733 10587 38782 10621
rect 38582 10549 38782 10587
rect 38840 10621 39040 10637
rect 38840 10587 38889 10621
rect 38923 10587 38957 10621
rect 38991 10587 39040 10621
rect 38840 10549 39040 10587
rect 39098 10621 39298 10637
rect 39098 10587 39147 10621
rect 39181 10587 39215 10621
rect 39249 10587 39298 10621
rect 39098 10549 39298 10587
rect 39356 10621 39556 10637
rect 39356 10587 39405 10621
rect 39439 10587 39473 10621
rect 39507 10587 39556 10621
rect 39356 10549 39556 10587
rect 39614 10621 39814 10637
rect 39614 10587 39663 10621
rect 39697 10587 39731 10621
rect 39765 10587 39814 10621
rect 39614 10549 39814 10587
rect 39872 10621 40072 10637
rect 39872 10587 39921 10621
rect 39955 10587 39989 10621
rect 40023 10587 40072 10621
rect 39872 10549 40072 10587
rect 40130 10621 40330 10637
rect 40130 10587 40179 10621
rect 40213 10587 40247 10621
rect 40281 10587 40330 10621
rect 40130 10549 40330 10587
rect 40388 10621 40588 10637
rect 40388 10587 40437 10621
rect 40471 10587 40505 10621
rect 40539 10587 40588 10621
rect 40388 10549 40588 10587
rect 40646 10621 40846 10637
rect 40646 10587 40695 10621
rect 40729 10587 40763 10621
rect 40797 10587 40846 10621
rect 40646 10549 40846 10587
rect 37858 9511 38058 9549
rect 37858 9477 37907 9511
rect 37941 9477 37975 9511
rect 38009 9477 38058 9511
rect 37858 9461 38058 9477
rect 38324 9511 38524 9549
rect 38324 9477 38373 9511
rect 38407 9477 38441 9511
rect 38475 9477 38524 9511
rect 38324 9461 38524 9477
rect 38582 9511 38782 9549
rect 38582 9477 38631 9511
rect 38665 9477 38699 9511
rect 38733 9477 38782 9511
rect 38582 9461 38782 9477
rect 38840 9511 39040 9549
rect 38840 9477 38889 9511
rect 38923 9477 38957 9511
rect 38991 9477 39040 9511
rect 38840 9461 39040 9477
rect 39098 9511 39298 9549
rect 39098 9477 39147 9511
rect 39181 9477 39215 9511
rect 39249 9477 39298 9511
rect 39098 9461 39298 9477
rect 39356 9511 39556 9549
rect 39356 9477 39405 9511
rect 39439 9477 39473 9511
rect 39507 9477 39556 9511
rect 39356 9461 39556 9477
rect 39614 9511 39814 9549
rect 39614 9477 39663 9511
rect 39697 9477 39731 9511
rect 39765 9477 39814 9511
rect 39614 9461 39814 9477
rect 39872 9511 40072 9549
rect 39872 9477 39921 9511
rect 39955 9477 39989 9511
rect 40023 9477 40072 9511
rect 39872 9461 40072 9477
rect 40130 9511 40330 9549
rect 40130 9477 40179 9511
rect 40213 9477 40247 9511
rect 40281 9477 40330 9511
rect 40130 9461 40330 9477
rect 40388 9511 40588 9549
rect 40388 9477 40437 9511
rect 40471 9477 40505 9511
rect 40539 9477 40588 9511
rect 40388 9461 40588 9477
rect 40646 9511 40846 9549
rect 40646 9477 40695 9511
rect 40729 9477 40763 9511
rect 40797 9477 40846 9511
rect 40646 9461 40846 9477
rect 37858 8360 38058 8376
rect 37858 8326 37907 8360
rect 37941 8326 37975 8360
rect 38009 8326 38058 8360
rect 37858 8288 38058 8326
rect 38116 8360 38316 8376
rect 38116 8326 38165 8360
rect 38199 8326 38233 8360
rect 38267 8326 38316 8360
rect 38116 8288 38316 8326
rect 38374 8360 38574 8376
rect 38374 8326 38423 8360
rect 38457 8326 38491 8360
rect 38525 8326 38574 8360
rect 38374 8288 38574 8326
rect 38632 8360 38832 8376
rect 38632 8326 38681 8360
rect 38715 8326 38749 8360
rect 38783 8326 38832 8360
rect 38632 8288 38832 8326
rect 38890 8360 39090 8376
rect 38890 8326 38939 8360
rect 38973 8326 39007 8360
rect 39041 8326 39090 8360
rect 38890 8288 39090 8326
rect 39148 8360 39348 8376
rect 39148 8326 39197 8360
rect 39231 8326 39265 8360
rect 39299 8326 39348 8360
rect 39148 8288 39348 8326
rect 39406 8360 39606 8376
rect 39406 8326 39455 8360
rect 39489 8326 39523 8360
rect 39557 8326 39606 8360
rect 39406 8288 39606 8326
rect 39664 8360 39864 8376
rect 39664 8326 39713 8360
rect 39747 8326 39781 8360
rect 39815 8326 39864 8360
rect 39664 8288 39864 8326
rect 39922 8360 40122 8376
rect 39922 8326 39971 8360
rect 40005 8326 40039 8360
rect 40073 8326 40122 8360
rect 39922 8288 40122 8326
rect 40180 8360 40380 8376
rect 40180 8326 40229 8360
rect 40263 8326 40297 8360
rect 40331 8326 40380 8360
rect 40180 8288 40380 8326
rect 40438 8360 40638 8376
rect 40438 8326 40487 8360
rect 40521 8326 40555 8360
rect 40589 8326 40638 8360
rect 40438 8288 40638 8326
rect 40696 8360 40896 8376
rect 40696 8326 40745 8360
rect 40779 8326 40813 8360
rect 40847 8326 40896 8360
rect 40696 8288 40896 8326
rect 40954 8360 41154 8376
rect 40954 8326 41003 8360
rect 41037 8326 41071 8360
rect 41105 8326 41154 8360
rect 40954 8288 41154 8326
rect 41212 8360 41412 8376
rect 41212 8326 41261 8360
rect 41295 8326 41329 8360
rect 41363 8326 41412 8360
rect 41212 8288 41412 8326
rect 41470 8360 41670 8376
rect 41470 8326 41519 8360
rect 41553 8326 41587 8360
rect 41621 8326 41670 8360
rect 41470 8288 41670 8326
rect 41728 8360 41928 8376
rect 41728 8326 41777 8360
rect 41811 8326 41845 8360
rect 41879 8326 41928 8360
rect 41728 8288 41928 8326
rect 37858 6250 38058 6288
rect 37858 6216 37907 6250
rect 37941 6216 37975 6250
rect 38009 6216 38058 6250
rect 37858 6200 38058 6216
rect 38116 6250 38316 6288
rect 38116 6216 38165 6250
rect 38199 6216 38233 6250
rect 38267 6216 38316 6250
rect 38116 6200 38316 6216
rect 38374 6250 38574 6288
rect 38374 6216 38423 6250
rect 38457 6216 38491 6250
rect 38525 6216 38574 6250
rect 38374 6200 38574 6216
rect 38632 6250 38832 6288
rect 38632 6216 38681 6250
rect 38715 6216 38749 6250
rect 38783 6216 38832 6250
rect 38632 6200 38832 6216
rect 38890 6250 39090 6288
rect 38890 6216 38939 6250
rect 38973 6216 39007 6250
rect 39041 6216 39090 6250
rect 38890 6200 39090 6216
rect 39148 6250 39348 6288
rect 39148 6216 39197 6250
rect 39231 6216 39265 6250
rect 39299 6216 39348 6250
rect 39148 6200 39348 6216
rect 39406 6250 39606 6288
rect 39406 6216 39455 6250
rect 39489 6216 39523 6250
rect 39557 6216 39606 6250
rect 39406 6200 39606 6216
rect 39664 6250 39864 6288
rect 39664 6216 39713 6250
rect 39747 6216 39781 6250
rect 39815 6216 39864 6250
rect 39664 6200 39864 6216
rect 39922 6250 40122 6288
rect 39922 6216 39971 6250
rect 40005 6216 40039 6250
rect 40073 6216 40122 6250
rect 39922 6200 40122 6216
rect 40180 6250 40380 6288
rect 40180 6216 40229 6250
rect 40263 6216 40297 6250
rect 40331 6216 40380 6250
rect 40180 6200 40380 6216
rect 40438 6250 40638 6288
rect 40438 6216 40487 6250
rect 40521 6216 40555 6250
rect 40589 6216 40638 6250
rect 40438 6200 40638 6216
rect 40696 6250 40896 6288
rect 40696 6216 40745 6250
rect 40779 6216 40813 6250
rect 40847 6216 40896 6250
rect 40696 6200 40896 6216
rect 40954 6250 41154 6288
rect 40954 6216 41003 6250
rect 41037 6216 41071 6250
rect 41105 6216 41154 6250
rect 40954 6200 41154 6216
rect 41212 6250 41412 6288
rect 41212 6216 41261 6250
rect 41295 6216 41329 6250
rect 41363 6216 41412 6250
rect 41212 6200 41412 6216
rect 41470 6250 41670 6288
rect 41470 6216 41519 6250
rect 41553 6216 41587 6250
rect 41621 6216 41670 6250
rect 41470 6200 41670 6216
rect 41728 6250 41928 6288
rect 41728 6216 41777 6250
rect 41811 6216 41845 6250
rect 41879 6216 41928 6250
rect 41728 6200 41928 6216
<< polycont >>
rect 23263 18794 23297 18828
rect 23331 18794 23365 18828
rect 23399 18794 23433 18828
rect 23467 18794 23501 18828
rect 23535 18794 23569 18828
rect 23603 18794 23637 18828
rect 23671 18794 23705 18828
rect 23739 18794 23773 18828
rect 23807 18794 23841 18828
rect 23875 18794 23909 18828
rect 23943 18794 23977 18828
rect 24011 18794 24045 18828
rect 24079 18794 24113 18828
rect 24147 18794 24181 18828
rect -2885 18140 -2851 18174
rect -2817 18140 -2783 18174
rect -2627 18140 -2593 18174
rect -2559 18140 -2525 18174
rect -2369 18140 -2335 18174
rect -2301 18140 -2267 18174
rect -2111 18140 -2077 18174
rect -2043 18140 -2009 18174
rect -1853 18140 -1819 18174
rect -1785 18140 -1751 18174
rect -1595 18140 -1561 18174
rect -1527 18140 -1493 18174
rect -1337 18140 -1303 18174
rect -1269 18140 -1235 18174
rect -1079 18140 -1045 18174
rect -1011 18140 -977 18174
rect -821 18140 -787 18174
rect -753 18140 -719 18174
rect -563 18140 -529 18174
rect -495 18140 -461 18174
rect -6353 17271 -6319 17305
rect -6285 17271 -6251 17305
rect -6095 17271 -6061 17305
rect -6027 17271 -5993 17305
rect -6353 16143 -6319 16177
rect -6285 16143 -6251 16177
rect -6095 16143 -6061 16177
rect -6027 16143 -5993 16177
rect 23263 17666 23297 17700
rect 23331 17666 23365 17700
rect 23399 17666 23433 17700
rect 23467 17666 23501 17700
rect 23535 17666 23569 17700
rect 23603 17666 23637 17700
rect 23671 17666 23705 17700
rect 23739 17666 23773 17700
rect 23807 17666 23841 17700
rect 23875 17666 23909 17700
rect 23943 17666 23977 17700
rect 24011 17666 24045 17700
rect 24079 17666 24113 17700
rect 24147 17666 24181 17700
rect 24779 18794 24813 18828
rect 24847 18794 24881 18828
rect 24915 18794 24949 18828
rect 24983 18794 25017 18828
rect 25051 18794 25085 18828
rect 25119 18794 25153 18828
rect 25187 18794 25221 18828
rect 25255 18794 25289 18828
rect 25323 18794 25357 18828
rect 25391 18794 25425 18828
rect 25459 18794 25493 18828
rect 25527 18794 25561 18828
rect 25595 18794 25629 18828
rect 25663 18794 25697 18828
rect 25837 18794 25871 18828
rect 25905 18794 25939 18828
rect 25973 18794 26007 18828
rect 26041 18794 26075 18828
rect 26109 18794 26143 18828
rect 26177 18794 26211 18828
rect 26245 18794 26279 18828
rect 26313 18794 26347 18828
rect 26381 18794 26415 18828
rect 26449 18794 26483 18828
rect 26517 18794 26551 18828
rect 26585 18794 26619 18828
rect 26653 18794 26687 18828
rect 26721 18794 26755 18828
rect 26895 18794 26929 18828
rect 26963 18794 26997 18828
rect 27031 18794 27065 18828
rect 27099 18794 27133 18828
rect 27167 18794 27201 18828
rect 27235 18794 27269 18828
rect 27303 18794 27337 18828
rect 27371 18794 27405 18828
rect 27439 18794 27473 18828
rect 27507 18794 27541 18828
rect 27575 18794 27609 18828
rect 27643 18794 27677 18828
rect 27711 18794 27745 18828
rect 27779 18794 27813 18828
rect -2885 16012 -2851 16046
rect -2817 16012 -2783 16046
rect -2627 16012 -2593 16046
rect -2559 16012 -2525 16046
rect -2369 16012 -2335 16046
rect -2301 16012 -2267 16046
rect -2111 16012 -2077 16046
rect -2043 16012 -2009 16046
rect -1853 16012 -1819 16046
rect -1785 16012 -1751 16046
rect -1595 16012 -1561 16046
rect -1527 16012 -1493 16046
rect -1337 16012 -1303 16046
rect -1269 16012 -1235 16046
rect -1079 16012 -1045 16046
rect -1011 16012 -977 16046
rect -821 16012 -787 16046
rect -753 16012 -719 16046
rect -563 16012 -529 16046
rect -495 16012 -461 16046
rect 23237 17174 23271 17208
rect 23305 17174 23339 17208
rect 23373 17174 23407 17208
rect 23441 17174 23475 17208
rect 23509 17174 23543 17208
rect 23577 17174 23611 17208
rect 23645 17174 23679 17208
rect 23713 17174 23747 17208
rect 23781 17174 23815 17208
rect 23849 17174 23883 17208
rect 23917 17174 23951 17208
rect 23985 17174 24019 17208
rect 24053 17174 24087 17208
rect 24121 17174 24155 17208
rect 42707 18890 42741 18924
rect 42775 18890 42809 18924
rect 42965 18890 42999 18924
rect 43033 18890 43067 18924
rect 43223 18890 43257 18924
rect 43291 18890 43325 18924
rect 43481 18890 43515 18924
rect 43549 18890 43583 18924
rect 43739 18890 43773 18924
rect 43807 18890 43841 18924
rect 43997 18890 44031 18924
rect 44065 18890 44099 18924
rect 44255 18890 44289 18924
rect 44323 18890 44357 18924
rect 44513 18890 44547 18924
rect 44581 18890 44615 18924
rect 44771 18890 44805 18924
rect 44839 18890 44873 18924
rect 45029 18890 45063 18924
rect 45097 18890 45131 18924
rect 24779 17066 24813 17100
rect 24847 17066 24881 17100
rect 24915 17066 24949 17100
rect 24983 17066 25017 17100
rect 25051 17066 25085 17100
rect 25119 17066 25153 17100
rect 25187 17066 25221 17100
rect 25255 17066 25289 17100
rect 25323 17066 25357 17100
rect 25391 17066 25425 17100
rect 25459 17066 25493 17100
rect 25527 17066 25561 17100
rect 25595 17066 25629 17100
rect 25663 17066 25697 17100
rect 25837 17066 25871 17100
rect 25905 17066 25939 17100
rect 25973 17066 26007 17100
rect 26041 17066 26075 17100
rect 26109 17066 26143 17100
rect 26177 17066 26211 17100
rect 26245 17066 26279 17100
rect 26313 17066 26347 17100
rect 26381 17066 26415 17100
rect 26449 17066 26483 17100
rect 26517 17066 26551 17100
rect 26585 17066 26619 17100
rect 26653 17066 26687 17100
rect 26721 17066 26755 17100
rect 26895 17066 26929 17100
rect 26963 17066 26997 17100
rect 27031 17066 27065 17100
rect 27099 17066 27133 17100
rect 27167 17066 27201 17100
rect 27235 17066 27269 17100
rect 27303 17066 27337 17100
rect 27371 17066 27405 17100
rect 27439 17066 27473 17100
rect 27507 17066 27541 17100
rect 27575 17066 27609 17100
rect 27643 17066 27677 17100
rect 27711 17066 27745 17100
rect 27779 17066 27813 17100
rect 39239 18021 39273 18055
rect 39307 18021 39341 18055
rect 39497 18021 39531 18055
rect 39565 18021 39599 18055
rect 39239 16893 39273 16927
rect 39307 16893 39341 16927
rect 39497 16893 39531 16927
rect 39565 16893 39599 16927
rect 23237 16064 23271 16098
rect 23305 16064 23339 16098
rect 23373 16064 23407 16098
rect 23441 16064 23475 16098
rect 23509 16064 23543 16098
rect 23577 16064 23611 16098
rect 23645 16064 23679 16098
rect 23713 16064 23747 16098
rect 23781 16064 23815 16098
rect 23849 16064 23883 16098
rect 23917 16064 23951 16098
rect 23985 16064 24019 16098
rect 24053 16064 24087 16098
rect 24121 16064 24155 16098
rect 42707 16762 42741 16796
rect 42775 16762 42809 16796
rect 42965 16762 42999 16796
rect 43033 16762 43067 16796
rect 43223 16762 43257 16796
rect 43291 16762 43325 16796
rect 43481 16762 43515 16796
rect 43549 16762 43583 16796
rect 43739 16762 43773 16796
rect 43807 16762 43841 16796
rect 43997 16762 44031 16796
rect 44065 16762 44099 16796
rect 44255 16762 44289 16796
rect 44323 16762 44357 16796
rect 44513 16762 44547 16796
rect 44581 16762 44615 16796
rect 44771 16762 44805 16796
rect 44839 16762 44873 16796
rect 45029 16762 45063 16796
rect 45097 16762 45131 16796
rect -7080 14934 -7046 14968
rect -6820 14934 -6786 14968
rect -6028 14923 -5994 14957
rect -5778 14910 -5744 14944
rect -5007 14914 -4973 14948
rect -7343 12687 -7309 12721
rect -6547 12695 -6513 12729
rect -6310 12690 -6276 12724
rect -5516 12692 -5482 12726
rect -5261 12692 -5227 12726
rect 13081 14814 13115 14848
rect 13149 14814 13183 14848
rect 13217 14814 13251 14848
rect 13285 14814 13319 14848
rect 13353 14814 13387 14848
rect 13421 14814 13455 14848
rect 13489 14814 13523 14848
rect 13557 14814 13591 14848
rect 13625 14814 13659 14848
rect 13693 14814 13727 14848
rect 13761 14814 13795 14848
rect 13829 14814 13863 14848
rect 13897 14814 13931 14848
rect 13965 14814 13999 14848
rect 14139 14814 14173 14848
rect 14207 14814 14241 14848
rect 14275 14814 14309 14848
rect 14343 14814 14377 14848
rect 14411 14814 14445 14848
rect 14479 14814 14513 14848
rect 14547 14814 14581 14848
rect 14615 14814 14649 14848
rect 14683 14814 14717 14848
rect 14751 14814 14785 14848
rect 14819 14814 14853 14848
rect 14887 14814 14921 14848
rect 14955 14814 14989 14848
rect 15023 14814 15057 14848
rect 13081 11686 13115 11720
rect 13149 11686 13183 11720
rect 13217 11686 13251 11720
rect 13285 11686 13319 11720
rect 13353 11686 13387 11720
rect 13421 11686 13455 11720
rect 13489 11686 13523 11720
rect 13557 11686 13591 11720
rect 13625 11686 13659 11720
rect 13693 11686 13727 11720
rect 13761 11686 13795 11720
rect 13829 11686 13863 11720
rect 13897 11686 13931 11720
rect 13965 11686 13999 11720
rect 14139 11686 14173 11720
rect 14207 11686 14241 11720
rect 14275 11686 14309 11720
rect 14343 11686 14377 11720
rect 14411 11686 14445 11720
rect 14479 11686 14513 11720
rect 14547 11686 14581 11720
rect 14615 11686 14649 11720
rect 14683 11686 14717 11720
rect 14751 11686 14785 11720
rect 14819 11686 14853 11720
rect 14887 11686 14921 11720
rect 14955 11686 14989 11720
rect 15023 11686 15057 11720
rect 15651 14814 15685 14848
rect 15719 14814 15753 14848
rect 15787 14814 15821 14848
rect 15855 14814 15889 14848
rect 15923 14814 15957 14848
rect 15991 14814 16025 14848
rect 16059 14814 16093 14848
rect 16127 14814 16161 14848
rect 16195 14814 16229 14848
rect 16263 14814 16297 14848
rect 16331 14814 16365 14848
rect 16399 14814 16433 14848
rect 16467 14814 16501 14848
rect 16535 14814 16569 14848
rect 15651 11686 15685 11720
rect 15719 11686 15753 11720
rect 15787 11686 15821 11720
rect 15855 11686 15889 11720
rect 15923 11686 15957 11720
rect 15991 11686 16025 11720
rect 16059 11686 16093 11720
rect 16127 11686 16161 11720
rect 16195 11686 16229 11720
rect 16263 11686 16297 11720
rect 16331 11686 16365 11720
rect 16399 11686 16433 11720
rect 16467 11686 16501 11720
rect 16535 11686 16569 11720
rect 17161 14824 17195 14858
rect 17229 14824 17263 14858
rect 17297 14824 17331 14858
rect 17365 14824 17399 14858
rect 17433 14824 17467 14858
rect 17501 14824 17535 14858
rect 17569 14824 17603 14858
rect 17637 14824 17671 14858
rect 17705 14824 17739 14858
rect 17773 14824 17807 14858
rect 17841 14824 17875 14858
rect 17909 14824 17943 14858
rect 17977 14824 18011 14858
rect 18045 14824 18079 14858
rect 17161 11696 17195 11730
rect 17229 11696 17263 11730
rect 17297 11696 17331 11730
rect 17365 11696 17399 11730
rect 17433 11696 17467 11730
rect 17501 11696 17535 11730
rect 17569 11696 17603 11730
rect 17637 11696 17671 11730
rect 17705 11696 17739 11730
rect 17773 11696 17807 11730
rect 17841 11696 17875 11730
rect 17909 11696 17943 11730
rect 17977 11696 18011 11730
rect 18045 11696 18079 11730
rect 18625 14808 18659 14842
rect 18693 14808 18727 14842
rect 18761 14808 18795 14842
rect 18829 14808 18863 14842
rect 18897 14808 18931 14842
rect 18965 14808 18999 14842
rect 19033 14808 19067 14842
rect 19101 14808 19135 14842
rect 19169 14808 19203 14842
rect 19237 14808 19271 14842
rect 19305 14808 19339 14842
rect 19373 14808 19407 14842
rect 19441 14808 19475 14842
rect 19509 14808 19543 14842
rect 38512 15684 38546 15718
rect 38772 15684 38806 15718
rect 39564 15673 39598 15707
rect 39814 15660 39848 15694
rect 40585 15664 40619 15698
rect 18625 11680 18659 11714
rect 18693 11680 18727 11714
rect 18761 11680 18795 11714
rect 18829 11680 18863 11714
rect 18897 11680 18931 11714
rect 18965 11680 18999 11714
rect 19033 11680 19067 11714
rect 19101 11680 19135 11714
rect 19169 11680 19203 11714
rect 19237 11680 19271 11714
rect 19305 11680 19339 11714
rect 19373 11680 19407 11714
rect 19441 11680 19475 11714
rect 19509 11680 19543 11714
rect -8720 11202 -8686 11236
rect -8652 11202 -8618 11236
rect -8462 11202 -8428 11236
rect -8394 11202 -8360 11236
rect -8204 11202 -8170 11236
rect -8136 11202 -8102 11236
rect -7946 11202 -7912 11236
rect -7878 11202 -7844 11236
rect -7688 11202 -7654 11236
rect -7620 11202 -7586 11236
rect -7430 11202 -7396 11236
rect -7362 11202 -7328 11236
rect -7172 11202 -7138 11236
rect -7104 11202 -7070 11236
rect -6914 11202 -6880 11236
rect -6846 11202 -6812 11236
rect -6656 11202 -6622 11236
rect -6588 11202 -6554 11236
rect -6398 11202 -6364 11236
rect -6330 11202 -6296 11236
rect -6140 11202 -6106 11236
rect -6072 11202 -6038 11236
rect -5882 11202 -5848 11236
rect -5814 11202 -5780 11236
rect -5624 11202 -5590 11236
rect -5556 11202 -5522 11236
rect -5366 11202 -5332 11236
rect -5298 11202 -5264 11236
rect -5108 11202 -5074 11236
rect -5040 11202 -5006 11236
rect -4850 11202 -4816 11236
rect -4782 11202 -4748 11236
rect -4592 11202 -4558 11236
rect -4524 11202 -4490 11236
rect -4334 11202 -4300 11236
rect -4266 11202 -4232 11236
rect -4076 11202 -4042 11236
rect -4008 11202 -3974 11236
rect -3818 11202 -3784 11236
rect -3750 11202 -3716 11236
rect -8720 10092 -8686 10126
rect -8652 10092 -8618 10126
rect -8462 10092 -8428 10126
rect -8394 10092 -8360 10126
rect -8204 10092 -8170 10126
rect -8136 10092 -8102 10126
rect -7946 10092 -7912 10126
rect -7878 10092 -7844 10126
rect -7688 10092 -7654 10126
rect -7620 10092 -7586 10126
rect -7430 10092 -7396 10126
rect -7362 10092 -7328 10126
rect -7172 10092 -7138 10126
rect -7104 10092 -7070 10126
rect -6914 10092 -6880 10126
rect -6846 10092 -6812 10126
rect -6656 10092 -6622 10126
rect -6588 10092 -6554 10126
rect -6398 10092 -6364 10126
rect -6330 10092 -6296 10126
rect -6140 10092 -6106 10126
rect -6072 10092 -6038 10126
rect -5882 10092 -5848 10126
rect -5814 10092 -5780 10126
rect -5624 10092 -5590 10126
rect -5556 10092 -5522 10126
rect -5366 10092 -5332 10126
rect -5298 10092 -5264 10126
rect -5108 10092 -5074 10126
rect -5040 10092 -5006 10126
rect -4850 10092 -4816 10126
rect -4782 10092 -4748 10126
rect -4592 10092 -4558 10126
rect -4524 10092 -4490 10126
rect -4334 10092 -4300 10126
rect -4266 10092 -4232 10126
rect -4076 10092 -4042 10126
rect -4008 10092 -3974 10126
rect -3818 10092 -3784 10126
rect -3750 10092 -3716 10126
rect 15041 11294 15075 11328
rect 15109 11294 15143 11328
rect 15177 11294 15211 11328
rect 15245 11294 15279 11328
rect 15313 11294 15347 11328
rect 15381 11294 15415 11328
rect 15449 11294 15483 11328
rect 15517 11294 15551 11328
rect 15585 11294 15619 11328
rect 15653 11294 15687 11328
rect 15721 11294 15755 11328
rect 15789 11294 15823 11328
rect 15857 11294 15891 11328
rect 15925 11294 15959 11328
rect 16099 11294 16133 11328
rect 16167 11294 16201 11328
rect 16235 11294 16269 11328
rect 16303 11294 16337 11328
rect 16371 11294 16405 11328
rect 16439 11294 16473 11328
rect 16507 11294 16541 11328
rect 16575 11294 16609 11328
rect 16643 11294 16677 11328
rect 16711 11294 16745 11328
rect 16779 11294 16813 11328
rect 16847 11294 16881 11328
rect 16915 11294 16949 11328
rect 16983 11294 17017 11328
rect -7685 9837 -7651 9871
rect -7617 9837 -7583 9871
rect -7219 9837 -7185 9871
rect -7151 9837 -7117 9871
rect -6961 9837 -6927 9871
rect -6893 9837 -6859 9871
rect -6703 9837 -6669 9871
rect -6635 9837 -6601 9871
rect -6445 9837 -6411 9871
rect -6377 9837 -6343 9871
rect -6187 9837 -6153 9871
rect -6119 9837 -6085 9871
rect -5929 9837 -5895 9871
rect -5861 9837 -5827 9871
rect -5671 9837 -5637 9871
rect -5603 9837 -5569 9871
rect -5413 9837 -5379 9871
rect -5345 9837 -5311 9871
rect -5155 9837 -5121 9871
rect -5087 9837 -5053 9871
rect -4897 9837 -4863 9871
rect -4829 9837 -4795 9871
rect -7685 8727 -7651 8761
rect -7617 8727 -7583 8761
rect -7219 8727 -7185 8761
rect -7151 8727 -7117 8761
rect -6961 8727 -6927 8761
rect -6893 8727 -6859 8761
rect -6703 8727 -6669 8761
rect -6635 8727 -6601 8761
rect -6445 8727 -6411 8761
rect -6377 8727 -6343 8761
rect -6187 8727 -6153 8761
rect -6119 8727 -6085 8761
rect -5929 8727 -5895 8761
rect -5861 8727 -5827 8761
rect -5671 8727 -5637 8761
rect -5603 8727 -5569 8761
rect -5413 8727 -5379 8761
rect -5345 8727 -5311 8761
rect -5155 8727 -5121 8761
rect -5087 8727 -5053 8761
rect -4897 8727 -4863 8761
rect -4829 8727 -4795 8761
rect -7685 7576 -7651 7610
rect -7617 7576 -7583 7610
rect -7427 7576 -7393 7610
rect -7359 7576 -7325 7610
rect -7169 7576 -7135 7610
rect -7101 7576 -7067 7610
rect -6911 7576 -6877 7610
rect -6843 7576 -6809 7610
rect -6653 7576 -6619 7610
rect -6585 7576 -6551 7610
rect -6395 7576 -6361 7610
rect -6327 7576 -6293 7610
rect -6137 7576 -6103 7610
rect -6069 7576 -6035 7610
rect -5879 7576 -5845 7610
rect -5811 7576 -5777 7610
rect -5621 7576 -5587 7610
rect -5553 7576 -5519 7610
rect -5363 7576 -5329 7610
rect -5295 7576 -5261 7610
rect -5105 7576 -5071 7610
rect -5037 7576 -5003 7610
rect -4847 7576 -4813 7610
rect -4779 7576 -4745 7610
rect -4589 7576 -4555 7610
rect -4521 7576 -4487 7610
rect -4331 7576 -4297 7610
rect -4263 7576 -4229 7610
rect -4073 7576 -4039 7610
rect -4005 7576 -3971 7610
rect -3815 7576 -3781 7610
rect -3747 7576 -3713 7610
rect 15041 8166 15075 8200
rect 15109 8166 15143 8200
rect 15177 8166 15211 8200
rect 15245 8166 15279 8200
rect 15313 8166 15347 8200
rect 15381 8166 15415 8200
rect 15449 8166 15483 8200
rect 15517 8166 15551 8200
rect 15585 8166 15619 8200
rect 15653 8166 15687 8200
rect 15721 8166 15755 8200
rect 15789 8166 15823 8200
rect 15857 8166 15891 8200
rect 15925 8166 15959 8200
rect 16099 8166 16133 8200
rect 16167 8166 16201 8200
rect 16235 8166 16269 8200
rect 16303 8166 16337 8200
rect 16371 8166 16405 8200
rect 16439 8166 16473 8200
rect 16507 8166 16541 8200
rect 16575 8166 16609 8200
rect 16643 8166 16677 8200
rect 16711 8166 16745 8200
rect 16779 8166 16813 8200
rect 16847 8166 16881 8200
rect 16915 8166 16949 8200
rect 16983 8166 17017 8200
rect 17565 11268 17599 11302
rect 17633 11268 17667 11302
rect 17701 11268 17735 11302
rect 17769 11268 17803 11302
rect 17837 11268 17871 11302
rect 17905 11268 17939 11302
rect 17973 11268 18007 11302
rect 18041 11268 18075 11302
rect 18109 11268 18143 11302
rect 18177 11268 18211 11302
rect 18245 11268 18279 11302
rect 18313 11268 18347 11302
rect 18381 11268 18415 11302
rect 18449 11268 18483 11302
rect 18623 11268 18657 11302
rect 18691 11268 18725 11302
rect 18759 11268 18793 11302
rect 18827 11268 18861 11302
rect 18895 11268 18929 11302
rect 18963 11268 18997 11302
rect 19031 11268 19065 11302
rect 19099 11268 19133 11302
rect 19167 11268 19201 11302
rect 19235 11268 19269 11302
rect 19303 11268 19337 11302
rect 19371 11268 19405 11302
rect 19439 11268 19473 11302
rect 19507 11268 19541 11302
rect 17565 8140 17599 8174
rect 17633 8140 17667 8174
rect 17701 8140 17735 8174
rect 17769 8140 17803 8174
rect 17837 8140 17871 8174
rect 17905 8140 17939 8174
rect 17973 8140 18007 8174
rect 18041 8140 18075 8174
rect 18109 8140 18143 8174
rect 18177 8140 18211 8174
rect 18245 8140 18279 8174
rect 18313 8140 18347 8174
rect 18381 8140 18415 8174
rect 18449 8140 18483 8174
rect 18623 8140 18657 8174
rect 18691 8140 18725 8174
rect 18759 8140 18793 8174
rect 18827 8140 18861 8174
rect 18895 8140 18929 8174
rect 18963 8140 18997 8174
rect 19031 8140 19065 8174
rect 19099 8140 19133 8174
rect 19167 8140 19201 8174
rect 19235 8140 19269 8174
rect 19303 8140 19337 8174
rect 19371 8140 19405 8174
rect 19439 8140 19473 8174
rect 19507 8140 19541 8174
rect 17521 7586 17555 7620
rect 17589 7586 17623 7620
rect 17657 7586 17691 7620
rect 17725 7586 17759 7620
rect 17793 7586 17827 7620
rect 17861 7586 17895 7620
rect 17929 7586 17963 7620
rect 17997 7586 18031 7620
rect 18065 7586 18099 7620
rect 18133 7586 18167 7620
rect 18201 7586 18235 7620
rect 18269 7586 18303 7620
rect 18337 7586 18371 7620
rect 18405 7586 18439 7620
rect -7685 5466 -7651 5500
rect -7617 5466 -7583 5500
rect -7427 5466 -7393 5500
rect -7359 5466 -7325 5500
rect -7169 5466 -7135 5500
rect -7101 5466 -7067 5500
rect -6911 5466 -6877 5500
rect -6843 5466 -6809 5500
rect -6653 5466 -6619 5500
rect -6585 5466 -6551 5500
rect -6395 5466 -6361 5500
rect -6327 5466 -6293 5500
rect -6137 5466 -6103 5500
rect -6069 5466 -6035 5500
rect -5879 5466 -5845 5500
rect -5811 5466 -5777 5500
rect -5621 5466 -5587 5500
rect -5553 5466 -5519 5500
rect -5363 5466 -5329 5500
rect -5295 5466 -5261 5500
rect -5105 5466 -5071 5500
rect -5037 5466 -5003 5500
rect -4847 5466 -4813 5500
rect -4779 5466 -4745 5500
rect -4589 5466 -4555 5500
rect -4521 5466 -4487 5500
rect -4331 5466 -4297 5500
rect -4263 5466 -4229 5500
rect -4073 5466 -4039 5500
rect -4005 5466 -3971 5500
rect -3815 5466 -3781 5500
rect -3747 5466 -3713 5500
rect 17521 4476 17555 4510
rect 17589 4476 17623 4510
rect 17657 4476 17691 4510
rect 17725 4476 17759 4510
rect 17793 4476 17827 4510
rect 17861 4476 17895 4510
rect 17929 4476 17963 4510
rect 17997 4476 18031 4510
rect 18065 4476 18099 4510
rect 18133 4476 18167 4510
rect 18201 4476 18235 4510
rect 18269 4476 18303 4510
rect 18337 4476 18371 4510
rect 18405 4476 18439 4510
rect 18971 7586 19005 7620
rect 19039 7586 19073 7620
rect 19107 7586 19141 7620
rect 19175 7586 19209 7620
rect 19243 7586 19277 7620
rect 19311 7586 19345 7620
rect 19379 7586 19413 7620
rect 19447 7586 19481 7620
rect 19515 7586 19549 7620
rect 19583 7586 19617 7620
rect 19651 7586 19685 7620
rect 19719 7586 19753 7620
rect 19787 7586 19821 7620
rect 19855 7586 19889 7620
rect 23128 13235 23162 13269
rect 23128 13167 23162 13201
rect 23128 13099 23162 13133
rect 23128 13031 23162 13065
rect 23128 12963 23162 12997
rect 23128 12895 23162 12929
rect 23128 12827 23162 12861
rect 23128 12759 23162 12793
rect 23128 12691 23162 12725
rect 23128 12623 23162 12657
rect 23128 12555 23162 12589
rect 23128 12487 23162 12521
rect 23128 12419 23162 12453
rect 23128 12351 23162 12385
rect 24256 13235 24290 13269
rect 24256 13167 24290 13201
rect 24256 13099 24290 13133
rect 24256 13031 24290 13065
rect 24256 12963 24290 12997
rect 24256 12895 24290 12929
rect 24256 12827 24290 12861
rect 24256 12759 24290 12793
rect 24256 12691 24290 12725
rect 24256 12623 24290 12657
rect 24256 12555 24290 12589
rect 24256 12487 24290 12521
rect 24256 12419 24290 12453
rect 24256 12351 24290 12385
rect 24688 13229 24722 13263
rect 24688 13161 24722 13195
rect 24688 13093 24722 13127
rect 24688 13025 24722 13059
rect 24688 12957 24722 12991
rect 24688 12889 24722 12923
rect 24688 12821 24722 12855
rect 24688 12753 24722 12787
rect 24688 12685 24722 12719
rect 24688 12617 24722 12651
rect 24688 12549 24722 12583
rect 24688 12481 24722 12515
rect 24688 12413 24722 12447
rect 24688 12345 24722 12379
rect 25816 13229 25850 13263
rect 25816 13161 25850 13195
rect 25816 13093 25850 13127
rect 25816 13025 25850 13059
rect 25816 12957 25850 12991
rect 25816 12889 25850 12923
rect 25816 12821 25850 12855
rect 25816 12753 25850 12787
rect 25816 12685 25850 12719
rect 25816 12617 25850 12651
rect 25816 12549 25850 12583
rect 25816 12481 25850 12515
rect 25816 12413 25850 12447
rect 25816 12345 25850 12379
rect 23058 11695 23092 11729
rect 23058 11627 23092 11661
rect 23058 11559 23092 11593
rect 23058 11491 23092 11525
rect 23058 11423 23092 11457
rect 23058 11355 23092 11389
rect 23058 11287 23092 11321
rect 23058 11219 23092 11253
rect 23058 11151 23092 11185
rect 23058 11083 23092 11117
rect 23058 11015 23092 11049
rect 23058 10947 23092 10981
rect 23058 10879 23092 10913
rect 23058 10811 23092 10845
rect 24168 11695 24202 11729
rect 24168 11627 24202 11661
rect 24168 11559 24202 11593
rect 24168 11491 24202 11525
rect 24168 11423 24202 11457
rect 24168 11355 24202 11389
rect 24168 11287 24202 11321
rect 24168 11219 24202 11253
rect 24168 11151 24202 11185
rect 24168 11083 24202 11117
rect 24168 11015 24202 11049
rect 24168 10947 24202 10981
rect 24168 10879 24202 10913
rect 24168 10811 24202 10845
rect 24688 12171 24722 12205
rect 24688 12103 24722 12137
rect 24688 12035 24722 12069
rect 24688 11967 24722 12001
rect 24688 11899 24722 11933
rect 24688 11831 24722 11865
rect 24688 11763 24722 11797
rect 24688 11695 24722 11729
rect 24688 11627 24722 11661
rect 24688 11559 24722 11593
rect 24688 11491 24722 11525
rect 24688 11423 24722 11457
rect 24688 11355 24722 11389
rect 24688 11287 24722 11321
rect 25816 12171 25850 12205
rect 25816 12103 25850 12137
rect 25816 12035 25850 12069
rect 25816 11967 25850 12001
rect 25816 11899 25850 11933
rect 25816 11831 25850 11865
rect 25816 11763 25850 11797
rect 25816 11695 25850 11729
rect 25816 11627 25850 11661
rect 25816 11559 25850 11593
rect 25816 11491 25850 11525
rect 25816 11423 25850 11457
rect 25816 11355 25850 11389
rect 25816 11287 25850 11321
rect 24688 11113 24722 11147
rect 24688 11045 24722 11079
rect 24688 10977 24722 11011
rect 24688 10909 24722 10943
rect 24688 10841 24722 10875
rect 24688 10773 24722 10807
rect 24688 10705 24722 10739
rect 24688 10637 24722 10671
rect 24688 10569 24722 10603
rect 24688 10501 24722 10535
rect 24688 10433 24722 10467
rect 24688 10365 24722 10399
rect 24688 10297 24722 10331
rect 24688 10229 24722 10263
rect 25816 11113 25850 11147
rect 25816 11045 25850 11079
rect 25816 10977 25850 11011
rect 25816 10909 25850 10943
rect 25816 10841 25850 10875
rect 25816 10773 25850 10807
rect 25816 10705 25850 10739
rect 25816 10637 25850 10671
rect 25816 10569 25850 10603
rect 25816 10501 25850 10535
rect 25816 10433 25850 10467
rect 25816 10365 25850 10399
rect 25816 10297 25850 10331
rect 25816 10229 25850 10263
rect 24688 10055 24722 10089
rect 24688 9987 24722 10021
rect 24688 9919 24722 9953
rect 24688 9851 24722 9885
rect 24688 9783 24722 9817
rect 24688 9715 24722 9749
rect 24688 9647 24722 9681
rect 24688 9579 24722 9613
rect 24688 9511 24722 9545
rect 24688 9443 24722 9477
rect 24688 9375 24722 9409
rect 24688 9307 24722 9341
rect 24688 9239 24722 9273
rect 24688 9171 24722 9205
rect 25816 10055 25850 10089
rect 25816 9987 25850 10021
rect 25816 9919 25850 9953
rect 25816 9851 25850 9885
rect 25816 9783 25850 9817
rect 25816 9715 25850 9749
rect 25816 9647 25850 9681
rect 25816 9579 25850 9613
rect 25816 9511 25850 9545
rect 25816 9443 25850 9477
rect 25816 9375 25850 9409
rect 25816 9307 25850 9341
rect 25816 9239 25850 9273
rect 25816 9171 25850 9205
rect 23538 7759 23572 7793
rect 23538 7691 23572 7725
rect 23538 7623 23572 7657
rect 23538 7555 23572 7589
rect 23538 7487 23572 7521
rect 23538 7419 23572 7453
rect 23538 7351 23572 7385
rect 23538 7283 23572 7317
rect 23538 7215 23572 7249
rect 23538 7147 23572 7181
rect 23538 7079 23572 7113
rect 23538 7011 23572 7045
rect 23538 6943 23572 6977
rect 23538 6875 23572 6909
rect 24648 7759 24682 7793
rect 24648 7691 24682 7725
rect 24648 7623 24682 7657
rect 24648 7555 24682 7589
rect 24648 7487 24682 7521
rect 24648 7419 24682 7453
rect 24648 7351 24682 7385
rect 24648 7283 24682 7317
rect 24648 7215 24682 7249
rect 24648 7147 24682 7181
rect 24648 7079 24682 7113
rect 24648 7011 24682 7045
rect 24648 6943 24682 6977
rect 24648 6875 24682 6909
rect 23538 6701 23572 6735
rect 23538 6633 23572 6667
rect 23538 6565 23572 6599
rect 23538 6497 23572 6531
rect 23538 6429 23572 6463
rect 23538 6361 23572 6395
rect 23538 6293 23572 6327
rect 23538 6225 23572 6259
rect 23538 6157 23572 6191
rect 23538 6089 23572 6123
rect 23538 6021 23572 6055
rect 23538 5953 23572 5987
rect 23538 5885 23572 5919
rect 23538 5817 23572 5851
rect 24648 6701 24682 6735
rect 24648 6633 24682 6667
rect 24648 6565 24682 6599
rect 24648 6497 24682 6531
rect 24648 6429 24682 6463
rect 24648 6361 24682 6395
rect 24648 6293 24682 6327
rect 24648 6225 24682 6259
rect 24648 6157 24682 6191
rect 24648 6089 24682 6123
rect 24648 6021 24682 6055
rect 24648 5953 24682 5987
rect 24648 5885 24682 5919
rect 24648 5817 24682 5851
rect 23538 5643 23572 5677
rect 23538 5575 23572 5609
rect 23538 5507 23572 5541
rect 23538 5439 23572 5473
rect 23538 5371 23572 5405
rect 23538 5303 23572 5337
rect 23538 5235 23572 5269
rect 23538 5167 23572 5201
rect 23538 5099 23572 5133
rect 23538 5031 23572 5065
rect 23538 4963 23572 4997
rect 23538 4895 23572 4929
rect 23538 4827 23572 4861
rect 23538 4759 23572 4793
rect 24648 5643 24682 5677
rect 24648 5575 24682 5609
rect 24648 5507 24682 5541
rect 24648 5439 24682 5473
rect 24648 5371 24682 5405
rect 24648 5303 24682 5337
rect 24648 5235 24682 5269
rect 24648 5167 24682 5201
rect 24648 5099 24682 5133
rect 24648 5031 24682 5065
rect 24648 4963 24682 4997
rect 24648 4895 24682 4929
rect 24648 4827 24682 4861
rect 24648 4759 24682 4793
rect 18971 4476 19005 4510
rect 19039 4476 19073 4510
rect 19107 4476 19141 4510
rect 19175 4476 19209 4510
rect 19243 4476 19277 4510
rect 19311 4476 19345 4510
rect 19379 4476 19413 4510
rect 19447 4476 19481 4510
rect 19515 4476 19549 4510
rect 19583 4476 19617 4510
rect 19651 4476 19685 4510
rect 19719 4476 19753 4510
rect 19787 4476 19821 4510
rect 19855 4476 19889 4510
rect 23538 4585 23572 4619
rect 23538 4517 23572 4551
rect 23538 4449 23572 4483
rect 23538 4381 23572 4415
rect 23538 4313 23572 4347
rect 23538 4245 23572 4279
rect 23538 4177 23572 4211
rect 23538 4109 23572 4143
rect 23538 4041 23572 4075
rect 23538 3973 23572 4007
rect 23538 3905 23572 3939
rect 23538 3837 23572 3871
rect 23538 3769 23572 3803
rect 23538 3701 23572 3735
rect 24648 4585 24682 4619
rect 24648 4517 24682 4551
rect 24648 4449 24682 4483
rect 24648 4381 24682 4415
rect 24648 4313 24682 4347
rect 24648 4245 24682 4279
rect 24648 4177 24682 4211
rect 24648 4109 24682 4143
rect 24648 4041 24682 4075
rect 24648 3973 24682 4007
rect 24648 3905 24682 3939
rect 24648 3837 24682 3871
rect 24648 3769 24682 3803
rect 24648 3701 24682 3735
rect 25038 7759 25072 7793
rect 25038 7691 25072 7725
rect 25038 7623 25072 7657
rect 25038 7555 25072 7589
rect 25038 7487 25072 7521
rect 25038 7419 25072 7453
rect 25038 7351 25072 7385
rect 25038 7283 25072 7317
rect 25038 7215 25072 7249
rect 25038 7147 25072 7181
rect 25038 7079 25072 7113
rect 25038 7011 25072 7045
rect 25038 6943 25072 6977
rect 25038 6875 25072 6909
rect 26148 7759 26182 7793
rect 26148 7691 26182 7725
rect 26148 7623 26182 7657
rect 26148 7555 26182 7589
rect 26148 7487 26182 7521
rect 26148 7419 26182 7453
rect 26148 7351 26182 7385
rect 26148 7283 26182 7317
rect 26148 7215 26182 7249
rect 26148 7147 26182 7181
rect 26148 7079 26182 7113
rect 26148 7011 26182 7045
rect 26148 6943 26182 6977
rect 26148 6875 26182 6909
rect 25038 6701 25072 6735
rect 25038 6633 25072 6667
rect 25038 6565 25072 6599
rect 25038 6497 25072 6531
rect 25038 6429 25072 6463
rect 25038 6361 25072 6395
rect 25038 6293 25072 6327
rect 25038 6225 25072 6259
rect 25038 6157 25072 6191
rect 25038 6089 25072 6123
rect 25038 6021 25072 6055
rect 25038 5953 25072 5987
rect 25038 5885 25072 5919
rect 25038 5817 25072 5851
rect 26148 6701 26182 6735
rect 26148 6633 26182 6667
rect 26148 6565 26182 6599
rect 26148 6497 26182 6531
rect 26148 6429 26182 6463
rect 26148 6361 26182 6395
rect 26148 6293 26182 6327
rect 26148 6225 26182 6259
rect 26148 6157 26182 6191
rect 26148 6089 26182 6123
rect 26148 6021 26182 6055
rect 26148 5953 26182 5987
rect 26148 5885 26182 5919
rect 26148 5817 26182 5851
rect 25038 5643 25072 5677
rect 25038 5575 25072 5609
rect 25038 5507 25072 5541
rect 25038 5439 25072 5473
rect 25038 5371 25072 5405
rect 25038 5303 25072 5337
rect 25038 5235 25072 5269
rect 25038 5167 25072 5201
rect 25038 5099 25072 5133
rect 25038 5031 25072 5065
rect 25038 4963 25072 4997
rect 25038 4895 25072 4929
rect 25038 4827 25072 4861
rect 25038 4759 25072 4793
rect 26148 5643 26182 5677
rect 26148 5575 26182 5609
rect 26148 5507 26182 5541
rect 26148 5439 26182 5473
rect 26148 5371 26182 5405
rect 26148 5303 26182 5337
rect 26148 5235 26182 5269
rect 26148 5167 26182 5201
rect 26148 5099 26182 5133
rect 26148 5031 26182 5065
rect 26148 4963 26182 4997
rect 26148 4895 26182 4929
rect 26148 4827 26182 4861
rect 26148 4759 26182 4793
rect 25038 4585 25072 4619
rect 25038 4517 25072 4551
rect 25038 4449 25072 4483
rect 25038 4381 25072 4415
rect 25038 4313 25072 4347
rect 25038 4245 25072 4279
rect 25038 4177 25072 4211
rect 25038 4109 25072 4143
rect 25038 4041 25072 4075
rect 25038 3973 25072 4007
rect 25038 3905 25072 3939
rect 25038 3837 25072 3871
rect 25038 3769 25072 3803
rect 25038 3701 25072 3735
rect 26148 4585 26182 4619
rect 26148 4517 26182 4551
rect 26148 4449 26182 4483
rect 26148 4381 26182 4415
rect 26148 4313 26182 4347
rect 26148 4245 26182 4279
rect 26148 4177 26182 4211
rect 26148 4109 26182 4143
rect 26148 4041 26182 4075
rect 26148 3973 26182 4007
rect 26148 3905 26182 3939
rect 26148 3837 26182 3871
rect 26148 3769 26182 3803
rect 26148 3701 26182 3735
rect 38249 13437 38283 13471
rect 39045 13445 39079 13479
rect 39282 13440 39316 13474
rect 40076 13442 40110 13476
rect 40331 13442 40365 13476
rect 36872 11952 36906 11986
rect 36940 11952 36974 11986
rect 37130 11952 37164 11986
rect 37198 11952 37232 11986
rect 37388 11952 37422 11986
rect 37456 11952 37490 11986
rect 37646 11952 37680 11986
rect 37714 11952 37748 11986
rect 37904 11952 37938 11986
rect 37972 11952 38006 11986
rect 38162 11952 38196 11986
rect 38230 11952 38264 11986
rect 38420 11952 38454 11986
rect 38488 11952 38522 11986
rect 38678 11952 38712 11986
rect 38746 11952 38780 11986
rect 38936 11952 38970 11986
rect 39004 11952 39038 11986
rect 39194 11952 39228 11986
rect 39262 11952 39296 11986
rect 39452 11952 39486 11986
rect 39520 11952 39554 11986
rect 39710 11952 39744 11986
rect 39778 11952 39812 11986
rect 39968 11952 40002 11986
rect 40036 11952 40070 11986
rect 40226 11952 40260 11986
rect 40294 11952 40328 11986
rect 40484 11952 40518 11986
rect 40552 11952 40586 11986
rect 40742 11952 40776 11986
rect 40810 11952 40844 11986
rect 41000 11952 41034 11986
rect 41068 11952 41102 11986
rect 41258 11952 41292 11986
rect 41326 11952 41360 11986
rect 41516 11952 41550 11986
rect 41584 11952 41618 11986
rect 41774 11952 41808 11986
rect 41842 11952 41876 11986
rect 36872 10842 36906 10876
rect 36940 10842 36974 10876
rect 37130 10842 37164 10876
rect 37198 10842 37232 10876
rect 37388 10842 37422 10876
rect 37456 10842 37490 10876
rect 37646 10842 37680 10876
rect 37714 10842 37748 10876
rect 37904 10842 37938 10876
rect 37972 10842 38006 10876
rect 38162 10842 38196 10876
rect 38230 10842 38264 10876
rect 38420 10842 38454 10876
rect 38488 10842 38522 10876
rect 38678 10842 38712 10876
rect 38746 10842 38780 10876
rect 38936 10842 38970 10876
rect 39004 10842 39038 10876
rect 39194 10842 39228 10876
rect 39262 10842 39296 10876
rect 39452 10842 39486 10876
rect 39520 10842 39554 10876
rect 39710 10842 39744 10876
rect 39778 10842 39812 10876
rect 39968 10842 40002 10876
rect 40036 10842 40070 10876
rect 40226 10842 40260 10876
rect 40294 10842 40328 10876
rect 40484 10842 40518 10876
rect 40552 10842 40586 10876
rect 40742 10842 40776 10876
rect 40810 10842 40844 10876
rect 41000 10842 41034 10876
rect 41068 10842 41102 10876
rect 41258 10842 41292 10876
rect 41326 10842 41360 10876
rect 41516 10842 41550 10876
rect 41584 10842 41618 10876
rect 41774 10842 41808 10876
rect 41842 10842 41876 10876
rect 37907 10587 37941 10621
rect 37975 10587 38009 10621
rect 38373 10587 38407 10621
rect 38441 10587 38475 10621
rect 38631 10587 38665 10621
rect 38699 10587 38733 10621
rect 38889 10587 38923 10621
rect 38957 10587 38991 10621
rect 39147 10587 39181 10621
rect 39215 10587 39249 10621
rect 39405 10587 39439 10621
rect 39473 10587 39507 10621
rect 39663 10587 39697 10621
rect 39731 10587 39765 10621
rect 39921 10587 39955 10621
rect 39989 10587 40023 10621
rect 40179 10587 40213 10621
rect 40247 10587 40281 10621
rect 40437 10587 40471 10621
rect 40505 10587 40539 10621
rect 40695 10587 40729 10621
rect 40763 10587 40797 10621
rect 37907 9477 37941 9511
rect 37975 9477 38009 9511
rect 38373 9477 38407 9511
rect 38441 9477 38475 9511
rect 38631 9477 38665 9511
rect 38699 9477 38733 9511
rect 38889 9477 38923 9511
rect 38957 9477 38991 9511
rect 39147 9477 39181 9511
rect 39215 9477 39249 9511
rect 39405 9477 39439 9511
rect 39473 9477 39507 9511
rect 39663 9477 39697 9511
rect 39731 9477 39765 9511
rect 39921 9477 39955 9511
rect 39989 9477 40023 9511
rect 40179 9477 40213 9511
rect 40247 9477 40281 9511
rect 40437 9477 40471 9511
rect 40505 9477 40539 9511
rect 40695 9477 40729 9511
rect 40763 9477 40797 9511
rect 37907 8326 37941 8360
rect 37975 8326 38009 8360
rect 38165 8326 38199 8360
rect 38233 8326 38267 8360
rect 38423 8326 38457 8360
rect 38491 8326 38525 8360
rect 38681 8326 38715 8360
rect 38749 8326 38783 8360
rect 38939 8326 38973 8360
rect 39007 8326 39041 8360
rect 39197 8326 39231 8360
rect 39265 8326 39299 8360
rect 39455 8326 39489 8360
rect 39523 8326 39557 8360
rect 39713 8326 39747 8360
rect 39781 8326 39815 8360
rect 39971 8326 40005 8360
rect 40039 8326 40073 8360
rect 40229 8326 40263 8360
rect 40297 8326 40331 8360
rect 40487 8326 40521 8360
rect 40555 8326 40589 8360
rect 40745 8326 40779 8360
rect 40813 8326 40847 8360
rect 41003 8326 41037 8360
rect 41071 8326 41105 8360
rect 41261 8326 41295 8360
rect 41329 8326 41363 8360
rect 41519 8326 41553 8360
rect 41587 8326 41621 8360
rect 41777 8326 41811 8360
rect 41845 8326 41879 8360
rect 37907 6216 37941 6250
rect 37975 6216 38009 6250
rect 38165 6216 38199 6250
rect 38233 6216 38267 6250
rect 38423 6216 38457 6250
rect 38491 6216 38525 6250
rect 38681 6216 38715 6250
rect 38749 6216 38783 6250
rect 38939 6216 38973 6250
rect 39007 6216 39041 6250
rect 39197 6216 39231 6250
rect 39265 6216 39299 6250
rect 39455 6216 39489 6250
rect 39523 6216 39557 6250
rect 39713 6216 39747 6250
rect 39781 6216 39815 6250
rect 39971 6216 40005 6250
rect 40039 6216 40073 6250
rect 40229 6216 40263 6250
rect 40297 6216 40331 6250
rect 40487 6216 40521 6250
rect 40555 6216 40589 6250
rect 40745 6216 40779 6250
rect 40813 6216 40847 6250
rect 41003 6216 41037 6250
rect 41071 6216 41105 6250
rect 41261 6216 41295 6250
rect 41329 6216 41363 6250
rect 41519 6216 41553 6250
rect 41587 6216 41621 6250
rect 41777 6216 41811 6250
rect 41845 6216 41879 6250
<< xpolycontact >>
rect 24590 16550 25022 16620
rect 27122 16550 27554 16620
rect 24590 16232 25022 16302
rect 27122 16232 27554 16302
rect 24590 15914 25022 15984
rect 27122 15914 27554 15984
rect -3880 14473 -3810 14905
rect -3880 12441 -3810 12873
rect 24590 15596 25022 15666
rect 27122 15596 27554 15666
rect 24590 15278 25022 15348
rect 27122 15278 27554 15348
rect 16210 6678 16280 7110
rect 16210 4646 16280 5078
rect 16528 6678 16598 7110
rect 16528 4646 16598 5078
rect 16846 6678 16916 7110
rect 16846 4646 16916 5078
rect 20512 14038 20582 14470
rect 20512 4720 20582 5152
rect 20830 14038 20900 14470
rect 20830 4720 20900 5152
rect 21148 14038 21218 14470
rect 21148 4720 21218 5152
rect 21466 14038 21536 14470
rect 21466 4720 21536 5152
rect 28964 14830 29034 15262
rect 28964 13758 29034 14190
rect 29282 14830 29352 15262
rect 29282 13758 29352 14190
rect 29600 14830 29670 15262
rect 29600 13758 29670 14190
rect 26528 12912 26598 13344
rect 26528 3080 26598 3512
rect 26846 12912 26916 13344
rect 26846 3080 26916 3512
rect 27164 12912 27234 13344
rect 27164 3080 27234 3512
rect 27700 12896 27770 13328
rect 27700 6464 27770 6896
rect 28018 12896 28088 13328
rect 28018 6464 28088 6896
rect 28336 12896 28406 13328
rect 28336 6464 28406 6896
rect 28654 12896 28724 13328
rect 28654 6464 28724 6896
rect 28972 12896 29042 13328
rect 28972 6464 29042 6896
rect 29290 12896 29360 13328
rect 29290 6464 29360 6896
rect 29608 12896 29678 13328
rect 29608 6464 29678 6896
rect 41712 15223 41782 15655
rect 41712 13191 41782 13623
<< ppolyres >>
rect 25022 16550 27122 16620
rect 25022 16232 27122 16302
rect 25022 15914 27122 15984
rect -3880 12873 -3810 14473
rect 25022 15596 27122 15666
rect 25022 15278 27122 15348
rect 16210 5078 16280 6678
rect 16528 5078 16598 6678
rect 16846 5078 16916 6678
rect 20512 5152 20582 14038
rect 20830 5152 20900 14038
rect 21148 5152 21218 14038
rect 21466 5152 21536 14038
rect 28964 14190 29034 14830
rect 29282 14190 29352 14830
rect 29600 14190 29670 14830
rect 26528 3512 26598 12912
rect 26846 3512 26916 12912
rect 27164 3512 27234 12912
rect 27700 6896 27770 12896
rect 28018 6896 28088 12896
rect 28336 6896 28406 12896
rect 28654 6896 28724 12896
rect 28972 6896 29042 12896
rect 29290 6896 29360 12896
rect 29608 6896 29678 12896
rect 41712 13623 41782 15223
<< locali >>
rect 41308 22935 42036 22951
rect -4284 22185 -3556 22201
rect -4284 21359 -4261 22185
rect -3579 21359 -3556 22185
rect 41308 22109 41331 22935
rect 42013 22109 42036 22935
rect 41308 22093 42036 22109
rect -4284 21343 -3556 21359
rect 42341 19247 45374 19253
rect 40682 19215 45374 19247
rect 40682 19037 41520 19215
rect 41770 19199 45374 19215
rect 41770 19093 43604 19199
rect 43710 19093 45374 19199
rect 41770 19062 45374 19093
rect 41770 19037 42576 19062
rect 40682 19028 42576 19037
rect 42610 19028 42644 19062
rect 42678 19028 42712 19062
rect 42746 19028 42780 19062
rect 42814 19028 42848 19062
rect 42882 19028 42916 19062
rect 42950 19028 42984 19062
rect 43018 19028 43052 19062
rect 43086 19028 43120 19062
rect 43154 19028 43188 19062
rect 43222 19028 43256 19062
rect 43290 19028 43324 19062
rect 43358 19028 43392 19062
rect 43426 19028 43460 19062
rect 43494 19028 43528 19062
rect 43562 19028 43596 19062
rect 43630 19028 43664 19062
rect 43698 19028 43732 19062
rect 43766 19028 43800 19062
rect 43834 19028 43868 19062
rect 43902 19028 43936 19062
rect 43970 19028 44004 19062
rect 44038 19028 44072 19062
rect 44106 19028 44140 19062
rect 44174 19028 44208 19062
rect 44242 19028 44276 19062
rect 44310 19028 44344 19062
rect 44378 19028 44412 19062
rect 44446 19028 44480 19062
rect 44514 19028 44548 19062
rect 44582 19028 44616 19062
rect 44650 19028 44684 19062
rect 44718 19028 44752 19062
rect 44786 19028 44820 19062
rect 44854 19028 44888 19062
rect 44922 19028 44956 19062
rect 44990 19028 45024 19062
rect 45058 19028 45092 19062
rect 45126 19028 45160 19062
rect 45194 19028 45228 19062
rect 45262 19028 45374 19062
rect 40682 19006 45374 19028
rect 23042 18932 23161 18966
rect 23195 18932 23229 18966
rect 23263 18932 23297 18966
rect 23331 18932 23365 18966
rect 23399 18932 23433 18966
rect 23467 18932 23501 18966
rect 23535 18932 23569 18966
rect 23603 18932 23637 18966
rect 23671 18932 23705 18966
rect 23739 18932 23773 18966
rect 23807 18932 23841 18966
rect 23875 18932 23909 18966
rect 23943 18932 23977 18966
rect 24011 18932 24045 18966
rect 24079 18932 24113 18966
rect 24147 18932 24181 18966
rect 24215 18932 24249 18966
rect 24283 18932 24402 18966
rect 23042 18842 23076 18932
rect 24368 18842 24402 18932
rect 23042 18774 23076 18808
rect 23222 18794 23263 18828
rect 23307 18794 23331 18828
rect 23379 18794 23399 18828
rect 23451 18794 23467 18828
rect 23523 18794 23535 18828
rect 23595 18794 23603 18828
rect 23667 18794 23671 18828
rect 23773 18794 23777 18828
rect 23841 18794 23849 18828
rect 23909 18794 23921 18828
rect 23977 18794 23993 18828
rect 24045 18794 24065 18828
rect 24113 18794 24137 18828
rect 24181 18794 24222 18828
rect 24368 18774 24402 18808
rect 23042 18706 23076 18740
rect 21862 18659 22482 18660
rect 23042 18659 23076 18672
rect 23176 18732 23210 18751
rect 23176 18660 23210 18672
rect 21862 18638 23176 18659
rect 24234 18732 24268 18751
rect 24234 18660 24268 18672
rect 21862 18604 23042 18638
rect 23076 18604 23176 18638
rect 23210 18604 23213 18659
rect 21862 18588 23213 18604
rect 21862 18570 23176 18588
rect 21862 18536 23042 18570
rect 23076 18536 23176 18570
rect 23210 18569 23213 18588
rect 24234 18588 24268 18604
rect 23210 18536 23222 18569
rect 21862 18516 23222 18536
rect -3251 18497 -218 18503
rect -4910 18465 -218 18497
rect -4910 18287 -4072 18465
rect -3822 18449 -218 18465
rect -3822 18343 -1988 18449
rect -1882 18343 -218 18449
rect -3822 18312 -218 18343
rect -3822 18287 -3016 18312
rect -4910 18278 -3016 18287
rect -2982 18278 -2948 18312
rect -2914 18278 -2880 18312
rect -2846 18278 -2812 18312
rect -2778 18278 -2744 18312
rect -2710 18278 -2676 18312
rect -2642 18278 -2608 18312
rect -2574 18278 -2540 18312
rect -2506 18278 -2472 18312
rect -2438 18278 -2404 18312
rect -2370 18278 -2336 18312
rect -2302 18278 -2268 18312
rect -2234 18278 -2200 18312
rect -2166 18278 -2132 18312
rect -2098 18278 -2064 18312
rect -2030 18278 -1996 18312
rect -1962 18278 -1928 18312
rect -1894 18278 -1860 18312
rect -1826 18278 -1792 18312
rect -1758 18278 -1724 18312
rect -1690 18278 -1656 18312
rect -1622 18278 -1588 18312
rect -1554 18278 -1520 18312
rect -1486 18278 -1452 18312
rect -1418 18278 -1384 18312
rect -1350 18278 -1316 18312
rect -1282 18278 -1248 18312
rect -1214 18278 -1180 18312
rect -1146 18278 -1112 18312
rect -1078 18278 -1044 18312
rect -1010 18278 -976 18312
rect -942 18278 -908 18312
rect -874 18278 -840 18312
rect -806 18278 -772 18312
rect -738 18278 -704 18312
rect -670 18278 -636 18312
rect -602 18278 -568 18312
rect -534 18278 -500 18312
rect -466 18278 -432 18312
rect -398 18278 -364 18312
rect -330 18278 -218 18312
rect -4910 18256 -218 18278
rect -4910 17785 -4669 18256
rect -3251 18253 -218 18256
rect 21862 18502 23176 18516
rect 21862 18468 23042 18502
rect 23076 18468 23176 18502
rect 23210 18468 23222 18516
rect 21862 18444 23222 18468
rect 21862 18434 23176 18444
rect 21862 18400 23042 18434
rect 23076 18400 23176 18434
rect 23210 18400 23222 18444
rect 21862 18387 23222 18400
rect 24234 18516 24268 18536
rect 24234 18444 24268 18468
rect 21862 18372 23213 18387
rect 21862 18366 23176 18372
rect 21862 18332 23042 18366
rect 23076 18332 23176 18366
rect 23210 18332 23213 18372
rect 21862 18300 23213 18332
rect 21862 18298 23176 18300
rect 21862 18264 23042 18298
rect 23076 18264 23176 18298
rect 23210 18264 23213 18300
rect -6817 17544 -4669 17785
rect -3114 18198 -3080 18253
rect -266 18198 -232 18253
rect -3114 18130 -3080 18164
rect -2934 18140 -2887 18174
rect -2851 18140 -2817 18174
rect -2781 18140 -2734 18174
rect -2676 18140 -2629 18174
rect -2593 18140 -2559 18174
rect -2523 18140 -2476 18174
rect -2418 18140 -2371 18174
rect -2335 18140 -2301 18174
rect -2265 18140 -2218 18174
rect -2160 18140 -2113 18174
rect -2077 18140 -2043 18174
rect -2007 18140 -1960 18174
rect -1902 18140 -1855 18174
rect -1819 18140 -1785 18174
rect -1749 18140 -1702 18174
rect -1644 18140 -1597 18174
rect -1561 18140 -1527 18174
rect -1491 18140 -1444 18174
rect -1386 18140 -1339 18174
rect -1303 18140 -1269 18174
rect -1233 18140 -1186 18174
rect -1128 18140 -1081 18174
rect -1045 18140 -1011 18174
rect -975 18140 -928 18174
rect -870 18140 -823 18174
rect -787 18140 -753 18174
rect -717 18140 -670 18174
rect -612 18140 -565 18174
rect -529 18140 -495 18174
rect -459 18140 -412 18174
rect -266 18130 -232 18164
rect -3114 18062 -3080 18096
rect -3114 17994 -3080 18028
rect -3114 17926 -3080 17960
rect -3114 17858 -3080 17892
rect -3114 17790 -3080 17824
rect -3114 17722 -3080 17756
rect -3114 17654 -3080 17688
rect -3114 17586 -3080 17620
rect -6817 17541 -5446 17544
rect -6817 17536 -6239 17541
rect -6205 17536 -6167 17541
rect -6133 17536 -5446 17541
rect -6817 17502 -6702 17536
rect -6668 17502 -6634 17536
rect -6600 17502 -6566 17536
rect -6532 17502 -6498 17536
rect -6464 17502 -6430 17536
rect -6396 17502 -6362 17536
rect -6328 17502 -6294 17536
rect -6260 17507 -6239 17536
rect -6192 17507 -6167 17536
rect -6260 17502 -6226 17507
rect -6192 17502 -6158 17507
rect -6124 17502 -6090 17536
rect -6056 17502 -6022 17536
rect -5988 17502 -5954 17536
rect -5920 17502 -5886 17536
rect -5852 17502 -5818 17536
rect -5784 17502 -5750 17536
rect -5716 17502 -5682 17536
rect -5648 17502 -5614 17536
rect -5580 17502 -5446 17536
rect -6817 17478 -5446 17502
rect -6816 17441 -6736 17478
rect -6276 17454 -6096 17478
rect -5526 17461 -5446 17478
rect -6816 17407 -6798 17441
rect -6764 17407 -6736 17441
rect -6816 17373 -6736 17407
rect -6816 17339 -6798 17373
rect -6764 17339 -6736 17373
rect -6816 17305 -6736 17339
rect -5526 17427 -5508 17461
rect -5474 17427 -5446 17461
rect -5526 17393 -5446 17427
rect -5526 17359 -5508 17393
rect -5474 17359 -5446 17393
rect -5526 17325 -5446 17359
rect -6816 17271 -6798 17305
rect -6764 17271 -6736 17305
rect -6402 17271 -6355 17305
rect -6319 17271 -6285 17305
rect -6249 17271 -6202 17305
rect -6144 17271 -6097 17305
rect -6061 17271 -6027 17305
rect -5991 17271 -5944 17305
rect -5526 17291 -5508 17325
rect -5474 17291 -5446 17325
rect -6816 17237 -6736 17271
rect -6816 17203 -6798 17237
rect -6764 17203 -6736 17237
rect -5526 17257 -5446 17291
rect -6816 17169 -6736 17203
rect -6816 17135 -6798 17169
rect -6764 17135 -6736 17169
rect -6816 17101 -6736 17135
rect -6816 17067 -6798 17101
rect -6764 17067 -6736 17101
rect -6816 17033 -6736 17067
rect -6816 16999 -6798 17033
rect -6764 16999 -6736 17033
rect -6816 16965 -6736 16999
rect -6816 16931 -6798 16965
rect -6764 16931 -6736 16965
rect -6816 16897 -6736 16931
rect -6816 16863 -6798 16897
rect -6764 16863 -6736 16897
rect -6816 16829 -6736 16863
rect -6816 16795 -6798 16829
rect -6764 16795 -6736 16829
rect -6816 16761 -6736 16795
rect -6816 16727 -6798 16761
rect -6764 16727 -6736 16761
rect -6816 16693 -6736 16727
rect -6816 16659 -6798 16693
rect -6764 16659 -6736 16693
rect -6816 16625 -6736 16659
rect -6816 16591 -6798 16625
rect -6764 16591 -6736 16625
rect -6816 16557 -6736 16591
rect -6816 16523 -6798 16557
rect -6764 16523 -6736 16557
rect -6816 16489 -6736 16523
rect -6816 16455 -6798 16489
rect -6764 16455 -6736 16489
rect -6816 16421 -6736 16455
rect -6816 16387 -6798 16421
rect -6764 16387 -6736 16421
rect -6816 16353 -6736 16387
rect -6816 16319 -6798 16353
rect -6764 16319 -6736 16353
rect -6816 16285 -6736 16319
rect -6816 16251 -6798 16285
rect -6764 16251 -6736 16285
rect -6816 16217 -6736 16251
rect -6448 17209 -6414 17228
rect -6448 17137 -6414 17149
rect -6448 17065 -6414 17081
rect -6448 16993 -6414 17013
rect -6448 16921 -6414 16945
rect -6448 16849 -6414 16877
rect -6448 16777 -6414 16809
rect -6448 16707 -6414 16741
rect -6448 16639 -6414 16671
rect -6448 16571 -6414 16599
rect -6448 16503 -6414 16527
rect -6448 16435 -6414 16455
rect -6448 16367 -6414 16383
rect -6448 16299 -6414 16311
rect -6448 16220 -6414 16239
rect -6190 17209 -6156 17228
rect -6190 17137 -6156 17149
rect -6190 17065 -6156 17081
rect -6190 16993 -6156 17013
rect -6190 16921 -6156 16945
rect -6190 16849 -6156 16877
rect -6190 16777 -6156 16809
rect -6190 16707 -6156 16741
rect -6190 16639 -6156 16671
rect -6190 16571 -6156 16599
rect -6190 16503 -6156 16527
rect -6190 16435 -6156 16455
rect -6190 16367 -6156 16383
rect -6190 16299 -6156 16311
rect -6190 16220 -6156 16239
rect -5932 17209 -5898 17228
rect -5932 17137 -5898 17149
rect -5932 17065 -5898 17081
rect -5932 16993 -5898 17013
rect -5932 16921 -5898 16945
rect -5932 16849 -5898 16877
rect -5932 16777 -5898 16809
rect -5932 16707 -5898 16741
rect -5932 16639 -5898 16671
rect -5932 16571 -5898 16599
rect -5932 16503 -5898 16527
rect -5932 16435 -5898 16455
rect -5932 16367 -5898 16383
rect -5932 16299 -5898 16311
rect -5932 16220 -5898 16239
rect -5526 17223 -5508 17257
rect -5474 17223 -5446 17257
rect -5526 17189 -5446 17223
rect -5526 17155 -5508 17189
rect -5474 17155 -5446 17189
rect -5526 17121 -5446 17155
rect -5526 17087 -5508 17121
rect -5474 17087 -5446 17121
rect -5526 17053 -5446 17087
rect -5526 17019 -5508 17053
rect -5474 17019 -5446 17053
rect -5526 16985 -5446 17019
rect -5526 16951 -5508 16985
rect -5474 16951 -5446 16985
rect -5526 16917 -5446 16951
rect -5526 16883 -5508 16917
rect -5474 16883 -5446 16917
rect -5526 16849 -5446 16883
rect -5526 16815 -5508 16849
rect -5474 16815 -5446 16849
rect -5526 16781 -5446 16815
rect -5526 16747 -5508 16781
rect -5474 16747 -5446 16781
rect -5526 16713 -5446 16747
rect -5526 16679 -5508 16713
rect -5474 16679 -5446 16713
rect -5526 16645 -5446 16679
rect -5526 16611 -5508 16645
rect -5474 16611 -5446 16645
rect -5526 16577 -5446 16611
rect -5526 16543 -5508 16577
rect -5474 16543 -5446 16577
rect -5526 16509 -5446 16543
rect -5526 16475 -5508 16509
rect -5474 16475 -5446 16509
rect -5526 16441 -5446 16475
rect -5526 16407 -5508 16441
rect -5474 16407 -5446 16441
rect -5526 16373 -5446 16407
rect -5526 16339 -5508 16373
rect -5474 16339 -5446 16373
rect -5526 16305 -5446 16339
rect -5526 16271 -5508 16305
rect -5474 16271 -5446 16305
rect -5526 16237 -5446 16271
rect -6816 16183 -6798 16217
rect -6764 16183 -6736 16217
rect -6816 16149 -6736 16183
rect -5526 16203 -5508 16237
rect -5474 16203 -5446 16237
rect -6816 16115 -6798 16149
rect -6764 16115 -6736 16149
rect -6402 16143 -6355 16177
rect -6319 16143 -6285 16177
rect -6249 16143 -6202 16177
rect -6144 16143 -6097 16177
rect -6061 16143 -6027 16177
rect -5991 16143 -5944 16177
rect -5526 16169 -5446 16203
rect -6816 16081 -6736 16115
rect -6816 16047 -6798 16081
rect -6764 16047 -6736 16081
rect -6816 16024 -6736 16047
rect -5526 16135 -5508 16169
rect -5474 16135 -5446 16169
rect -5526 16101 -5446 16135
rect -5526 16067 -5508 16101
rect -5474 16067 -5446 16101
rect -5526 16024 -5446 16067
rect -6816 15996 -5446 16024
rect -6816 15962 -6682 15996
rect -6648 15962 -6614 15996
rect -6580 15962 -6546 15996
rect -6512 15962 -6478 15996
rect -6444 15962 -6410 15996
rect -6376 15962 -6342 15996
rect -6308 15962 -6274 15996
rect -6240 15962 -6206 15996
rect -6172 15962 -6138 15996
rect -6104 15962 -6070 15996
rect -6036 15962 -6002 15996
rect -5968 15962 -5934 15996
rect -5900 15962 -5866 15996
rect -5832 15962 -5798 15996
rect -5764 15962 -5730 15996
rect -5696 15962 -5662 15996
rect -5628 15962 -5594 15996
rect -5560 15962 -5446 15996
rect -6816 15944 -5446 15962
rect -3114 17518 -3080 17552
rect -3114 17450 -3080 17484
rect -3114 17382 -3080 17416
rect -3114 17314 -3080 17348
rect -3114 17246 -3080 17280
rect -3114 17178 -3080 17212
rect -3114 17110 -3080 17144
rect -3114 17042 -3080 17076
rect -3114 16974 -3080 17008
rect -3114 16906 -3080 16940
rect -3114 16838 -3080 16872
rect -3114 16770 -3080 16804
rect -3114 16702 -3080 16736
rect -3114 16634 -3080 16668
rect -3114 16566 -3080 16600
rect -3114 16498 -3080 16532
rect -3114 16430 -3080 16464
rect -3114 16362 -3080 16396
rect -3114 16294 -3080 16328
rect -3114 16226 -3080 16260
rect -3114 16158 -3080 16192
rect -3114 16090 -3080 16124
rect -2980 18062 -2946 18097
rect -2980 17994 -2946 18012
rect -2980 17926 -2946 17940
rect -2980 17858 -2946 17868
rect -2980 17790 -2946 17796
rect -2980 17722 -2946 17724
rect -2980 17686 -2946 17688
rect -2980 17614 -2946 17620
rect -2980 17542 -2946 17552
rect -2980 17470 -2946 17484
rect -2980 17398 -2946 17416
rect -2980 17326 -2946 17348
rect -2980 17254 -2946 17280
rect -2980 17182 -2946 17212
rect -2980 17110 -2946 17144
rect -2980 17042 -2946 17076
rect -2980 16974 -2946 17004
rect -2980 16906 -2946 16932
rect -2980 16838 -2946 16860
rect -2980 16770 -2946 16788
rect -2980 16702 -2946 16716
rect -2980 16634 -2946 16644
rect -2980 16566 -2946 16572
rect -2980 16498 -2946 16500
rect -2980 16462 -2946 16464
rect -2980 16390 -2946 16396
rect -2980 16318 -2946 16328
rect -2980 16246 -2946 16260
rect -2980 16174 -2946 16192
rect -2980 16089 -2946 16124
rect -2722 18062 -2688 18097
rect -2722 17994 -2688 18012
rect -2722 17926 -2688 17940
rect -2722 17858 -2688 17868
rect -2722 17790 -2688 17796
rect -2722 17722 -2688 17724
rect -2722 17686 -2688 17688
rect -2722 17614 -2688 17620
rect -2722 17542 -2688 17552
rect -2722 17470 -2688 17484
rect -2722 17398 -2688 17416
rect -2722 17326 -2688 17348
rect -2722 17254 -2688 17280
rect -2722 17182 -2688 17212
rect -2722 17110 -2688 17144
rect -2722 17042 -2688 17076
rect -2722 16974 -2688 17004
rect -2722 16906 -2688 16932
rect -2722 16838 -2688 16860
rect -2722 16770 -2688 16788
rect -2722 16702 -2688 16716
rect -2722 16634 -2688 16644
rect -2722 16566 -2688 16572
rect -2722 16498 -2688 16500
rect -2722 16462 -2688 16464
rect -2722 16390 -2688 16396
rect -2722 16318 -2688 16328
rect -2722 16246 -2688 16260
rect -2722 16174 -2688 16192
rect -2722 16089 -2688 16124
rect -2464 18062 -2430 18097
rect -2464 17994 -2430 18012
rect -2464 17926 -2430 17940
rect -2464 17858 -2430 17868
rect -2464 17790 -2430 17796
rect -2464 17722 -2430 17724
rect -2464 17686 -2430 17688
rect -2464 17614 -2430 17620
rect -2464 17542 -2430 17552
rect -2464 17470 -2430 17484
rect -2464 17398 -2430 17416
rect -2464 17326 -2430 17348
rect -2464 17254 -2430 17280
rect -2464 17182 -2430 17212
rect -2464 17110 -2430 17144
rect -2464 17042 -2430 17076
rect -2464 16974 -2430 17004
rect -2464 16906 -2430 16932
rect -2464 16838 -2430 16860
rect -2464 16770 -2430 16788
rect -2464 16702 -2430 16716
rect -2464 16634 -2430 16644
rect -2464 16566 -2430 16572
rect -2464 16498 -2430 16500
rect -2464 16462 -2430 16464
rect -2464 16390 -2430 16396
rect -2464 16318 -2430 16328
rect -2464 16246 -2430 16260
rect -2464 16174 -2430 16192
rect -2464 16089 -2430 16124
rect -2206 18062 -2172 18097
rect -2206 17994 -2172 18012
rect -2206 17926 -2172 17940
rect -2206 17858 -2172 17868
rect -2206 17790 -2172 17796
rect -2206 17722 -2172 17724
rect -2206 17686 -2172 17688
rect -2206 17614 -2172 17620
rect -2206 17542 -2172 17552
rect -2206 17470 -2172 17484
rect -2206 17398 -2172 17416
rect -2206 17326 -2172 17348
rect -2206 17254 -2172 17280
rect -2206 17182 -2172 17212
rect -2206 17110 -2172 17144
rect -2206 17042 -2172 17076
rect -2206 16974 -2172 17004
rect -2206 16906 -2172 16932
rect -2206 16838 -2172 16860
rect -2206 16770 -2172 16788
rect -2206 16702 -2172 16716
rect -2206 16634 -2172 16644
rect -2206 16566 -2172 16572
rect -2206 16498 -2172 16500
rect -2206 16462 -2172 16464
rect -2206 16390 -2172 16396
rect -2206 16318 -2172 16328
rect -2206 16246 -2172 16260
rect -2206 16174 -2172 16192
rect -2206 16089 -2172 16124
rect -1948 18062 -1914 18097
rect -1948 17994 -1914 18012
rect -1948 17926 -1914 17940
rect -1948 17858 -1914 17868
rect -1948 17790 -1914 17796
rect -1948 17722 -1914 17724
rect -1948 17686 -1914 17688
rect -1948 17614 -1914 17620
rect -1948 17542 -1914 17552
rect -1948 17470 -1914 17484
rect -1948 17398 -1914 17416
rect -1948 17326 -1914 17348
rect -1948 17254 -1914 17280
rect -1948 17182 -1914 17212
rect -1948 17110 -1914 17144
rect -1948 17042 -1914 17076
rect -1948 16974 -1914 17004
rect -1948 16906 -1914 16932
rect -1948 16838 -1914 16860
rect -1948 16770 -1914 16788
rect -1948 16702 -1914 16716
rect -1948 16634 -1914 16644
rect -1948 16566 -1914 16572
rect -1948 16498 -1914 16500
rect -1948 16462 -1914 16464
rect -1948 16390 -1914 16396
rect -1948 16318 -1914 16328
rect -1948 16246 -1914 16260
rect -1948 16174 -1914 16192
rect -1948 16089 -1914 16124
rect -1690 18062 -1656 18097
rect -1690 17994 -1656 18012
rect -1690 17926 -1656 17940
rect -1690 17858 -1656 17868
rect -1690 17790 -1656 17796
rect -1690 17722 -1656 17724
rect -1690 17686 -1656 17688
rect -1690 17614 -1656 17620
rect -1690 17542 -1656 17552
rect -1690 17470 -1656 17484
rect -1690 17398 -1656 17416
rect -1690 17326 -1656 17348
rect -1690 17254 -1656 17280
rect -1690 17182 -1656 17212
rect -1690 17110 -1656 17144
rect -1690 17042 -1656 17076
rect -1690 16974 -1656 17004
rect -1690 16906 -1656 16932
rect -1690 16838 -1656 16860
rect -1690 16770 -1656 16788
rect -1690 16702 -1656 16716
rect -1690 16634 -1656 16644
rect -1690 16566 -1656 16572
rect -1690 16498 -1656 16500
rect -1690 16462 -1656 16464
rect -1690 16390 -1656 16396
rect -1690 16318 -1656 16328
rect -1690 16246 -1656 16260
rect -1690 16174 -1656 16192
rect -1690 16089 -1656 16124
rect -1432 18062 -1398 18097
rect -1432 17994 -1398 18012
rect -1432 17926 -1398 17940
rect -1432 17858 -1398 17868
rect -1432 17790 -1398 17796
rect -1432 17722 -1398 17724
rect -1432 17686 -1398 17688
rect -1432 17614 -1398 17620
rect -1432 17542 -1398 17552
rect -1432 17470 -1398 17484
rect -1432 17398 -1398 17416
rect -1432 17326 -1398 17348
rect -1432 17254 -1398 17280
rect -1432 17182 -1398 17212
rect -1432 17110 -1398 17144
rect -1432 17042 -1398 17076
rect -1432 16974 -1398 17004
rect -1432 16906 -1398 16932
rect -1432 16838 -1398 16860
rect -1432 16770 -1398 16788
rect -1432 16702 -1398 16716
rect -1432 16634 -1398 16644
rect -1432 16566 -1398 16572
rect -1432 16498 -1398 16500
rect -1432 16462 -1398 16464
rect -1432 16390 -1398 16396
rect -1432 16318 -1398 16328
rect -1432 16246 -1398 16260
rect -1432 16174 -1398 16192
rect -1432 16089 -1398 16124
rect -1174 18062 -1140 18097
rect -1174 17994 -1140 18012
rect -1174 17926 -1140 17940
rect -1174 17858 -1140 17868
rect -1174 17790 -1140 17796
rect -1174 17722 -1140 17724
rect -1174 17686 -1140 17688
rect -1174 17614 -1140 17620
rect -1174 17542 -1140 17552
rect -1174 17470 -1140 17484
rect -1174 17398 -1140 17416
rect -1174 17326 -1140 17348
rect -1174 17254 -1140 17280
rect -1174 17182 -1140 17212
rect -1174 17110 -1140 17144
rect -1174 17042 -1140 17076
rect -1174 16974 -1140 17004
rect -1174 16906 -1140 16932
rect -1174 16838 -1140 16860
rect -1174 16770 -1140 16788
rect -1174 16702 -1140 16716
rect -1174 16634 -1140 16644
rect -1174 16566 -1140 16572
rect -1174 16498 -1140 16500
rect -1174 16462 -1140 16464
rect -1174 16390 -1140 16396
rect -1174 16318 -1140 16328
rect -1174 16246 -1140 16260
rect -1174 16174 -1140 16192
rect -1174 16089 -1140 16124
rect -916 18062 -882 18097
rect -916 17994 -882 18012
rect -916 17926 -882 17940
rect -916 17858 -882 17868
rect -916 17790 -882 17796
rect -916 17722 -882 17724
rect -916 17686 -882 17688
rect -916 17614 -882 17620
rect -916 17542 -882 17552
rect -916 17470 -882 17484
rect -916 17398 -882 17416
rect -916 17326 -882 17348
rect -916 17254 -882 17280
rect -916 17182 -882 17212
rect -916 17110 -882 17144
rect -916 17042 -882 17076
rect -916 16974 -882 17004
rect -916 16906 -882 16932
rect -916 16838 -882 16860
rect -916 16770 -882 16788
rect -916 16702 -882 16716
rect -916 16634 -882 16644
rect -916 16566 -882 16572
rect -916 16498 -882 16500
rect -916 16462 -882 16464
rect -916 16390 -882 16396
rect -916 16318 -882 16328
rect -916 16246 -882 16260
rect -916 16174 -882 16192
rect -916 16089 -882 16124
rect -658 18062 -624 18097
rect -658 17994 -624 18012
rect -658 17926 -624 17940
rect -658 17858 -624 17868
rect -658 17790 -624 17796
rect -658 17722 -624 17724
rect -658 17686 -624 17688
rect -658 17614 -624 17620
rect -658 17542 -624 17552
rect -658 17470 -624 17484
rect -658 17398 -624 17416
rect -658 17326 -624 17348
rect -658 17254 -624 17280
rect -658 17182 -624 17212
rect -658 17110 -624 17144
rect -658 17042 -624 17076
rect -658 16974 -624 17004
rect -658 16906 -624 16932
rect -658 16838 -624 16860
rect -658 16770 -624 16788
rect -658 16702 -624 16716
rect -658 16634 -624 16644
rect -658 16566 -624 16572
rect -658 16498 -624 16500
rect -658 16462 -624 16464
rect -658 16390 -624 16396
rect -658 16318 -624 16328
rect -658 16246 -624 16260
rect -658 16174 -624 16192
rect -658 16089 -624 16124
rect -400 18062 -366 18097
rect -400 17994 -366 18012
rect -400 17926 -366 17940
rect -400 17858 -366 17868
rect -400 17790 -366 17796
rect -400 17722 -366 17724
rect -400 17686 -366 17688
rect -400 17614 -366 17620
rect -400 17542 -366 17552
rect -400 17470 -366 17484
rect -400 17398 -366 17416
rect -400 17326 -366 17348
rect -400 17254 -366 17280
rect -400 17182 -366 17212
rect -400 17110 -366 17144
rect -400 17042 -366 17076
rect -400 16974 -366 17004
rect -400 16906 -366 16932
rect -400 16838 -366 16860
rect -400 16770 -366 16788
rect -400 16702 -366 16716
rect -400 16634 -366 16644
rect -400 16566 -366 16572
rect -400 16498 -366 16500
rect -400 16462 -366 16464
rect -400 16390 -366 16396
rect -400 16318 -366 16328
rect -400 16246 -366 16260
rect -400 16174 -366 16192
rect -400 16089 -366 16124
rect -266 18062 -232 18096
rect -266 17994 -232 18028
rect -266 17926 -232 17960
rect -266 17858 -232 17892
rect -266 17790 -232 17824
rect -266 17722 -232 17756
rect -266 17654 -232 17688
rect -266 17586 -232 17620
rect -266 17518 -232 17552
rect -266 17450 -232 17484
rect -266 17382 -232 17416
rect -266 17314 -232 17348
rect -266 17246 -232 17280
rect -266 17178 -232 17212
rect -266 17110 -232 17144
rect 21862 18230 23213 18264
rect 21862 18196 23042 18230
rect 23076 18196 23176 18230
rect 21862 18194 23176 18196
rect 23210 18194 23213 18230
rect 21862 18162 23213 18194
rect 21862 18128 23042 18162
rect 23076 18128 23176 18162
rect 21862 18122 23176 18128
rect 23210 18122 23213 18162
rect 21862 18094 23213 18122
rect 21862 18060 23042 18094
rect 23076 18060 23176 18094
rect 21862 18050 23176 18060
rect 23210 18050 23213 18094
rect 21862 18032 23213 18050
rect 24234 18372 24268 18400
rect 24234 18300 24268 18332
rect 24234 18230 24268 18264
rect 24234 18162 24268 18194
rect 24234 18094 24268 18122
rect 21862 17122 22482 18032
rect 23042 18026 23076 18032
rect 23042 17958 23076 17992
rect 23042 17890 23076 17924
rect 23042 17822 23076 17856
rect 23042 17754 23076 17788
rect 23176 18026 23210 18032
rect 23176 17958 23210 17978
rect 23176 17890 23210 17906
rect 23176 17822 23210 17834
rect 23176 17743 23210 17762
rect 24234 18026 24268 18050
rect 24234 17958 24268 17978
rect 24234 17890 24268 17906
rect 24234 17822 24268 17834
rect 24234 17743 24268 17762
rect 24368 18706 24402 18740
rect 24368 18638 24402 18672
rect 24368 18570 24402 18604
rect 24558 18932 24681 18966
rect 24715 18932 24749 18966
rect 24783 18932 24817 18966
rect 24851 18932 24885 18966
rect 24919 18932 24953 18966
rect 24987 18932 25021 18966
rect 25055 18932 25089 18966
rect 25123 18932 25157 18966
rect 25191 18932 25225 18966
rect 25259 18932 25293 18966
rect 25327 18932 25361 18966
rect 25395 18932 25429 18966
rect 25463 18932 25497 18966
rect 25531 18932 25565 18966
rect 25599 18932 25633 18966
rect 25667 18932 25701 18966
rect 25735 18932 25769 18966
rect 25803 18932 25837 18966
rect 25871 18932 25905 18966
rect 25939 18932 25973 18966
rect 26007 18932 26041 18966
rect 26075 18932 26109 18966
rect 26143 18932 26177 18966
rect 26211 18932 26245 18966
rect 26279 18932 26313 18966
rect 26347 18932 26381 18966
rect 26415 18932 26449 18966
rect 26483 18932 26517 18966
rect 26551 18932 26585 18966
rect 26619 18932 26653 18966
rect 26687 18932 26721 18966
rect 26755 18932 26789 18966
rect 26823 18932 26857 18966
rect 26891 18932 26925 18966
rect 26959 18932 26993 18966
rect 27027 18932 27061 18966
rect 27095 18932 27129 18966
rect 27163 18932 27197 18966
rect 27231 18932 27265 18966
rect 27299 18932 27333 18966
rect 27367 18932 27401 18966
rect 27435 18932 27469 18966
rect 27503 18932 27537 18966
rect 27571 18932 27605 18966
rect 27639 18932 27673 18966
rect 27707 18932 27741 18966
rect 27775 18932 27809 18966
rect 27843 18932 27877 18966
rect 27911 18932 28034 18966
rect 24558 18848 24592 18932
rect 28000 18848 28034 18932
rect 24558 18780 24592 18814
rect 24738 18794 24779 18828
rect 24823 18794 24847 18828
rect 24895 18794 24915 18828
rect 24967 18794 24983 18828
rect 25039 18794 25051 18828
rect 25111 18794 25119 18828
rect 25183 18794 25187 18828
rect 25289 18794 25293 18828
rect 25357 18794 25365 18828
rect 25425 18794 25437 18828
rect 25493 18794 25509 18828
rect 25561 18794 25581 18828
rect 25629 18794 25653 18828
rect 25697 18794 25738 18828
rect 25796 18794 25837 18828
rect 25881 18794 25905 18828
rect 25953 18794 25973 18828
rect 26025 18794 26041 18828
rect 26097 18794 26109 18828
rect 26169 18794 26177 18828
rect 26241 18794 26245 18828
rect 26347 18794 26351 18828
rect 26415 18794 26423 18828
rect 26483 18794 26495 18828
rect 26551 18794 26567 18828
rect 26619 18794 26639 18828
rect 26687 18794 26711 18828
rect 26755 18794 26796 18828
rect 26854 18794 26895 18828
rect 26939 18794 26963 18828
rect 27011 18794 27031 18828
rect 27083 18794 27099 18828
rect 27155 18794 27167 18828
rect 27227 18794 27235 18828
rect 27299 18794 27303 18828
rect 27405 18794 27409 18828
rect 27473 18794 27481 18828
rect 27541 18794 27553 18828
rect 27609 18794 27625 18828
rect 27677 18794 27697 18828
rect 27745 18794 27769 18828
rect 27813 18794 27854 18828
rect 28000 18780 28034 18814
rect 24558 18712 24592 18746
rect 24558 18644 24592 18678
rect 24558 18576 24592 18610
rect 24368 18502 24402 18536
rect 24368 18434 24402 18468
rect 24368 18366 24402 18400
rect 24546 18542 24558 18544
rect 24692 18720 24726 18751
rect 24692 18648 24726 18678
rect 24692 18576 24726 18610
rect 24592 18542 24692 18544
rect 25750 18720 25784 18751
rect 25750 18648 25784 18678
rect 25750 18576 25784 18610
rect 24726 18542 24738 18544
rect 24546 18508 24738 18542
rect 24546 18474 24558 18508
rect 24592 18474 24692 18508
rect 24546 18470 24692 18474
rect 24726 18470 24738 18508
rect 24546 18440 24738 18470
rect 24546 18406 24558 18440
rect 24592 18406 24692 18440
rect 24546 18398 24692 18406
rect 24726 18398 24738 18440
rect 24546 18372 24738 18398
rect 24546 18362 24558 18372
rect 24368 18298 24402 18332
rect 24368 18230 24402 18264
rect 24368 18162 24402 18196
rect 24368 18094 24402 18128
rect 24368 18026 24402 18060
rect 24368 17958 24402 17992
rect 24368 17890 24402 17924
rect 24368 17822 24402 17856
rect 24368 17754 24402 17788
rect 23042 17686 23076 17720
rect 23222 17666 23263 17700
rect 23307 17666 23331 17700
rect 23379 17666 23399 17700
rect 23451 17666 23467 17700
rect 23523 17666 23535 17700
rect 23595 17666 23603 17700
rect 23667 17666 23671 17700
rect 23773 17666 23777 17700
rect 23841 17666 23849 17700
rect 23909 17666 23921 17700
rect 23977 17666 23993 17700
rect 24045 17666 24065 17700
rect 24113 17666 24137 17700
rect 24181 17666 24222 17700
rect 24368 17686 24402 17720
rect 23042 17562 23076 17652
rect 24368 17562 24402 17652
rect 23042 17528 23161 17562
rect 23195 17528 23229 17562
rect 23263 17528 23297 17562
rect 23331 17528 23365 17562
rect 23399 17528 23433 17562
rect 23467 17528 23501 17562
rect 23535 17528 23569 17562
rect 23603 17528 23637 17562
rect 23671 17528 23705 17562
rect 23739 17528 23773 17562
rect 23807 17528 23841 17562
rect 23875 17528 23909 17562
rect 23943 17528 23977 17562
rect 24011 17528 24045 17562
rect 24079 17528 24113 17562
rect 24147 17528 24181 17562
rect 24215 17528 24249 17562
rect 24283 17528 24402 17562
rect 24592 18362 24692 18372
rect 24558 18304 24592 18338
rect 24558 18236 24592 18270
rect 24558 18168 24592 18202
rect 24558 18100 24592 18134
rect 24558 18032 24592 18066
rect 24558 17964 24592 17998
rect 24558 17896 24592 17930
rect 24558 17828 24592 17862
rect 24558 17760 24592 17794
rect 24558 17692 24592 17726
rect 24558 17624 24592 17658
rect 24558 17556 24592 17590
rect 24558 17488 24592 17522
rect 24558 17420 24592 17454
rect 24558 17352 24592 17386
rect -266 17042 -232 17076
rect -266 16974 -232 17008
rect -266 16906 -232 16940
rect -266 16838 -232 16872
rect -266 16770 -232 16804
rect -266 16702 -232 16736
rect -266 16634 -232 16668
rect -266 16566 -232 16600
rect -266 16498 -232 16532
rect -266 16430 -232 16464
rect -266 16362 -232 16396
rect -266 16294 -232 16328
rect -266 16226 -232 16260
rect -266 16158 -232 16192
rect -266 16090 -232 16124
rect -3114 16022 -3080 16056
rect -2934 16012 -2887 16046
rect -2851 16012 -2817 16046
rect -2781 16012 -2734 16046
rect -2676 16012 -2629 16046
rect -2593 16012 -2559 16046
rect -2523 16012 -2476 16046
rect -2418 16012 -2371 16046
rect -2335 16012 -2301 16046
rect -2265 16012 -2218 16046
rect -2160 16012 -2113 16046
rect -2077 16012 -2043 16046
rect -2007 16012 -1960 16046
rect -1902 16012 -1855 16046
rect -1819 16012 -1785 16046
rect -1749 16012 -1702 16046
rect -1644 16012 -1597 16046
rect -1561 16012 -1527 16046
rect -1491 16012 -1444 16046
rect -1386 16012 -1339 16046
rect -1303 16012 -1269 16046
rect -1233 16012 -1186 16046
rect -1128 16012 -1081 16046
rect -1045 16012 -1011 16046
rect -975 16012 -928 16046
rect -870 16012 -823 16046
rect -787 16012 -753 16046
rect -717 16012 -670 16046
rect -612 16012 -565 16046
rect -529 16012 -495 16046
rect -459 16012 -412 16046
rect -266 16022 -232 16056
rect -3114 15908 -3080 15988
rect -266 15908 -232 15988
rect -3114 15874 -3016 15908
rect -2982 15874 -2948 15908
rect -2914 15874 -2880 15908
rect -2846 15874 -2812 15908
rect -2778 15874 -2744 15908
rect -2710 15874 -2676 15908
rect -2642 15874 -2608 15908
rect -2574 15874 -2540 15908
rect -2506 15874 -2472 15908
rect -2438 15874 -2404 15908
rect -2370 15874 -2336 15908
rect -2302 15874 -2268 15908
rect -2234 15874 -2200 15908
rect -2166 15874 -2132 15908
rect -2098 15874 -2064 15908
rect -2030 15874 -1996 15908
rect -1962 15874 -1928 15908
rect -1894 15874 -1860 15908
rect -1826 15874 -1792 15908
rect -1758 15874 -1724 15908
rect -1690 15874 -1656 15908
rect -1622 15874 -1588 15908
rect -1554 15874 -1520 15908
rect -1486 15874 -1452 15908
rect -1418 15874 -1384 15908
rect -1350 15874 -1316 15908
rect -1282 15874 -1248 15908
rect -1214 15874 -1180 15908
rect -1146 15874 -1112 15908
rect -1078 15874 -1044 15908
rect -1010 15874 -976 15908
rect -942 15874 -908 15908
rect -874 15874 -840 15908
rect -806 15874 -772 15908
rect -738 15874 -704 15908
rect -670 15874 -636 15908
rect -602 15874 -568 15908
rect -534 15874 -500 15908
rect -466 15874 -432 15908
rect -398 15874 -364 15908
rect -330 15874 -232 15908
rect 10297 17061 22482 17122
rect -7886 15466 -4427 15515
rect -7886 15432 -7630 15466
rect -7596 15432 -7562 15466
rect -7528 15432 -7494 15466
rect -7460 15432 -7426 15466
rect -7392 15432 -7358 15466
rect -7324 15432 -7290 15466
rect -7256 15432 -7222 15466
rect -7188 15432 -7154 15466
rect -7120 15432 -7086 15466
rect -7052 15432 -7018 15466
rect -6984 15432 -6950 15466
rect -6916 15432 -6882 15466
rect -6848 15432 -6814 15466
rect -6780 15432 -6746 15466
rect -6712 15432 -6678 15466
rect -6644 15432 -6610 15466
rect -6576 15432 -6542 15466
rect -6508 15432 -6474 15466
rect -6440 15432 -6406 15466
rect -6372 15432 -6338 15466
rect -6304 15432 -6270 15466
rect -6236 15432 -6202 15466
rect -6168 15432 -6134 15466
rect -6100 15432 -6066 15466
rect -6032 15432 -5998 15466
rect -5964 15432 -5930 15466
rect -5896 15432 -5862 15466
rect -5828 15432 -5794 15466
rect -5760 15432 -5726 15466
rect -5692 15432 -5658 15466
rect -5624 15432 -5590 15466
rect -5556 15432 -5522 15466
rect -5488 15432 -5454 15466
rect -5420 15432 -5386 15466
rect -5352 15432 -5318 15466
rect -5284 15432 -5250 15466
rect -5216 15432 -5182 15466
rect -5148 15432 -5114 15466
rect -5080 15432 -5046 15466
rect -5012 15432 -4978 15466
rect -4944 15432 -4910 15466
rect -4876 15432 -4842 15466
rect -4808 15432 -4774 15466
rect -4740 15432 -4706 15466
rect -4672 15432 -4427 15466
rect -7886 15381 -4427 15432
rect -7886 15308 -7753 15381
rect -7886 15274 -7843 15308
rect -7809 15274 -7753 15308
rect -7886 15240 -7753 15274
rect -7886 15206 -7843 15240
rect -7809 15206 -7753 15240
rect -4545 15268 -4427 15381
rect -4545 15234 -4503 15268
rect -4469 15234 -4427 15268
rect -7886 15172 -7753 15206
rect -7886 15138 -7843 15172
rect -7809 15138 -7753 15172
rect -7886 15104 -7753 15138
rect -7886 15070 -7843 15104
rect -7809 15070 -7753 15104
rect -7886 15036 -7753 15070
rect -7886 15002 -7843 15036
rect -7809 15002 -7753 15036
rect -7886 14968 -7753 15002
rect -7886 14934 -7843 14968
rect -7809 14934 -7753 14968
rect -7886 14900 -7753 14934
rect -7138 15163 -6726 15212
rect -7138 15057 -7075 15163
rect -6825 15057 -6726 15163
rect -7138 14968 -6726 15057
rect -7138 14934 -7080 14968
rect -7046 14934 -6820 14968
rect -6786 14934 -6726 14968
rect -6095 15162 -5697 15213
rect -6095 15056 -6059 15162
rect -5737 15056 -5697 15162
rect -6095 14981 -5697 15056
rect -5061 15171 -4913 15212
rect -5061 15137 -5006 15171
rect -4972 15137 -4913 15171
rect -5061 15099 -4913 15137
rect -5061 15065 -5006 15099
rect -4972 15065 -4913 15099
rect -6095 14957 -5696 14981
rect -7138 14902 -6726 14934
rect -6689 14912 -6129 14956
rect -7886 14866 -7843 14900
rect -7809 14866 -7753 14900
rect -7886 14832 -7753 14866
rect -7886 14798 -7843 14832
rect -7809 14798 -7753 14832
rect -7886 14764 -7753 14798
rect -7886 14730 -7843 14764
rect -7809 14730 -7753 14764
rect -7886 14696 -7753 14730
rect -7886 14662 -7843 14696
rect -7809 14662 -7753 14696
rect -7886 14628 -7753 14662
rect -7886 14594 -7843 14628
rect -7809 14594 -7753 14628
rect -7886 14560 -7753 14594
rect -7886 14526 -7843 14560
rect -7809 14526 -7753 14560
rect -7886 14492 -7753 14526
rect -7886 14458 -7843 14492
rect -7809 14458 -7753 14492
rect -7886 14424 -7753 14458
rect -7886 14390 -7843 14424
rect -7809 14390 -7753 14424
rect -7886 14356 -7753 14390
rect -7886 14322 -7843 14356
rect -7809 14322 -7753 14356
rect -7886 14288 -7753 14322
rect -7886 14254 -7843 14288
rect -7809 14254 -7753 14288
rect -7886 14220 -7753 14254
rect -7886 14186 -7843 14220
rect -7809 14186 -7753 14220
rect -7886 14152 -7753 14186
rect -7886 14118 -7843 14152
rect -7809 14118 -7753 14152
rect -7886 14084 -7753 14118
rect -7886 14050 -7843 14084
rect -7809 14050 -7753 14084
rect -7886 14016 -7753 14050
rect -7886 13982 -7843 14016
rect -7809 13982 -7753 14016
rect -7886 13948 -7753 13982
rect -7886 13914 -7843 13948
rect -7809 13914 -7753 13948
rect -7886 13880 -7753 13914
rect -7886 13846 -7843 13880
rect -7809 13846 -7753 13880
rect -7886 13812 -7753 13846
rect -7886 13778 -7843 13812
rect -7809 13778 -7753 13812
rect -7886 13744 -7753 13778
rect -7886 13710 -7843 13744
rect -7809 13710 -7753 13744
rect -7886 13676 -7753 13710
rect -7886 13642 -7843 13676
rect -7809 13642 -7753 13676
rect -7886 13608 -7753 13642
rect -7886 13574 -7843 13608
rect -7809 13574 -7753 13608
rect -7886 13540 -7753 13574
rect -7886 13506 -7843 13540
rect -7809 13506 -7753 13540
rect -7886 13472 -7753 13506
rect -7886 13438 -7843 13472
rect -7809 13438 -7753 13472
rect -7886 13404 -7753 13438
rect -7886 13370 -7843 13404
rect -7809 13370 -7753 13404
rect -7886 13336 -7753 13370
rect -7886 13302 -7843 13336
rect -7809 13302 -7753 13336
rect -7886 13268 -7753 13302
rect -7886 13234 -7843 13268
rect -7809 13234 -7753 13268
rect -7886 13200 -7753 13234
rect -7886 13166 -7843 13200
rect -7809 13166 -7753 13200
rect -7886 13132 -7753 13166
rect -7886 13098 -7843 13132
rect -7809 13098 -7753 13132
rect -7886 13064 -7753 13098
rect -7886 13030 -7843 13064
rect -7809 13030 -7753 13064
rect -7886 12996 -7753 13030
rect -7886 12962 -7843 12996
rect -7809 12962 -7753 12996
rect -7886 12928 -7753 12962
rect -7886 12894 -7843 12928
rect -7809 12894 -7753 12928
rect -7886 12860 -7753 12894
rect -7886 12826 -7843 12860
rect -7809 12826 -7753 12860
rect -7459 14804 -7425 14839
rect -7459 14736 -7425 14754
rect -7459 14668 -7425 14682
rect -7459 14600 -7425 14610
rect -7459 14532 -7425 14538
rect -7459 14464 -7425 14466
rect -7459 14428 -7425 14430
rect -7459 14356 -7425 14362
rect -7459 14284 -7425 14294
rect -7459 14212 -7425 14226
rect -7459 14140 -7425 14158
rect -7459 14068 -7425 14090
rect -7459 13996 -7425 14022
rect -7459 13924 -7425 13954
rect -7459 13852 -7425 13886
rect -7459 13784 -7425 13818
rect -7459 13716 -7425 13746
rect -7459 13648 -7425 13674
rect -7459 13580 -7425 13602
rect -7459 13512 -7425 13530
rect -7459 13444 -7425 13458
rect -7459 13376 -7425 13386
rect -7459 13308 -7425 13314
rect -7459 13240 -7425 13242
rect -7459 13204 -7425 13206
rect -7459 13132 -7425 13138
rect -7459 13060 -7425 13070
rect -7459 12988 -7425 13002
rect -7459 12916 -7425 12934
rect -7201 14804 -7167 14839
rect -7201 14736 -7167 14754
rect -7201 14668 -7167 14682
rect -7201 14600 -7167 14610
rect -7201 14532 -7167 14538
rect -7201 14464 -7167 14466
rect -7201 14428 -7167 14430
rect -7201 14356 -7167 14362
rect -7201 14284 -7167 14294
rect -7201 14212 -7167 14226
rect -7201 14140 -7167 14158
rect -7201 14068 -7167 14090
rect -7201 13996 -7167 14022
rect -7201 13924 -7167 13954
rect -7201 13852 -7167 13886
rect -7201 13784 -7167 13818
rect -7201 13716 -7167 13746
rect -7201 13648 -7167 13674
rect -7201 13580 -7167 13602
rect -7201 13512 -7167 13530
rect -7201 13444 -7167 13458
rect -7201 13376 -7167 13386
rect -7201 13308 -7167 13314
rect -7201 13240 -7167 13242
rect -7201 13204 -7167 13206
rect -7201 13132 -7167 13138
rect -7201 13060 -7167 13070
rect -7201 12988 -7167 13002
rect -7201 12916 -7167 12934
rect -7459 12831 -7425 12866
rect -7207 12866 -7201 12871
rect -6943 14804 -6909 14839
rect -6943 14736 -6909 14754
rect -6943 14668 -6909 14682
rect -6943 14600 -6909 14610
rect -6943 14532 -6909 14538
rect -6943 14464 -6909 14466
rect -6943 14428 -6909 14430
rect -6943 14356 -6909 14362
rect -6943 14284 -6909 14294
rect -6943 14212 -6909 14226
rect -6943 14140 -6909 14158
rect -6943 14068 -6909 14090
rect -6943 13996 -6909 14022
rect -6943 13924 -6909 13954
rect -6943 13852 -6909 13886
rect -6943 13784 -6909 13818
rect -6943 13716 -6909 13746
rect -6943 13648 -6909 13674
rect -6943 13580 -6909 13602
rect -6943 13512 -6909 13530
rect -6943 13444 -6909 13458
rect -6943 13376 -6909 13386
rect -6943 13308 -6909 13314
rect -6943 13240 -6909 13242
rect -6943 13204 -6909 13206
rect -6943 13132 -6909 13138
rect -6943 13060 -6909 13070
rect -6943 12988 -6909 13002
rect -6943 12916 -6909 12934
rect -7167 12866 -7163 12871
rect -7886 12792 -7753 12826
rect -7886 12758 -7843 12792
rect -7809 12758 -7753 12792
rect -7886 12724 -7753 12758
rect -7207 12763 -7163 12866
rect -6943 12831 -6909 12866
rect -6689 14804 -6645 14912
rect -6689 14754 -6685 14804
rect -6651 14754 -6645 14804
rect -6689 14736 -6645 14754
rect -6689 14682 -6685 14736
rect -6651 14682 -6645 14736
rect -6689 14668 -6645 14682
rect -6689 14610 -6685 14668
rect -6651 14610 -6645 14668
rect -6689 14600 -6645 14610
rect -6689 14538 -6685 14600
rect -6651 14538 -6645 14600
rect -6689 14532 -6645 14538
rect -6689 14466 -6685 14532
rect -6651 14466 -6645 14532
rect -6689 14464 -6645 14466
rect -6689 14430 -6685 14464
rect -6651 14430 -6645 14464
rect -6689 14428 -6645 14430
rect -6689 14362 -6685 14428
rect -6651 14362 -6645 14428
rect -6689 14356 -6645 14362
rect -6689 14294 -6685 14356
rect -6651 14294 -6645 14356
rect -6689 14284 -6645 14294
rect -6689 14226 -6685 14284
rect -6651 14226 -6645 14284
rect -6689 14212 -6645 14226
rect -6689 14158 -6685 14212
rect -6651 14158 -6645 14212
rect -6689 14140 -6645 14158
rect -6689 14090 -6685 14140
rect -6651 14090 -6645 14140
rect -6689 14068 -6645 14090
rect -6689 14022 -6685 14068
rect -6651 14022 -6645 14068
rect -6689 13996 -6645 14022
rect -6689 13954 -6685 13996
rect -6651 13954 -6645 13996
rect -6689 13924 -6645 13954
rect -6689 13886 -6685 13924
rect -6651 13886 -6645 13924
rect -6689 13852 -6645 13886
rect -6689 13818 -6685 13852
rect -6651 13818 -6645 13852
rect -6689 13784 -6645 13818
rect -6689 13746 -6685 13784
rect -6651 13746 -6645 13784
rect -6689 13716 -6645 13746
rect -6689 13674 -6685 13716
rect -6651 13674 -6645 13716
rect -6689 13648 -6645 13674
rect -6689 13602 -6685 13648
rect -6651 13602 -6645 13648
rect -6689 13580 -6645 13602
rect -6689 13530 -6685 13580
rect -6651 13530 -6645 13580
rect -6689 13512 -6645 13530
rect -6689 13458 -6685 13512
rect -6651 13458 -6645 13512
rect -6689 13444 -6645 13458
rect -6689 13386 -6685 13444
rect -6651 13386 -6645 13444
rect -6689 13376 -6645 13386
rect -6689 13314 -6685 13376
rect -6651 13314 -6645 13376
rect -6689 13308 -6645 13314
rect -6689 13242 -6685 13308
rect -6651 13242 -6645 13308
rect -6689 13240 -6645 13242
rect -6689 13206 -6685 13240
rect -6651 13206 -6645 13240
rect -6689 13204 -6645 13206
rect -6689 13138 -6685 13204
rect -6651 13138 -6645 13204
rect -6689 13132 -6645 13138
rect -6689 13070 -6685 13132
rect -6651 13070 -6645 13132
rect -6689 13060 -6645 13070
rect -6689 13002 -6685 13060
rect -6651 13002 -6645 13060
rect -6689 12988 -6645 13002
rect -6689 12934 -6685 12988
rect -6651 12934 -6645 12988
rect -6689 12916 -6645 12934
rect -6689 12866 -6685 12916
rect -6651 12866 -6645 12916
rect -6689 12783 -6645 12866
rect -6427 14804 -6393 14839
rect -6427 14736 -6393 14754
rect -6427 14668 -6393 14682
rect -6427 14600 -6393 14610
rect -6427 14532 -6393 14538
rect -6427 14464 -6393 14466
rect -6427 14428 -6393 14430
rect -6427 14356 -6393 14362
rect -6427 14284 -6393 14294
rect -6427 14212 -6393 14226
rect -6427 14140 -6393 14158
rect -6427 14068 -6393 14090
rect -6427 13996 -6393 14022
rect -6427 13924 -6393 13954
rect -6427 13852 -6393 13886
rect -6427 13784 -6393 13818
rect -6427 13716 -6393 13746
rect -6427 13648 -6393 13674
rect -6427 13580 -6393 13602
rect -6427 13512 -6393 13530
rect -6427 13444 -6393 13458
rect -6427 13376 -6393 13386
rect -6427 13308 -6393 13314
rect -6427 13240 -6393 13242
rect -6427 13204 -6393 13206
rect -6427 13132 -6393 13138
rect -6427 13060 -6393 13070
rect -6427 12988 -6393 13002
rect -6427 12916 -6393 12934
rect -6427 12831 -6393 12866
rect -6173 14804 -6129 14912
rect -6095 14923 -6028 14957
rect -5994 14944 -5696 14957
rect -5466 14954 -5226 14964
rect -5994 14923 -5778 14944
rect -6095 14910 -5778 14923
rect -5744 14910 -5696 14944
rect -6095 14874 -5696 14910
rect -5660 14935 -5101 14954
rect -5660 14910 -5436 14935
rect -6173 14754 -6169 14804
rect -6135 14754 -6129 14804
rect -6173 14736 -6129 14754
rect -6173 14682 -6169 14736
rect -6135 14682 -6129 14736
rect -6173 14668 -6129 14682
rect -6173 14610 -6169 14668
rect -6135 14610 -6129 14668
rect -6173 14600 -6129 14610
rect -6173 14538 -6169 14600
rect -6135 14538 -6129 14600
rect -6173 14532 -6129 14538
rect -6173 14466 -6169 14532
rect -6135 14466 -6129 14532
rect -6173 14464 -6129 14466
rect -6173 14430 -6169 14464
rect -6135 14430 -6129 14464
rect -6173 14428 -6129 14430
rect -6173 14362 -6169 14428
rect -6135 14362 -6129 14428
rect -6173 14356 -6129 14362
rect -6173 14294 -6169 14356
rect -6135 14294 -6129 14356
rect -6173 14284 -6129 14294
rect -6173 14226 -6169 14284
rect -6135 14226 -6129 14284
rect -6173 14212 -6129 14226
rect -6173 14158 -6169 14212
rect -6135 14158 -6129 14212
rect -6173 14140 -6129 14158
rect -6173 14090 -6169 14140
rect -6135 14090 -6129 14140
rect -6173 14068 -6129 14090
rect -6173 14022 -6169 14068
rect -6135 14022 -6129 14068
rect -6173 13996 -6129 14022
rect -6173 13954 -6169 13996
rect -6135 13954 -6129 13996
rect -6173 13924 -6129 13954
rect -6173 13886 -6169 13924
rect -6135 13886 -6129 13924
rect -6173 13852 -6129 13886
rect -6173 13818 -6169 13852
rect -6135 13818 -6129 13852
rect -6173 13784 -6129 13818
rect -6173 13746 -6169 13784
rect -6135 13746 -6129 13784
rect -6173 13716 -6129 13746
rect -6173 13674 -6169 13716
rect -6135 13674 -6129 13716
rect -6173 13648 -6129 13674
rect -6173 13602 -6169 13648
rect -6135 13602 -6129 13648
rect -6173 13580 -6129 13602
rect -6173 13530 -6169 13580
rect -6135 13530 -6129 13580
rect -6173 13512 -6129 13530
rect -6173 13458 -6169 13512
rect -6135 13458 -6129 13512
rect -6173 13444 -6129 13458
rect -6173 13386 -6169 13444
rect -6135 13386 -6129 13444
rect -6173 13376 -6129 13386
rect -6173 13314 -6169 13376
rect -6135 13314 -6129 13376
rect -6173 13308 -6129 13314
rect -6173 13242 -6169 13308
rect -6135 13242 -6129 13308
rect -6173 13240 -6129 13242
rect -6173 13206 -6169 13240
rect -6135 13206 -6129 13240
rect -6173 13204 -6129 13206
rect -6173 13138 -6169 13204
rect -6135 13138 -6129 13204
rect -6173 13132 -6129 13138
rect -6173 13070 -6169 13132
rect -6135 13070 -6129 13132
rect -6173 13060 -6129 13070
rect -6173 13002 -6169 13060
rect -6135 13002 -6129 13060
rect -6173 12988 -6129 13002
rect -6173 12934 -6169 12988
rect -6135 12934 -6129 12988
rect -6173 12916 -6129 12934
rect -6173 12866 -6169 12916
rect -6135 12866 -6129 12916
rect -6874 12763 -6645 12783
rect -7207 12758 -6645 12763
rect -7886 12690 -7843 12724
rect -7809 12690 -7753 12724
rect -7886 12656 -7753 12690
rect -7886 12622 -7843 12656
rect -7809 12622 -7753 12656
rect -7392 12721 -7246 12754
rect -7392 12687 -7343 12721
rect -7309 12687 -7246 12721
rect -7207 12724 -6840 12758
rect -6806 12724 -6768 12758
rect -6734 12724 -6645 12758
rect -6173 12762 -6129 12866
rect -5911 14804 -5877 14839
rect -5911 14736 -5877 14754
rect -5911 14668 -5877 14682
rect -5911 14600 -5877 14610
rect -5911 14532 -5877 14538
rect -5911 14464 -5877 14466
rect -5911 14428 -5877 14430
rect -5911 14356 -5877 14362
rect -5911 14284 -5877 14294
rect -5911 14212 -5877 14226
rect -5911 14140 -5877 14158
rect -5911 14068 -5877 14090
rect -5911 13996 -5877 14022
rect -5911 13924 -5877 13954
rect -5911 13852 -5877 13886
rect -5911 13784 -5877 13818
rect -5911 13716 -5877 13746
rect -5911 13648 -5877 13674
rect -5911 13580 -5877 13602
rect -5911 13512 -5877 13530
rect -5911 13444 -5877 13458
rect -5911 13376 -5877 13386
rect -5911 13308 -5877 13314
rect -5911 13240 -5877 13242
rect -5911 13204 -5877 13206
rect -5911 13132 -5877 13138
rect -5911 13060 -5877 13070
rect -5911 12988 -5877 13002
rect -5911 12916 -5877 12934
rect -5911 12831 -5877 12866
rect -5660 14804 -5616 14910
rect -5466 14901 -5436 14910
rect -5402 14901 -5364 14935
rect -5330 14901 -5292 14935
rect -5258 14910 -5101 14935
rect -5258 14901 -5226 14910
rect -5466 14874 -5226 14901
rect -5660 14754 -5653 14804
rect -5619 14754 -5616 14804
rect -5660 14736 -5616 14754
rect -5660 14682 -5653 14736
rect -5619 14682 -5616 14736
rect -5660 14668 -5616 14682
rect -5660 14610 -5653 14668
rect -5619 14610 -5616 14668
rect -5660 14600 -5616 14610
rect -5660 14538 -5653 14600
rect -5619 14538 -5616 14600
rect -5660 14532 -5616 14538
rect -5660 14466 -5653 14532
rect -5619 14466 -5616 14532
rect -5660 14464 -5616 14466
rect -5660 14430 -5653 14464
rect -5619 14430 -5616 14464
rect -5660 14428 -5616 14430
rect -5660 14362 -5653 14428
rect -5619 14362 -5616 14428
rect -5660 14356 -5616 14362
rect -5660 14294 -5653 14356
rect -5619 14294 -5616 14356
rect -5660 14284 -5616 14294
rect -5660 14226 -5653 14284
rect -5619 14226 -5616 14284
rect -5660 14212 -5616 14226
rect -5660 14158 -5653 14212
rect -5619 14158 -5616 14212
rect -5660 14140 -5616 14158
rect -5660 14090 -5653 14140
rect -5619 14090 -5616 14140
rect -5660 14068 -5616 14090
rect -5660 14022 -5653 14068
rect -5619 14022 -5616 14068
rect -5660 13996 -5616 14022
rect -5660 13954 -5653 13996
rect -5619 13954 -5616 13996
rect -5660 13924 -5616 13954
rect -5660 13886 -5653 13924
rect -5619 13886 -5616 13924
rect -5660 13852 -5616 13886
rect -5660 13818 -5653 13852
rect -5619 13818 -5616 13852
rect -5660 13784 -5616 13818
rect -5660 13746 -5653 13784
rect -5619 13746 -5616 13784
rect -5660 13716 -5616 13746
rect -5660 13674 -5653 13716
rect -5619 13674 -5616 13716
rect -5660 13648 -5616 13674
rect -5660 13602 -5653 13648
rect -5619 13602 -5616 13648
rect -5660 13580 -5616 13602
rect -5660 13530 -5653 13580
rect -5619 13530 -5616 13580
rect -5660 13512 -5616 13530
rect -5660 13458 -5653 13512
rect -5619 13458 -5616 13512
rect -5660 13444 -5616 13458
rect -5660 13386 -5653 13444
rect -5619 13386 -5616 13444
rect -5660 13376 -5616 13386
rect -5660 13314 -5653 13376
rect -5619 13314 -5616 13376
rect -5660 13308 -5616 13314
rect -5660 13242 -5653 13308
rect -5619 13242 -5616 13308
rect -5660 13240 -5616 13242
rect -5660 13206 -5653 13240
rect -5619 13206 -5616 13240
rect -5660 13204 -5616 13206
rect -5660 13138 -5653 13204
rect -5619 13138 -5616 13204
rect -5660 13132 -5616 13138
rect -5660 13070 -5653 13132
rect -5619 13070 -5616 13132
rect -5660 13060 -5616 13070
rect -5660 13002 -5653 13060
rect -5619 13002 -5616 13060
rect -5660 12988 -5616 13002
rect -5660 12934 -5653 12988
rect -5619 12934 -5616 12988
rect -5660 12916 -5616 12934
rect -5660 12866 -5653 12916
rect -5619 12866 -5616 12916
rect -5660 12762 -5616 12866
rect -5395 14804 -5361 14839
rect -5145 14804 -5101 14910
rect -5061 14948 -4913 15065
rect -5061 14914 -5007 14948
rect -4973 14914 -4913 14948
rect -5061 14909 -4913 14914
rect -4545 15200 -4427 15234
rect -4545 15166 -4503 15200
rect -4469 15166 -4427 15200
rect -4545 15132 -4427 15166
rect -4545 15098 -4503 15132
rect -4469 15098 -4427 15132
rect -4545 15064 -4427 15098
rect -4545 15030 -4503 15064
rect -4469 15030 -4427 15064
rect -4545 14996 -4427 15030
rect -4545 14962 -4503 14996
rect -4469 14962 -4427 14996
rect -4545 14928 -4427 14962
rect -5061 14874 -4921 14909
rect -4545 14894 -4503 14928
rect -4469 14894 -4427 14928
rect -4545 14860 -4427 14894
rect -5145 14777 -5137 14804
rect -5395 14736 -5361 14754
rect -5395 14668 -5361 14682
rect -5395 14600 -5361 14610
rect -5395 14532 -5361 14538
rect -5395 14464 -5361 14466
rect -5395 14428 -5361 14430
rect -5395 14356 -5361 14362
rect -5395 14284 -5361 14294
rect -5395 14212 -5361 14226
rect -5395 14140 -5361 14158
rect -5395 14068 -5361 14090
rect -5395 13996 -5361 14022
rect -5395 13924 -5361 13954
rect -5395 13852 -5361 13886
rect -5395 13784 -5361 13818
rect -5395 13716 -5361 13746
rect -5395 13648 -5361 13674
rect -5395 13580 -5361 13602
rect -5395 13512 -5361 13530
rect -5395 13444 -5361 13458
rect -5395 13376 -5361 13386
rect -5395 13308 -5361 13314
rect -5395 13240 -5361 13242
rect -5395 13204 -5361 13206
rect -5395 13132 -5361 13138
rect -5395 13060 -5361 13070
rect -5395 12988 -5361 13002
rect -5395 12916 -5361 12934
rect -5395 12831 -5361 12866
rect -5103 14777 -5101 14804
rect -4879 14804 -4845 14839
rect -5137 14736 -5103 14754
rect -5137 14668 -5103 14682
rect -5137 14600 -5103 14610
rect -5137 14532 -5103 14538
rect -5137 14464 -5103 14466
rect -5137 14428 -5103 14430
rect -5137 14356 -5103 14362
rect -5137 14284 -5103 14294
rect -5137 14212 -5103 14226
rect -5137 14140 -5103 14158
rect -5137 14068 -5103 14090
rect -5137 13996 -5103 14022
rect -5137 13924 -5103 13954
rect -5137 13852 -5103 13886
rect -5137 13784 -5103 13818
rect -5137 13716 -5103 13746
rect -5137 13648 -5103 13674
rect -5137 13580 -5103 13602
rect -5137 13512 -5103 13530
rect -5137 13444 -5103 13458
rect -5137 13376 -5103 13386
rect -5137 13308 -5103 13314
rect -5137 13240 -5103 13242
rect -5137 13204 -5103 13206
rect -5137 13132 -5103 13138
rect -5137 13060 -5103 13070
rect -5137 12988 -5103 13002
rect -5137 12916 -5103 12934
rect -5137 12831 -5103 12866
rect -4879 14736 -4845 14754
rect -4879 14668 -4845 14682
rect -4879 14600 -4845 14610
rect -4879 14532 -4845 14538
rect -4879 14464 -4845 14466
rect -4879 14428 -4845 14430
rect -4879 14356 -4845 14362
rect -4879 14284 -4845 14294
rect -4879 14212 -4845 14226
rect -4879 14140 -4845 14158
rect -4879 14068 -4845 14090
rect -4879 13996 -4845 14022
rect -4879 13924 -4845 13954
rect -4879 13852 -4845 13886
rect -4879 13784 -4845 13818
rect -4879 13716 -4845 13746
rect -4879 13648 -4845 13674
rect -4879 13580 -4845 13602
rect -4879 13512 -4845 13530
rect -4879 13444 -4845 13458
rect -4879 13376 -4845 13386
rect -4879 13308 -4845 13314
rect -4879 13240 -4845 13242
rect -4879 13204 -4845 13206
rect -4879 13132 -4845 13138
rect -4879 13060 -4845 13070
rect -4879 12988 -4845 13002
rect -4879 12916 -4845 12934
rect -4879 12831 -4845 12866
rect -4545 14826 -4503 14860
rect -4469 14826 -4427 14860
rect -4545 14792 -4427 14826
rect -4545 14758 -4503 14792
rect -4469 14758 -4427 14792
rect -4545 14724 -4427 14758
rect -4545 14690 -4503 14724
rect -4469 14690 -4427 14724
rect -4545 14656 -4427 14690
rect -4545 14622 -4503 14656
rect -4469 14622 -4427 14656
rect -4545 14588 -4427 14622
rect -4545 14554 -4503 14588
rect -4469 14554 -4427 14588
rect -4545 14520 -4427 14554
rect -4545 14486 -4503 14520
rect -4469 14486 -4427 14520
rect -4545 14452 -4427 14486
rect -4545 14418 -4503 14452
rect -4469 14418 -4427 14452
rect -4545 14384 -4427 14418
rect -4545 14350 -4503 14384
rect -4469 14350 -4427 14384
rect -4545 14316 -4427 14350
rect -4545 14282 -4503 14316
rect -4469 14282 -4427 14316
rect -4545 14248 -4427 14282
rect -4545 14214 -4503 14248
rect -4469 14214 -4427 14248
rect -4545 14180 -4427 14214
rect -4545 14146 -4503 14180
rect -4469 14146 -4427 14180
rect -4545 14112 -4427 14146
rect -4545 14078 -4503 14112
rect -4469 14078 -4427 14112
rect -4545 14044 -4427 14078
rect -4545 14010 -4503 14044
rect -4469 14010 -4427 14044
rect -4545 13976 -4427 14010
rect -4545 13942 -4503 13976
rect -4469 13942 -4427 13976
rect -4545 13908 -4427 13942
rect -4545 13874 -4503 13908
rect -4469 13874 -4427 13908
rect -4545 13840 -4427 13874
rect -4545 13806 -4503 13840
rect -4469 13806 -4427 13840
rect -4545 13772 -4427 13806
rect -4545 13738 -4503 13772
rect -4469 13738 -4427 13772
rect -4545 13704 -4427 13738
rect -4545 13670 -4503 13704
rect -4469 13670 -4427 13704
rect -4545 13636 -4427 13670
rect -4545 13602 -4503 13636
rect -4469 13602 -4427 13636
rect -4545 13568 -4427 13602
rect -4545 13534 -4503 13568
rect -4469 13534 -4427 13568
rect -4545 13500 -4427 13534
rect -4545 13466 -4503 13500
rect -4469 13466 -4427 13500
rect -4545 13432 -4427 13466
rect -4545 13398 -4503 13432
rect -4469 13398 -4427 13432
rect -4545 13364 -4427 13398
rect -4545 13330 -4503 13364
rect -4469 13330 -4427 13364
rect -4545 13296 -4427 13330
rect -4545 13262 -4503 13296
rect -4469 13262 -4427 13296
rect -4545 13228 -4427 13262
rect -4545 13194 -4503 13228
rect -4469 13194 -4427 13228
rect -4545 13160 -4427 13194
rect -4545 13126 -4503 13160
rect -4469 13126 -4427 13160
rect -4545 13092 -4427 13126
rect -4545 13058 -4503 13092
rect -4469 13058 -4427 13092
rect -4545 13024 -4427 13058
rect -4545 12990 -4503 13024
rect -4469 12990 -4427 13024
rect -4545 12956 -4427 12990
rect -4545 12922 -4503 12956
rect -4469 12922 -4427 12956
rect -4545 12888 -4427 12922
rect -4545 12854 -4503 12888
rect -4469 12854 -4427 12888
rect -7207 12719 -6645 12724
rect -6608 12729 -6457 12755
rect -6874 12707 -6646 12719
rect -7392 12637 -7246 12687
rect -6608 12695 -6547 12729
rect -6513 12695 -6457 12729
rect -7886 12588 -7753 12622
rect -7886 12554 -7843 12588
rect -7809 12554 -7753 12588
rect -7886 12520 -7753 12554
rect -7886 12486 -7843 12520
rect -7809 12486 -7753 12520
rect -7886 12452 -7753 12486
rect -7886 12418 -7843 12452
rect -7809 12418 -7753 12452
rect -7886 12384 -7753 12418
rect -7393 12552 -7245 12637
rect -7393 12518 -7339 12552
rect -7305 12518 -7245 12552
rect -7393 12480 -7245 12518
rect -7393 12446 -7339 12480
rect -7305 12446 -7245 12480
rect -7393 12400 -7245 12446
rect -6608 12560 -6457 12695
rect -6608 12526 -6550 12560
rect -6516 12526 -6457 12560
rect -6608 12488 -6457 12526
rect -6608 12454 -6550 12488
rect -6516 12454 -6457 12488
rect -6608 12401 -6457 12454
rect -6359 12724 -6211 12754
rect -6359 12690 -6310 12724
rect -6276 12690 -6211 12724
rect -6173 12718 -5616 12762
rect -4545 12820 -4427 12854
rect -4545 12786 -4503 12820
rect -4469 12786 -4427 12820
rect -5573 12726 -5428 12755
rect -4545 12752 -4427 12786
rect -6359 12562 -6211 12690
rect -6359 12528 -6310 12562
rect -6276 12528 -6211 12562
rect -6359 12490 -6211 12528
rect -6359 12456 -6310 12490
rect -6276 12456 -6211 12490
rect -6359 12403 -6211 12456
rect -5573 12692 -5516 12726
rect -5482 12692 -5428 12726
rect -5573 12557 -5428 12692
rect -5573 12523 -5531 12557
rect -5497 12523 -5428 12557
rect -5573 12485 -5428 12523
rect -5573 12451 -5531 12485
rect -5497 12451 -5428 12485
rect -5573 12403 -5428 12451
rect -5321 12726 -5165 12751
rect -5321 12692 -5261 12726
rect -5227 12692 -5165 12726
rect -5321 12570 -5165 12692
rect -5321 12536 -5262 12570
rect -5228 12536 -5165 12570
rect -5321 12498 -5165 12536
rect -5321 12464 -5262 12498
rect -5228 12464 -5165 12498
rect -5321 12403 -5165 12464
rect -4545 12718 -4503 12752
rect -4469 12718 -4427 12752
rect -4545 12684 -4427 12718
rect -4545 12650 -4503 12684
rect -4469 12650 -4427 12684
rect -4545 12616 -4427 12650
rect -4545 12582 -4503 12616
rect -4469 12582 -4427 12616
rect -4545 12548 -4427 12582
rect -4545 12514 -4503 12548
rect -4469 12514 -4427 12548
rect -4545 12480 -4427 12514
rect -4545 12446 -4503 12480
rect -4469 12446 -4427 12480
rect -4545 12412 -4427 12446
rect -7886 12350 -7843 12384
rect -7809 12350 -7753 12384
rect -7886 12278 -7753 12350
rect -4545 12378 -4503 12412
rect -4469 12378 -4427 12412
rect -4545 12344 -4427 12378
rect -4010 15001 -3896 15035
rect -3862 15001 -3828 15035
rect -3794 15001 -3680 15035
rect -4010 14914 -3976 15001
rect -3714 14914 -3680 15001
rect 10297 15011 10358 17061
rect 11256 15011 22482 17061
rect 23016 17312 23135 17346
rect 23169 17312 23203 17346
rect 23237 17312 23271 17346
rect 23305 17312 23339 17346
rect 23373 17312 23407 17346
rect 23441 17312 23475 17346
rect 23509 17312 23543 17346
rect 23577 17312 23611 17346
rect 23645 17312 23679 17346
rect 23713 17312 23747 17346
rect 23781 17312 23815 17346
rect 23849 17312 23883 17346
rect 23917 17312 23951 17346
rect 23985 17312 24019 17346
rect 24053 17312 24087 17346
rect 24121 17312 24155 17346
rect 24189 17312 24223 17346
rect 24257 17312 24376 17346
rect 23016 17231 23050 17312
rect 24342 17231 24376 17312
rect 23016 17163 23050 17197
rect 23196 17174 23237 17208
rect 23281 17174 23305 17208
rect 23353 17174 23373 17208
rect 23425 17174 23441 17208
rect 23497 17174 23509 17208
rect 23569 17174 23577 17208
rect 23641 17174 23645 17208
rect 23747 17174 23751 17208
rect 23815 17174 23823 17208
rect 23883 17174 23895 17208
rect 23951 17174 23967 17208
rect 24019 17174 24039 17208
rect 24087 17174 24111 17208
rect 24155 17174 24196 17208
rect 24342 17163 24376 17197
rect 23016 17095 23050 17129
rect 23016 17027 23050 17061
rect 23004 16993 23016 17004
rect 23150 17121 23184 17140
rect 23150 17049 23184 17061
rect 23050 16993 23150 17004
rect 24208 17121 24242 17140
rect 24208 17049 24242 17061
rect 23184 16993 23190 17004
rect 23004 16977 23190 16993
rect 23004 16959 23150 16977
rect 23004 16925 23016 16959
rect 23050 16925 23150 16959
rect 23184 16925 23190 16977
rect 23004 16905 23190 16925
rect 23004 16891 23150 16905
rect 23004 16863 23016 16891
rect 23050 16863 23150 16891
rect 23016 16823 23050 16857
rect 23016 16755 23050 16789
rect 23016 16687 23050 16721
rect 23016 16619 23050 16653
rect 23016 16551 23050 16585
rect 23004 16517 23016 16541
rect 23184 16863 23190 16905
rect 24208 16977 24242 16993
rect 24208 16905 24242 16925
rect 23150 16833 23184 16857
rect 23150 16761 23184 16789
rect 23150 16689 23184 16721
rect 23150 16619 23184 16653
rect 23150 16551 23184 16583
rect 23050 16517 23150 16541
rect 24208 16833 24242 16857
rect 24208 16761 24242 16789
rect 24342 17095 24376 17129
rect 24342 17027 24376 17061
rect 24342 16959 24376 16993
rect 24558 17284 24592 17318
rect 24558 17216 24592 17250
rect 24558 17148 24592 17182
rect 24726 18362 24738 18372
rect 25750 18508 25784 18542
rect 25750 18440 25784 18470
rect 25750 18372 25784 18398
rect 24692 18304 24726 18326
rect 24692 18236 24726 18254
rect 24692 18168 24726 18182
rect 24692 18100 24726 18110
rect 24692 18032 24726 18038
rect 24692 17964 24726 17966
rect 24692 17928 24726 17930
rect 24692 17856 24726 17862
rect 24692 17784 24726 17794
rect 24692 17712 24726 17726
rect 24692 17640 24726 17658
rect 24692 17568 24726 17590
rect 24692 17496 24726 17522
rect 24692 17424 24726 17454
rect 24692 17352 24726 17386
rect 24692 17284 24726 17318
rect 24692 17216 24726 17246
rect 24692 17143 24726 17174
rect 25750 18304 25784 18326
rect 25750 18236 25784 18254
rect 25750 18168 25784 18182
rect 25750 18100 25784 18110
rect 25750 18032 25784 18038
rect 25750 17964 25784 17966
rect 25750 17928 25784 17930
rect 25750 17856 25784 17862
rect 25750 17784 25784 17794
rect 25750 17712 25784 17726
rect 25750 17640 25784 17658
rect 25750 17568 25784 17590
rect 25750 17496 25784 17522
rect 25750 17424 25784 17454
rect 25750 17352 25784 17386
rect 25750 17284 25784 17318
rect 25750 17216 25784 17246
rect 25750 17143 25784 17174
rect 26808 18720 26842 18751
rect 26808 18648 26842 18678
rect 26808 18576 26842 18610
rect 26808 18508 26842 18542
rect 26808 18440 26842 18470
rect 26808 18372 26842 18398
rect 26808 18304 26842 18326
rect 26808 18236 26842 18254
rect 26808 18168 26842 18182
rect 26808 18100 26842 18110
rect 26808 18032 26842 18038
rect 26808 17964 26842 17966
rect 26808 17928 26842 17930
rect 26808 17856 26842 17862
rect 26808 17784 26842 17794
rect 26808 17712 26842 17726
rect 26808 17640 26842 17658
rect 26808 17568 26842 17590
rect 26808 17496 26842 17522
rect 26808 17424 26842 17454
rect 26808 17352 26842 17386
rect 26808 17284 26842 17318
rect 26808 17216 26842 17246
rect 26808 17143 26842 17174
rect 27866 18720 27900 18751
rect 27866 18648 27900 18678
rect 27866 18576 27900 18610
rect 27866 18508 27900 18542
rect 27866 18440 27900 18470
rect 27866 18372 27900 18398
rect 27866 18304 27900 18326
rect 27866 18236 27900 18254
rect 27866 18168 27900 18182
rect 27866 18100 27900 18110
rect 27866 18032 27900 18038
rect 27866 17964 27900 17966
rect 27866 17928 27900 17930
rect 27866 17856 27900 17862
rect 27866 17784 27900 17794
rect 27866 17712 27900 17726
rect 27866 17640 27900 17658
rect 27866 17568 27900 17590
rect 27866 17496 27900 17522
rect 27866 17424 27900 17454
rect 27866 17352 27900 17386
rect 27866 17284 27900 17318
rect 27866 17216 27900 17246
rect 27866 17143 27900 17174
rect 28000 18712 28034 18746
rect 28000 18644 28034 18678
rect 28000 18576 28034 18610
rect 28000 18508 28034 18542
rect 40682 18535 40923 19006
rect 42341 19003 45374 19006
rect 28000 18440 28034 18474
rect 28000 18372 28034 18406
rect 28000 18304 28034 18338
rect 28000 18236 28034 18270
rect 38775 18294 40923 18535
rect 42478 18948 42512 19003
rect 45326 18948 45360 19003
rect 42478 18880 42512 18914
rect 42658 18890 42705 18924
rect 42741 18890 42775 18924
rect 42811 18890 42858 18924
rect 42916 18890 42963 18924
rect 42999 18890 43033 18924
rect 43069 18890 43116 18924
rect 43174 18890 43221 18924
rect 43257 18890 43291 18924
rect 43327 18890 43374 18924
rect 43432 18890 43479 18924
rect 43515 18890 43549 18924
rect 43585 18890 43632 18924
rect 43690 18890 43737 18924
rect 43773 18890 43807 18924
rect 43843 18890 43890 18924
rect 43948 18890 43995 18924
rect 44031 18890 44065 18924
rect 44101 18890 44148 18924
rect 44206 18890 44253 18924
rect 44289 18890 44323 18924
rect 44359 18890 44406 18924
rect 44464 18890 44511 18924
rect 44547 18890 44581 18924
rect 44617 18890 44664 18924
rect 44722 18890 44769 18924
rect 44805 18890 44839 18924
rect 44875 18890 44922 18924
rect 44980 18890 45027 18924
rect 45063 18890 45097 18924
rect 45133 18890 45180 18924
rect 45326 18880 45360 18914
rect 42478 18812 42512 18846
rect 42478 18744 42512 18778
rect 42478 18676 42512 18710
rect 42478 18608 42512 18642
rect 42478 18540 42512 18574
rect 42478 18472 42512 18506
rect 42478 18404 42512 18438
rect 42478 18336 42512 18370
rect 38775 18291 40146 18294
rect 38775 18286 39353 18291
rect 39387 18286 39425 18291
rect 39459 18286 40146 18291
rect 38775 18252 38890 18286
rect 38924 18252 38958 18286
rect 38992 18252 39026 18286
rect 39060 18252 39094 18286
rect 39128 18252 39162 18286
rect 39196 18252 39230 18286
rect 39264 18252 39298 18286
rect 39332 18257 39353 18286
rect 39400 18257 39425 18286
rect 39332 18252 39366 18257
rect 39400 18252 39434 18257
rect 39468 18252 39502 18286
rect 39536 18252 39570 18286
rect 39604 18252 39638 18286
rect 39672 18252 39706 18286
rect 39740 18252 39774 18286
rect 39808 18252 39842 18286
rect 39876 18252 39910 18286
rect 39944 18252 39978 18286
rect 40012 18252 40146 18286
rect 38775 18228 40146 18252
rect 28000 18168 28034 18202
rect 28000 18100 28034 18134
rect 28000 18032 28034 18066
rect 28000 17964 28034 17998
rect 28000 17896 28034 17930
rect 28000 17828 28034 17862
rect 28000 17760 28034 17794
rect 28000 17692 28034 17726
rect 28000 17624 28034 17658
rect 28000 17556 28034 17590
rect 28000 17488 28034 17522
rect 28000 17420 28034 17454
rect 28000 17352 28034 17386
rect 28000 17284 28034 17318
rect 28000 17216 28034 17250
rect 28000 17148 28034 17182
rect 24558 17080 24592 17114
rect 24738 17066 24779 17100
rect 24823 17066 24847 17100
rect 24895 17066 24915 17100
rect 24967 17066 24983 17100
rect 25039 17066 25051 17100
rect 25111 17066 25119 17100
rect 25183 17066 25187 17100
rect 25289 17066 25293 17100
rect 25357 17066 25365 17100
rect 25425 17066 25437 17100
rect 25493 17066 25509 17100
rect 25561 17066 25581 17100
rect 25629 17066 25653 17100
rect 25697 17066 25738 17100
rect 25796 17066 25837 17100
rect 25881 17066 25905 17100
rect 25953 17066 25973 17100
rect 26025 17066 26041 17100
rect 26097 17066 26109 17100
rect 26169 17066 26177 17100
rect 26241 17066 26245 17100
rect 26347 17066 26351 17100
rect 26415 17066 26423 17100
rect 26483 17066 26495 17100
rect 26551 17066 26567 17100
rect 26619 17066 26639 17100
rect 26687 17066 26711 17100
rect 26755 17066 26796 17100
rect 26854 17066 26895 17100
rect 26939 17066 26963 17100
rect 27011 17066 27031 17100
rect 27083 17066 27099 17100
rect 27155 17066 27167 17100
rect 27227 17066 27235 17100
rect 27299 17066 27303 17100
rect 27405 17066 27409 17100
rect 27473 17066 27481 17100
rect 27541 17066 27553 17100
rect 27609 17066 27625 17100
rect 27677 17066 27697 17100
rect 27745 17066 27769 17100
rect 27813 17066 27854 17100
rect 28000 17080 28034 17114
rect 24558 16962 24592 17046
rect 28000 16962 28034 17046
rect 24558 16928 24681 16962
rect 24715 16928 24749 16962
rect 24783 16928 24817 16962
rect 24851 16928 24885 16962
rect 24919 16928 24953 16962
rect 24987 16928 25021 16962
rect 25055 16928 25089 16962
rect 25123 16928 25157 16962
rect 25191 16928 25225 16962
rect 25259 16928 25293 16962
rect 25327 16928 25361 16962
rect 25395 16928 25429 16962
rect 25463 16928 25497 16962
rect 25531 16928 25565 16962
rect 25599 16928 25633 16962
rect 25667 16928 25701 16962
rect 25735 16928 25769 16962
rect 25803 16928 25837 16962
rect 25871 16928 25905 16962
rect 25939 16928 25973 16962
rect 26007 16928 26041 16962
rect 26075 16928 26109 16962
rect 26143 16928 26177 16962
rect 26211 16928 26245 16962
rect 26279 16928 26313 16962
rect 26347 16928 26381 16962
rect 26415 16928 26449 16962
rect 26483 16928 26517 16962
rect 26551 16928 26585 16962
rect 26619 16928 26653 16962
rect 26687 16928 26721 16962
rect 26755 16928 26789 16962
rect 26823 16928 26857 16962
rect 26891 16928 26925 16962
rect 26959 16928 26993 16962
rect 27027 16928 27061 16962
rect 27095 16928 27129 16962
rect 27163 16928 27197 16962
rect 27231 16928 27265 16962
rect 27299 16928 27333 16962
rect 27367 16928 27401 16962
rect 27435 16928 27469 16962
rect 27503 16928 27537 16962
rect 27571 16928 27605 16962
rect 27639 16928 27673 16962
rect 27707 16928 27741 16962
rect 27775 16928 27809 16962
rect 27843 16928 27877 16962
rect 27911 16928 28034 16962
rect 38776 18191 38856 18228
rect 39316 18204 39496 18228
rect 40066 18211 40146 18228
rect 38776 18157 38794 18191
rect 38828 18157 38856 18191
rect 38776 18123 38856 18157
rect 38776 18089 38794 18123
rect 38828 18089 38856 18123
rect 38776 18055 38856 18089
rect 40066 18177 40084 18211
rect 40118 18177 40146 18211
rect 40066 18143 40146 18177
rect 40066 18109 40084 18143
rect 40118 18109 40146 18143
rect 40066 18075 40146 18109
rect 38776 18021 38794 18055
rect 38828 18021 38856 18055
rect 39190 18021 39237 18055
rect 39273 18021 39307 18055
rect 39343 18021 39390 18055
rect 39448 18021 39495 18055
rect 39531 18021 39565 18055
rect 39601 18021 39648 18055
rect 40066 18041 40084 18075
rect 40118 18041 40146 18075
rect 38776 17987 38856 18021
rect 38776 17953 38794 17987
rect 38828 17953 38856 17987
rect 40066 18007 40146 18041
rect 38776 17919 38856 17953
rect 38776 17885 38794 17919
rect 38828 17885 38856 17919
rect 38776 17851 38856 17885
rect 38776 17817 38794 17851
rect 38828 17817 38856 17851
rect 38776 17783 38856 17817
rect 38776 17749 38794 17783
rect 38828 17749 38856 17783
rect 38776 17715 38856 17749
rect 38776 17681 38794 17715
rect 38828 17681 38856 17715
rect 38776 17647 38856 17681
rect 38776 17613 38794 17647
rect 38828 17613 38856 17647
rect 38776 17579 38856 17613
rect 38776 17545 38794 17579
rect 38828 17545 38856 17579
rect 38776 17511 38856 17545
rect 38776 17477 38794 17511
rect 38828 17477 38856 17511
rect 38776 17443 38856 17477
rect 38776 17409 38794 17443
rect 38828 17409 38856 17443
rect 38776 17375 38856 17409
rect 38776 17341 38794 17375
rect 38828 17341 38856 17375
rect 38776 17307 38856 17341
rect 38776 17273 38794 17307
rect 38828 17273 38856 17307
rect 38776 17239 38856 17273
rect 38776 17205 38794 17239
rect 38828 17205 38856 17239
rect 38776 17171 38856 17205
rect 38776 17137 38794 17171
rect 38828 17137 38856 17171
rect 38776 17103 38856 17137
rect 38776 17069 38794 17103
rect 38828 17069 38856 17103
rect 38776 17035 38856 17069
rect 38776 17001 38794 17035
rect 38828 17001 38856 17035
rect 38776 16967 38856 17001
rect 39144 17959 39178 17978
rect 39144 17887 39178 17899
rect 39144 17815 39178 17831
rect 39144 17743 39178 17763
rect 39144 17671 39178 17695
rect 39144 17599 39178 17627
rect 39144 17527 39178 17559
rect 39144 17457 39178 17491
rect 39144 17389 39178 17421
rect 39144 17321 39178 17349
rect 39144 17253 39178 17277
rect 39144 17185 39178 17205
rect 39144 17117 39178 17133
rect 39144 17049 39178 17061
rect 39144 16970 39178 16989
rect 39402 17959 39436 17978
rect 39402 17887 39436 17899
rect 39402 17815 39436 17831
rect 39402 17743 39436 17763
rect 39402 17671 39436 17695
rect 39402 17599 39436 17627
rect 39402 17527 39436 17559
rect 39402 17457 39436 17491
rect 39402 17389 39436 17421
rect 39402 17321 39436 17349
rect 39402 17253 39436 17277
rect 39402 17185 39436 17205
rect 39402 17117 39436 17133
rect 39402 17049 39436 17061
rect 39402 16970 39436 16989
rect 39660 17959 39694 17978
rect 39660 17887 39694 17899
rect 39660 17815 39694 17831
rect 39660 17743 39694 17763
rect 39660 17671 39694 17695
rect 39660 17599 39694 17627
rect 39660 17527 39694 17559
rect 39660 17457 39694 17491
rect 39660 17389 39694 17421
rect 39660 17321 39694 17349
rect 39660 17253 39694 17277
rect 39660 17185 39694 17205
rect 39660 17117 39694 17133
rect 39660 17049 39694 17061
rect 39660 16970 39694 16989
rect 40066 17973 40084 18007
rect 40118 17973 40146 18007
rect 40066 17939 40146 17973
rect 40066 17905 40084 17939
rect 40118 17905 40146 17939
rect 40066 17871 40146 17905
rect 40066 17837 40084 17871
rect 40118 17837 40146 17871
rect 40066 17803 40146 17837
rect 40066 17769 40084 17803
rect 40118 17769 40146 17803
rect 40066 17735 40146 17769
rect 40066 17701 40084 17735
rect 40118 17701 40146 17735
rect 40066 17667 40146 17701
rect 40066 17633 40084 17667
rect 40118 17633 40146 17667
rect 40066 17599 40146 17633
rect 40066 17565 40084 17599
rect 40118 17565 40146 17599
rect 40066 17531 40146 17565
rect 40066 17497 40084 17531
rect 40118 17497 40146 17531
rect 40066 17463 40146 17497
rect 40066 17429 40084 17463
rect 40118 17429 40146 17463
rect 40066 17395 40146 17429
rect 40066 17361 40084 17395
rect 40118 17361 40146 17395
rect 40066 17327 40146 17361
rect 40066 17293 40084 17327
rect 40118 17293 40146 17327
rect 40066 17259 40146 17293
rect 40066 17225 40084 17259
rect 40118 17225 40146 17259
rect 40066 17191 40146 17225
rect 40066 17157 40084 17191
rect 40118 17157 40146 17191
rect 40066 17123 40146 17157
rect 40066 17089 40084 17123
rect 40118 17089 40146 17123
rect 40066 17055 40146 17089
rect 40066 17021 40084 17055
rect 40118 17021 40146 17055
rect 40066 16987 40146 17021
rect 38776 16933 38794 16967
rect 38828 16933 38856 16967
rect 24342 16891 24376 16925
rect 24342 16823 24376 16857
rect 24342 16755 24376 16789
rect 24208 16689 24242 16721
rect 24208 16619 24242 16653
rect 24208 16551 24242 16583
rect 24330 16721 24342 16750
rect 38776 16899 38856 16933
rect 40066 16953 40084 16987
rect 40118 16953 40146 16987
rect 38776 16865 38794 16899
rect 38828 16865 38856 16899
rect 39190 16893 39237 16927
rect 39273 16893 39307 16927
rect 39343 16893 39390 16927
rect 39448 16893 39495 16927
rect 39531 16893 39565 16927
rect 39601 16893 39648 16927
rect 40066 16919 40146 16953
rect 38776 16831 38856 16865
rect 38776 16797 38794 16831
rect 38828 16797 38856 16831
rect 38776 16774 38856 16797
rect 40066 16885 40084 16919
rect 40118 16885 40146 16919
rect 40066 16851 40146 16885
rect 40066 16817 40084 16851
rect 40118 16817 40146 16851
rect 40066 16774 40146 16817
rect 24376 16721 24559 16750
rect 24330 16716 24559 16721
rect 24593 16716 24627 16750
rect 24661 16716 24695 16750
rect 24729 16716 24763 16750
rect 24797 16716 24831 16750
rect 24865 16716 24899 16750
rect 24933 16716 24967 16750
rect 25001 16716 25035 16750
rect 25069 16716 25103 16750
rect 25137 16716 25171 16750
rect 25205 16716 25239 16750
rect 25273 16716 25307 16750
rect 25341 16716 25375 16750
rect 25409 16716 25443 16750
rect 25477 16716 25511 16750
rect 25545 16716 25579 16750
rect 25613 16716 25647 16750
rect 25681 16716 25715 16750
rect 25749 16716 25783 16750
rect 25817 16716 25851 16750
rect 25885 16716 25919 16750
rect 25953 16716 25987 16750
rect 26021 16716 26055 16750
rect 26089 16716 26123 16750
rect 26157 16716 26191 16750
rect 26225 16716 26259 16750
rect 26293 16716 26327 16750
rect 26361 16716 26395 16750
rect 26429 16716 26463 16750
rect 26497 16716 26531 16750
rect 26565 16716 26599 16750
rect 26633 16716 26667 16750
rect 26701 16716 26735 16750
rect 26769 16716 26803 16750
rect 26837 16716 26871 16750
rect 26905 16716 26939 16750
rect 26973 16716 27007 16750
rect 27041 16716 27075 16750
rect 27109 16716 27143 16750
rect 27177 16716 27211 16750
rect 27245 16716 27279 16750
rect 27313 16716 27347 16750
rect 27381 16716 27415 16750
rect 27449 16716 27483 16750
rect 27517 16716 27551 16750
rect 27585 16716 27684 16750
rect 24330 16687 25021 16716
rect 24330 16653 24342 16687
rect 24376 16653 25021 16687
rect 24330 16646 25021 16653
rect 24330 16619 24460 16646
rect 24330 16585 24342 16619
rect 24376 16612 24460 16619
rect 24494 16620 25021 16646
rect 27122 16620 27554 16716
rect 24494 16612 24590 16620
rect 24376 16585 24590 16612
rect 24330 16578 24590 16585
rect 24330 16551 24460 16578
rect 24330 16550 24342 16551
rect 23004 16511 23150 16517
rect 23184 16511 23190 16541
rect 23004 16483 23190 16511
rect 23004 16449 23016 16483
rect 23050 16449 23150 16483
rect 23004 16439 23150 16449
rect 23184 16439 23190 16483
rect 23004 16415 23190 16439
rect 23004 16400 23016 16415
rect 23050 16400 23150 16415
rect 23016 16347 23050 16381
rect 23016 16279 23050 16313
rect 23016 16211 23050 16245
rect 23016 16143 23050 16177
rect 23184 16400 23190 16415
rect 24208 16483 24242 16511
rect 24208 16415 24242 16439
rect 23150 16347 23184 16367
rect 23150 16279 23184 16295
rect 23150 16211 23184 16223
rect 23150 16132 23184 16151
rect 24208 16347 24242 16367
rect 24208 16279 24242 16295
rect 24208 16211 24242 16223
rect 24208 16132 24242 16151
rect 24376 16550 24460 16551
rect 24342 16483 24376 16517
rect 24342 16415 24376 16449
rect 24342 16347 24376 16381
rect 24342 16279 24376 16313
rect 24342 16211 24376 16245
rect 24342 16143 24376 16177
rect 23016 16075 23050 16109
rect 23196 16064 23237 16098
rect 23281 16064 23305 16098
rect 23353 16064 23373 16098
rect 23425 16064 23441 16098
rect 23497 16064 23509 16098
rect 23569 16064 23577 16098
rect 23641 16064 23645 16098
rect 23747 16064 23751 16098
rect 23815 16064 23823 16098
rect 23883 16064 23895 16098
rect 23951 16064 23967 16098
rect 24019 16064 24039 16098
rect 24087 16064 24111 16098
rect 24155 16064 24196 16098
rect 24342 16075 24376 16109
rect 23016 15960 23050 16041
rect 24342 15960 24376 16041
rect 23016 15926 23135 15960
rect 23169 15926 23203 15960
rect 23237 15926 23271 15960
rect 23305 15926 23339 15960
rect 23373 15926 23407 15960
rect 23441 15926 23475 15960
rect 23509 15926 23543 15960
rect 23577 15926 23611 15960
rect 23645 15926 23679 15960
rect 23713 15926 23747 15960
rect 23781 15926 23815 15960
rect 23849 15926 23883 15960
rect 23917 15926 23951 15960
rect 23985 15926 24019 15960
rect 24053 15926 24087 15960
rect 24121 15926 24155 15960
rect 24189 15926 24223 15960
rect 24257 15926 24376 15960
rect 24494 16550 24590 16578
rect 27650 16646 27684 16716
rect 38776 16746 40146 16774
rect 38776 16712 38910 16746
rect 38944 16712 38978 16746
rect 39012 16712 39046 16746
rect 39080 16712 39114 16746
rect 39148 16712 39182 16746
rect 39216 16712 39250 16746
rect 39284 16712 39318 16746
rect 39352 16712 39386 16746
rect 39420 16712 39454 16746
rect 39488 16712 39522 16746
rect 39556 16712 39590 16746
rect 39624 16712 39658 16746
rect 39692 16712 39726 16746
rect 39760 16712 39794 16746
rect 39828 16712 39862 16746
rect 39896 16712 39930 16746
rect 39964 16712 39998 16746
rect 40032 16712 40146 16746
rect 38776 16694 40146 16712
rect 42478 18268 42512 18302
rect 42478 18200 42512 18234
rect 42478 18132 42512 18166
rect 42478 18064 42512 18098
rect 42478 17996 42512 18030
rect 42478 17928 42512 17962
rect 42478 17860 42512 17894
rect 42478 17792 42512 17826
rect 42478 17724 42512 17758
rect 42478 17656 42512 17690
rect 42478 17588 42512 17622
rect 42478 17520 42512 17554
rect 42478 17452 42512 17486
rect 42478 17384 42512 17418
rect 42478 17316 42512 17350
rect 42478 17248 42512 17282
rect 42478 17180 42512 17214
rect 42478 17112 42512 17146
rect 42478 17044 42512 17078
rect 42478 16976 42512 17010
rect 42478 16908 42512 16942
rect 42478 16840 42512 16874
rect 42612 18812 42646 18847
rect 42612 18744 42646 18762
rect 42612 18676 42646 18690
rect 42612 18608 42646 18618
rect 42612 18540 42646 18546
rect 42612 18472 42646 18474
rect 42612 18436 42646 18438
rect 42612 18364 42646 18370
rect 42612 18292 42646 18302
rect 42612 18220 42646 18234
rect 42612 18148 42646 18166
rect 42612 18076 42646 18098
rect 42612 18004 42646 18030
rect 42612 17932 42646 17962
rect 42612 17860 42646 17894
rect 42612 17792 42646 17826
rect 42612 17724 42646 17754
rect 42612 17656 42646 17682
rect 42612 17588 42646 17610
rect 42612 17520 42646 17538
rect 42612 17452 42646 17466
rect 42612 17384 42646 17394
rect 42612 17316 42646 17322
rect 42612 17248 42646 17250
rect 42612 17212 42646 17214
rect 42612 17140 42646 17146
rect 42612 17068 42646 17078
rect 42612 16996 42646 17010
rect 42612 16924 42646 16942
rect 42612 16839 42646 16874
rect 42870 18812 42904 18847
rect 42870 18744 42904 18762
rect 42870 18676 42904 18690
rect 42870 18608 42904 18618
rect 42870 18540 42904 18546
rect 42870 18472 42904 18474
rect 42870 18436 42904 18438
rect 42870 18364 42904 18370
rect 42870 18292 42904 18302
rect 42870 18220 42904 18234
rect 42870 18148 42904 18166
rect 42870 18076 42904 18098
rect 42870 18004 42904 18030
rect 42870 17932 42904 17962
rect 42870 17860 42904 17894
rect 42870 17792 42904 17826
rect 42870 17724 42904 17754
rect 42870 17656 42904 17682
rect 42870 17588 42904 17610
rect 42870 17520 42904 17538
rect 42870 17452 42904 17466
rect 42870 17384 42904 17394
rect 42870 17316 42904 17322
rect 42870 17248 42904 17250
rect 42870 17212 42904 17214
rect 42870 17140 42904 17146
rect 42870 17068 42904 17078
rect 42870 16996 42904 17010
rect 42870 16924 42904 16942
rect 42870 16839 42904 16874
rect 43128 18812 43162 18847
rect 43128 18744 43162 18762
rect 43128 18676 43162 18690
rect 43128 18608 43162 18618
rect 43128 18540 43162 18546
rect 43128 18472 43162 18474
rect 43128 18436 43162 18438
rect 43128 18364 43162 18370
rect 43128 18292 43162 18302
rect 43128 18220 43162 18234
rect 43128 18148 43162 18166
rect 43128 18076 43162 18098
rect 43128 18004 43162 18030
rect 43128 17932 43162 17962
rect 43128 17860 43162 17894
rect 43128 17792 43162 17826
rect 43128 17724 43162 17754
rect 43128 17656 43162 17682
rect 43128 17588 43162 17610
rect 43128 17520 43162 17538
rect 43128 17452 43162 17466
rect 43128 17384 43162 17394
rect 43128 17316 43162 17322
rect 43128 17248 43162 17250
rect 43128 17212 43162 17214
rect 43128 17140 43162 17146
rect 43128 17068 43162 17078
rect 43128 16996 43162 17010
rect 43128 16924 43162 16942
rect 43128 16839 43162 16874
rect 43386 18812 43420 18847
rect 43386 18744 43420 18762
rect 43386 18676 43420 18690
rect 43386 18608 43420 18618
rect 43386 18540 43420 18546
rect 43386 18472 43420 18474
rect 43386 18436 43420 18438
rect 43386 18364 43420 18370
rect 43386 18292 43420 18302
rect 43386 18220 43420 18234
rect 43386 18148 43420 18166
rect 43386 18076 43420 18098
rect 43386 18004 43420 18030
rect 43386 17932 43420 17962
rect 43386 17860 43420 17894
rect 43386 17792 43420 17826
rect 43386 17724 43420 17754
rect 43386 17656 43420 17682
rect 43386 17588 43420 17610
rect 43386 17520 43420 17538
rect 43386 17452 43420 17466
rect 43386 17384 43420 17394
rect 43386 17316 43420 17322
rect 43386 17248 43420 17250
rect 43386 17212 43420 17214
rect 43386 17140 43420 17146
rect 43386 17068 43420 17078
rect 43386 16996 43420 17010
rect 43386 16924 43420 16942
rect 43386 16839 43420 16874
rect 43644 18812 43678 18847
rect 43644 18744 43678 18762
rect 43644 18676 43678 18690
rect 43644 18608 43678 18618
rect 43644 18540 43678 18546
rect 43644 18472 43678 18474
rect 43644 18436 43678 18438
rect 43644 18364 43678 18370
rect 43644 18292 43678 18302
rect 43644 18220 43678 18234
rect 43644 18148 43678 18166
rect 43644 18076 43678 18098
rect 43644 18004 43678 18030
rect 43644 17932 43678 17962
rect 43644 17860 43678 17894
rect 43644 17792 43678 17826
rect 43644 17724 43678 17754
rect 43644 17656 43678 17682
rect 43644 17588 43678 17610
rect 43644 17520 43678 17538
rect 43644 17452 43678 17466
rect 43644 17384 43678 17394
rect 43644 17316 43678 17322
rect 43644 17248 43678 17250
rect 43644 17212 43678 17214
rect 43644 17140 43678 17146
rect 43644 17068 43678 17078
rect 43644 16996 43678 17010
rect 43644 16924 43678 16942
rect 43644 16839 43678 16874
rect 43902 18812 43936 18847
rect 43902 18744 43936 18762
rect 43902 18676 43936 18690
rect 43902 18608 43936 18618
rect 43902 18540 43936 18546
rect 43902 18472 43936 18474
rect 43902 18436 43936 18438
rect 43902 18364 43936 18370
rect 43902 18292 43936 18302
rect 43902 18220 43936 18234
rect 43902 18148 43936 18166
rect 43902 18076 43936 18098
rect 43902 18004 43936 18030
rect 43902 17932 43936 17962
rect 43902 17860 43936 17894
rect 43902 17792 43936 17826
rect 43902 17724 43936 17754
rect 43902 17656 43936 17682
rect 43902 17588 43936 17610
rect 43902 17520 43936 17538
rect 43902 17452 43936 17466
rect 43902 17384 43936 17394
rect 43902 17316 43936 17322
rect 43902 17248 43936 17250
rect 43902 17212 43936 17214
rect 43902 17140 43936 17146
rect 43902 17068 43936 17078
rect 43902 16996 43936 17010
rect 43902 16924 43936 16942
rect 43902 16839 43936 16874
rect 44160 18812 44194 18847
rect 44160 18744 44194 18762
rect 44160 18676 44194 18690
rect 44160 18608 44194 18618
rect 44160 18540 44194 18546
rect 44160 18472 44194 18474
rect 44160 18436 44194 18438
rect 44160 18364 44194 18370
rect 44160 18292 44194 18302
rect 44160 18220 44194 18234
rect 44160 18148 44194 18166
rect 44160 18076 44194 18098
rect 44160 18004 44194 18030
rect 44160 17932 44194 17962
rect 44160 17860 44194 17894
rect 44160 17792 44194 17826
rect 44160 17724 44194 17754
rect 44160 17656 44194 17682
rect 44160 17588 44194 17610
rect 44160 17520 44194 17538
rect 44160 17452 44194 17466
rect 44160 17384 44194 17394
rect 44160 17316 44194 17322
rect 44160 17248 44194 17250
rect 44160 17212 44194 17214
rect 44160 17140 44194 17146
rect 44160 17068 44194 17078
rect 44160 16996 44194 17010
rect 44160 16924 44194 16942
rect 44160 16839 44194 16874
rect 44418 18812 44452 18847
rect 44418 18744 44452 18762
rect 44418 18676 44452 18690
rect 44418 18608 44452 18618
rect 44418 18540 44452 18546
rect 44418 18472 44452 18474
rect 44418 18436 44452 18438
rect 44418 18364 44452 18370
rect 44418 18292 44452 18302
rect 44418 18220 44452 18234
rect 44418 18148 44452 18166
rect 44418 18076 44452 18098
rect 44418 18004 44452 18030
rect 44418 17932 44452 17962
rect 44418 17860 44452 17894
rect 44418 17792 44452 17826
rect 44418 17724 44452 17754
rect 44418 17656 44452 17682
rect 44418 17588 44452 17610
rect 44418 17520 44452 17538
rect 44418 17452 44452 17466
rect 44418 17384 44452 17394
rect 44418 17316 44452 17322
rect 44418 17248 44452 17250
rect 44418 17212 44452 17214
rect 44418 17140 44452 17146
rect 44418 17068 44452 17078
rect 44418 16996 44452 17010
rect 44418 16924 44452 16942
rect 44418 16839 44452 16874
rect 44676 18812 44710 18847
rect 44676 18744 44710 18762
rect 44676 18676 44710 18690
rect 44676 18608 44710 18618
rect 44676 18540 44710 18546
rect 44676 18472 44710 18474
rect 44676 18436 44710 18438
rect 44676 18364 44710 18370
rect 44676 18292 44710 18302
rect 44676 18220 44710 18234
rect 44676 18148 44710 18166
rect 44676 18076 44710 18098
rect 44676 18004 44710 18030
rect 44676 17932 44710 17962
rect 44676 17860 44710 17894
rect 44676 17792 44710 17826
rect 44676 17724 44710 17754
rect 44676 17656 44710 17682
rect 44676 17588 44710 17610
rect 44676 17520 44710 17538
rect 44676 17452 44710 17466
rect 44676 17384 44710 17394
rect 44676 17316 44710 17322
rect 44676 17248 44710 17250
rect 44676 17212 44710 17214
rect 44676 17140 44710 17146
rect 44676 17068 44710 17078
rect 44676 16996 44710 17010
rect 44676 16924 44710 16942
rect 44676 16839 44710 16874
rect 44934 18812 44968 18847
rect 44934 18744 44968 18762
rect 44934 18676 44968 18690
rect 44934 18608 44968 18618
rect 44934 18540 44968 18546
rect 44934 18472 44968 18474
rect 44934 18436 44968 18438
rect 44934 18364 44968 18370
rect 44934 18292 44968 18302
rect 44934 18220 44968 18234
rect 44934 18148 44968 18166
rect 44934 18076 44968 18098
rect 44934 18004 44968 18030
rect 44934 17932 44968 17962
rect 44934 17860 44968 17894
rect 44934 17792 44968 17826
rect 44934 17724 44968 17754
rect 44934 17656 44968 17682
rect 44934 17588 44968 17610
rect 44934 17520 44968 17538
rect 44934 17452 44968 17466
rect 44934 17384 44968 17394
rect 44934 17316 44968 17322
rect 44934 17248 44968 17250
rect 44934 17212 44968 17214
rect 44934 17140 44968 17146
rect 44934 17068 44968 17078
rect 44934 16996 44968 17010
rect 44934 16924 44968 16942
rect 44934 16839 44968 16874
rect 45192 18812 45226 18847
rect 45192 18744 45226 18762
rect 45192 18676 45226 18690
rect 45192 18608 45226 18618
rect 45192 18540 45226 18546
rect 45192 18472 45226 18474
rect 45192 18436 45226 18438
rect 45192 18364 45226 18370
rect 45192 18292 45226 18302
rect 45192 18220 45226 18234
rect 45192 18148 45226 18166
rect 45192 18076 45226 18098
rect 45192 18004 45226 18030
rect 45192 17932 45226 17962
rect 45192 17860 45226 17894
rect 45192 17792 45226 17826
rect 45192 17724 45226 17754
rect 45192 17656 45226 17682
rect 45192 17588 45226 17610
rect 45192 17520 45226 17538
rect 45192 17452 45226 17466
rect 45192 17384 45226 17394
rect 45192 17316 45226 17322
rect 45192 17248 45226 17250
rect 45192 17212 45226 17214
rect 45192 17140 45226 17146
rect 45192 17068 45226 17078
rect 45192 16996 45226 17010
rect 45192 16924 45226 16942
rect 45192 16839 45226 16874
rect 45326 18812 45360 18846
rect 45326 18744 45360 18778
rect 45326 18676 45360 18710
rect 45326 18608 45360 18642
rect 45326 18540 45360 18574
rect 45326 18472 45360 18506
rect 45326 18404 45360 18438
rect 45326 18336 45360 18370
rect 45326 18268 45360 18302
rect 45326 18200 45360 18234
rect 45326 18132 45360 18166
rect 45326 18064 45360 18098
rect 45326 17996 45360 18030
rect 45326 17928 45360 17962
rect 45326 17860 45360 17894
rect 45326 17792 45360 17826
rect 45326 17724 45360 17758
rect 45326 17656 45360 17690
rect 45326 17588 45360 17622
rect 45326 17520 45360 17554
rect 45326 17452 45360 17486
rect 45326 17384 45360 17418
rect 45326 17316 45360 17350
rect 45326 17248 45360 17282
rect 45326 17180 45360 17214
rect 45326 17112 45360 17146
rect 45326 17044 45360 17078
rect 45326 16976 45360 17010
rect 45326 16908 45360 16942
rect 45326 16840 45360 16874
rect 42478 16772 42512 16806
rect 42658 16762 42705 16796
rect 42741 16762 42775 16796
rect 42811 16762 42858 16796
rect 42916 16762 42963 16796
rect 42999 16762 43033 16796
rect 43069 16762 43116 16796
rect 43174 16762 43221 16796
rect 43257 16762 43291 16796
rect 43327 16762 43374 16796
rect 43432 16762 43479 16796
rect 43515 16762 43549 16796
rect 43585 16762 43632 16796
rect 43690 16762 43737 16796
rect 43773 16762 43807 16796
rect 43843 16762 43890 16796
rect 43948 16762 43995 16796
rect 44031 16762 44065 16796
rect 44101 16762 44148 16796
rect 44206 16762 44253 16796
rect 44289 16762 44323 16796
rect 44359 16762 44406 16796
rect 44464 16762 44511 16796
rect 44547 16762 44581 16796
rect 44617 16762 44664 16796
rect 44722 16762 44769 16796
rect 44805 16762 44839 16796
rect 44875 16762 44922 16796
rect 44980 16762 45027 16796
rect 45063 16762 45097 16796
rect 45133 16762 45180 16796
rect 45326 16772 45360 16806
rect 42478 16658 42512 16738
rect 45326 16658 45360 16738
rect 42478 16624 42576 16658
rect 42610 16624 42644 16658
rect 42678 16624 42712 16658
rect 42746 16624 42780 16658
rect 42814 16624 42848 16658
rect 42882 16624 42916 16658
rect 42950 16624 42984 16658
rect 43018 16624 43052 16658
rect 43086 16624 43120 16658
rect 43154 16624 43188 16658
rect 43222 16624 43256 16658
rect 43290 16624 43324 16658
rect 43358 16624 43392 16658
rect 43426 16624 43460 16658
rect 43494 16624 43528 16658
rect 43562 16624 43596 16658
rect 43630 16624 43664 16658
rect 43698 16624 43732 16658
rect 43766 16624 43800 16658
rect 43834 16624 43868 16658
rect 43902 16624 43936 16658
rect 43970 16624 44004 16658
rect 44038 16624 44072 16658
rect 44106 16624 44140 16658
rect 44174 16624 44208 16658
rect 44242 16624 44276 16658
rect 44310 16624 44344 16658
rect 44378 16624 44412 16658
rect 44446 16624 44480 16658
rect 44514 16624 44548 16658
rect 44582 16624 44616 16658
rect 44650 16624 44684 16658
rect 44718 16624 44752 16658
rect 44786 16624 44820 16658
rect 44854 16624 44888 16658
rect 44922 16624 44956 16658
rect 44990 16624 45024 16658
rect 45058 16624 45092 16658
rect 45126 16624 45160 16658
rect 45194 16624 45228 16658
rect 45262 16624 45360 16658
rect 27650 16578 27684 16612
rect 24460 16510 24494 16544
rect 24460 16442 24494 16476
rect 24460 16374 24494 16408
rect 24460 16306 24494 16340
rect 27650 16510 27684 16544
rect 27650 16442 27684 16476
rect 27650 16374 27684 16408
rect 27650 16306 27684 16340
rect 24460 16238 24494 16272
rect 27650 16238 27684 16272
rect 24460 16170 24494 16204
rect 24460 16102 24494 16136
rect 24460 16034 24494 16068
rect 24460 15966 24494 16000
rect 27650 16170 27684 16204
rect 27650 16102 27684 16136
rect 27650 16034 27684 16068
rect 24460 15898 24494 15932
rect 27650 15966 27684 16000
rect 10297 14996 22482 15011
rect 10297 14986 17059 14996
rect 10297 14952 12964 14986
rect 12998 14952 13032 14986
rect 13066 14952 13100 14986
rect 13134 14952 13168 14986
rect 13202 14952 13236 14986
rect 13270 14952 13304 14986
rect 13338 14952 13372 14986
rect 13406 14952 13440 14986
rect 13474 14952 13508 14986
rect 13542 14952 13576 14986
rect 13610 14952 13644 14986
rect 13678 14952 13712 14986
rect 13746 14952 13780 14986
rect 13814 14952 13848 14986
rect 13882 14952 13916 14986
rect 13950 14952 13984 14986
rect 14018 14952 14052 14986
rect 14086 14952 14120 14986
rect 14154 14952 14188 14986
rect 14222 14952 14256 14986
rect 14290 14952 14324 14986
rect 14358 14952 14392 14986
rect 14426 14952 14460 14986
rect 14494 14952 14528 14986
rect 14562 14952 14596 14986
rect 14630 14952 14664 14986
rect 14698 14952 14732 14986
rect 14766 14952 14800 14986
rect 14834 14952 14868 14986
rect 14902 14952 14936 14986
rect 14970 14952 15004 14986
rect 15038 14952 15072 14986
rect 15106 14952 15140 14986
rect 15174 14952 15549 14986
rect 15583 14952 15617 14986
rect 15651 14952 15685 14986
rect 15719 14952 15753 14986
rect 15787 14952 15821 14986
rect 15855 14952 15889 14986
rect 15923 14952 15957 14986
rect 15991 14952 16025 14986
rect 16059 14952 16093 14986
rect 16127 14952 16161 14986
rect 16195 14952 16229 14986
rect 16263 14952 16297 14986
rect 16331 14952 16365 14986
rect 16399 14952 16433 14986
rect 16467 14952 16501 14986
rect 16535 14952 16569 14986
rect 16603 14952 16637 14986
rect 16671 14962 17059 14986
rect 17093 14962 17127 14996
rect 17161 14962 17195 14996
rect 17229 14962 17263 14996
rect 17297 14962 17331 14996
rect 17365 14962 17399 14996
rect 17433 14962 17467 14996
rect 17501 14962 17535 14996
rect 17569 14962 17603 14996
rect 17637 14962 17671 14996
rect 17705 14962 17739 14996
rect 17773 14962 17807 14996
rect 17841 14962 17875 14996
rect 17909 14962 17943 14996
rect 17977 14962 18011 14996
rect 18045 14962 18079 14996
rect 18113 14962 18147 14996
rect 18181 14980 22482 14996
rect 18181 14962 18523 14980
rect 16671 14952 18523 14962
rect -4010 14846 -3976 14880
rect -4010 14778 -3976 14812
rect -4010 14710 -3976 14744
rect -4010 14642 -3976 14676
rect -4010 14574 -3976 14608
rect -4010 14506 -3976 14540
rect -3714 14846 -3680 14880
rect -3714 14778 -3680 14812
rect -3714 14710 -3680 14744
rect -3714 14642 -3680 14676
rect -3714 14574 -3680 14608
rect -3714 14506 -3680 14540
rect -4010 14438 -3976 14472
rect -4010 14370 -3976 14404
rect -4010 14302 -3976 14336
rect -4010 14234 -3976 14268
rect -4010 14166 -3976 14200
rect -4010 14098 -3976 14132
rect -4010 14030 -3976 14064
rect -4010 13962 -3976 13996
rect -4010 13894 -3976 13928
rect -4010 13826 -3976 13860
rect -4010 13758 -3976 13792
rect -4010 13690 -3976 13724
rect -4010 13622 -3976 13656
rect -4010 13554 -3976 13588
rect -4010 13486 -3976 13520
rect -4010 13418 -3976 13452
rect -4010 13350 -3976 13384
rect -4010 13282 -3976 13316
rect -4010 13214 -3976 13248
rect -4010 13146 -3976 13180
rect -4010 13078 -3976 13112
rect -4010 13010 -3976 13044
rect -4010 12942 -3976 12976
rect -4010 12874 -3976 12908
rect -3714 14438 -3680 14472
rect -3714 14370 -3680 14404
rect -3714 14302 -3680 14336
rect -3714 14234 -3680 14268
rect -3714 14166 -3680 14200
rect -3714 14098 -3680 14132
rect -3714 14030 -3680 14064
rect -3714 13962 -3680 13996
rect -3714 13894 -3680 13928
rect -3714 13826 -3680 13860
rect -3714 13758 -3680 13792
rect -3714 13690 -3680 13724
rect -3714 13622 -3680 13656
rect -3714 13554 -3680 13588
rect -3714 13486 -3680 13520
rect -3714 13418 -3680 13452
rect -3714 13350 -3680 13384
rect -3714 13282 -3680 13316
rect -3714 13214 -3680 13248
rect -3714 13146 -3680 13180
rect -3714 13078 -3680 13112
rect -3714 13010 -3680 13044
rect -3714 12942 -3680 12976
rect -3714 12874 -3680 12908
rect -4010 12806 -3976 12840
rect -4010 12738 -3976 12772
rect -4010 12670 -3976 12704
rect -4010 12602 -3976 12636
rect -4010 12534 -3976 12568
rect -4010 12466 -3976 12500
rect -3714 12806 -3680 12840
rect -3714 12738 -3680 12772
rect -3714 12670 -3680 12704
rect -3714 12602 -3680 12636
rect -3714 12534 -3680 12568
rect -3714 12466 -3680 12500
rect -4010 12355 -3976 12432
rect -3714 12355 -3680 12432
rect 12860 14882 12894 14952
rect 15244 14882 15278 14952
rect 13942 14848 14202 14870
rect 12860 14814 12894 14848
rect 13040 14814 13081 14848
rect 13125 14814 13149 14848
rect 13197 14814 13217 14848
rect 13269 14814 13285 14848
rect 13341 14814 13353 14848
rect 13413 14814 13421 14848
rect 13485 14814 13489 14848
rect 13591 14814 13595 14848
rect 13659 14814 13667 14848
rect 13727 14814 13739 14848
rect 13795 14814 13811 14848
rect 13863 14814 13883 14848
rect 13931 14814 13955 14848
rect 13999 14814 14139 14848
rect 14183 14814 14207 14848
rect 14255 14814 14275 14848
rect 14327 14814 14343 14848
rect 14399 14814 14411 14848
rect 14471 14814 14479 14848
rect 14543 14814 14547 14848
rect 14649 14814 14653 14848
rect 14717 14814 14725 14848
rect 14785 14814 14797 14848
rect 14853 14814 14869 14848
rect 14921 14814 14941 14848
rect 14989 14814 15013 14848
rect 15057 14814 15098 14848
rect 15244 14814 15278 14848
rect 13942 14810 14202 14814
rect 12860 14746 12894 14780
rect 12860 14678 12894 14712
rect 12860 14610 12894 14644
rect 12860 14542 12894 14576
rect 12860 14474 12894 14508
rect 12860 14406 12894 14440
rect 12860 14338 12894 14372
rect 12860 14270 12894 14304
rect 12860 14202 12894 14236
rect 12860 14134 12894 14168
rect 12860 14066 12894 14100
rect 12860 13998 12894 14032
rect 12860 13930 12894 13964
rect 12860 13862 12894 13896
rect 12860 13794 12894 13828
rect 12860 13726 12894 13760
rect 12860 13658 12894 13692
rect 12860 13590 12894 13624
rect 12860 13522 12894 13556
rect 12860 13454 12894 13488
rect 12860 13386 12894 13420
rect 12860 13318 12894 13352
rect 12860 13250 12894 13284
rect 12860 13182 12894 13216
rect 12860 13114 12894 13148
rect 12860 13046 12894 13080
rect 12860 12978 12894 13012
rect 12860 12910 12894 12944
rect 12860 12842 12894 12876
rect 12860 12774 12894 12808
rect 12860 12706 12894 12740
rect 12860 12638 12894 12672
rect 12860 12570 12894 12604
rect 12860 12502 12894 12536
rect 12860 12434 12894 12468
rect 12860 12366 12894 12400
rect -4545 12310 -4503 12344
rect -4469 12310 -4427 12344
rect -4082 12345 -3626 12355
rect -4082 12326 -3896 12345
rect -4545 12278 -4427 12310
rect -4086 12311 -3896 12326
rect -3862 12311 -3828 12345
rect -3794 12311 -3626 12345
rect -7888 12236 -4421 12278
rect -7888 12202 -7570 12236
rect -7536 12202 -7502 12236
rect -7468 12202 -7434 12236
rect -7400 12202 -7366 12236
rect -7332 12202 -7298 12236
rect -7264 12202 -7230 12236
rect -7196 12202 -7162 12236
rect -7128 12202 -7094 12236
rect -7060 12202 -7026 12236
rect -6992 12202 -6958 12236
rect -6924 12202 -6890 12236
rect -6856 12202 -6822 12236
rect -6788 12202 -6754 12236
rect -6720 12202 -6686 12236
rect -6652 12202 -6618 12236
rect -6584 12202 -6550 12236
rect -6516 12202 -6482 12236
rect -6448 12202 -6414 12236
rect -6380 12202 -6346 12236
rect -6312 12202 -6278 12236
rect -6244 12202 -6210 12236
rect -6176 12202 -6142 12236
rect -6108 12202 -6074 12236
rect -6040 12202 -6006 12236
rect -5972 12202 -5938 12236
rect -5904 12202 -5870 12236
rect -5836 12202 -5802 12236
rect -5768 12202 -5734 12236
rect -5700 12202 -5666 12236
rect -5632 12202 -5598 12236
rect -5564 12202 -5530 12236
rect -5496 12202 -5462 12236
rect -5428 12202 -5394 12236
rect -5360 12202 -5326 12236
rect -5292 12202 -5258 12236
rect -5224 12202 -5190 12236
rect -5156 12202 -5122 12236
rect -5088 12202 -5054 12236
rect -5020 12202 -4986 12236
rect -4952 12202 -4918 12236
rect -4884 12202 -4850 12236
rect -4816 12202 -4782 12236
rect -4748 12202 -4714 12236
rect -4680 12202 -4646 12236
rect -4612 12202 -4421 12236
rect -7888 12184 -4421 12202
rect -4086 12184 -3626 12311
rect -7888 12163 -3626 12184
rect -7906 11913 -3626 12163
rect -7906 11595 -4406 11913
rect -4082 11911 -3626 11913
rect 12860 12298 12894 12332
rect 12860 12230 12894 12264
rect 12860 12162 12894 12196
rect 12860 12094 12894 12128
rect 12860 12026 12894 12060
rect 12860 11958 12894 11992
rect 12860 11890 12894 11924
rect 12860 11822 12894 11856
rect 12860 11754 12894 11788
rect 12994 14746 13028 14771
rect 12994 14678 13028 14690
rect 12994 14610 13028 14618
rect 12994 14542 13028 14546
rect 12994 14436 13028 14440
rect 12994 14364 13028 14372
rect 12994 14292 13028 14304
rect 12994 14220 13028 14236
rect 12994 14148 13028 14168
rect 12994 14076 13028 14100
rect 12994 14004 13028 14032
rect 12994 13932 13028 13964
rect 12994 13862 13028 13896
rect 12994 13794 13028 13826
rect 12994 13726 13028 13754
rect 12994 13658 13028 13682
rect 12994 13590 13028 13610
rect 12994 13522 13028 13538
rect 12994 13454 13028 13466
rect 12994 13386 13028 13394
rect 12994 13318 13028 13322
rect 12994 13212 13028 13216
rect 12994 13140 13028 13148
rect 12994 13068 13028 13080
rect 12994 12996 13028 13012
rect 12994 12924 13028 12944
rect 12994 12852 13028 12876
rect 12994 12780 13028 12808
rect 12994 12708 13028 12740
rect 12994 12638 13028 12672
rect 12994 12570 13028 12602
rect 12994 12502 13028 12530
rect 12994 12434 13028 12458
rect 12994 12366 13028 12386
rect 12994 12298 13028 12314
rect 12994 12230 13028 12242
rect 12994 12162 13028 12170
rect 12994 12094 13028 12098
rect 12994 11988 13028 11992
rect 12994 11916 13028 11924
rect 12994 11844 13028 11856
rect 12994 11763 13028 11788
rect 14052 14746 14086 14771
rect 14052 14678 14086 14690
rect 14052 14610 14086 14618
rect 14052 14542 14086 14546
rect 14052 14436 14086 14440
rect 14052 14364 14086 14372
rect 14052 14292 14086 14304
rect 14052 14220 14086 14236
rect 14052 14148 14086 14168
rect 14052 14076 14086 14100
rect 14052 14004 14086 14032
rect 14052 13932 14086 13964
rect 14052 13862 14086 13896
rect 14052 13794 14086 13826
rect 14052 13726 14086 13754
rect 14052 13658 14086 13682
rect 14052 13590 14086 13610
rect 14052 13522 14086 13538
rect 14052 13454 14086 13466
rect 14052 13386 14086 13394
rect 14052 13318 14086 13322
rect 14052 13212 14086 13216
rect 14052 13140 14086 13148
rect 14052 13068 14086 13080
rect 14052 12996 14086 13012
rect 14052 12924 14086 12944
rect 14052 12852 14086 12876
rect 14052 12780 14086 12808
rect 14052 12708 14086 12740
rect 14052 12638 14086 12672
rect 14052 12570 14086 12602
rect 14052 12502 14086 12530
rect 14052 12434 14086 12458
rect 14052 12366 14086 12386
rect 14052 12298 14086 12314
rect 14052 12230 14086 12242
rect 14052 12162 14086 12170
rect 14052 12094 14086 12098
rect 14052 11988 14086 11992
rect 14052 11916 14086 11924
rect 14052 11844 14086 11856
rect 14052 11763 14086 11788
rect 15110 14746 15144 14771
rect 15110 14678 15144 14690
rect 15110 14610 15144 14618
rect 15110 14542 15144 14546
rect 15110 14436 15144 14440
rect 15110 14364 15144 14372
rect 15110 14292 15144 14304
rect 15110 14220 15144 14236
rect 15110 14148 15144 14168
rect 15110 14076 15144 14100
rect 15110 14004 15144 14032
rect 15110 13932 15144 13964
rect 15110 13862 15144 13896
rect 15110 13794 15144 13826
rect 15110 13726 15144 13754
rect 15110 13658 15144 13682
rect 15110 13590 15144 13610
rect 15110 13522 15144 13538
rect 15110 13454 15144 13466
rect 15110 13386 15144 13394
rect 15110 13318 15144 13322
rect 15110 13212 15144 13216
rect 15110 13140 15144 13148
rect 15110 13068 15144 13080
rect 15110 12996 15144 13012
rect 15110 12924 15144 12944
rect 15110 12852 15144 12876
rect 15110 12780 15144 12808
rect 15110 12708 15144 12740
rect 15110 12638 15144 12672
rect 15110 12570 15144 12602
rect 15110 12502 15144 12530
rect 15110 12434 15144 12458
rect 15110 12366 15144 12386
rect 15110 12298 15144 12314
rect 15110 12230 15144 12242
rect 15110 12162 15144 12170
rect 15110 12094 15144 12098
rect 15110 11988 15144 11992
rect 15110 11916 15144 11924
rect 15110 11844 15144 11856
rect 15110 11763 15144 11788
rect 15244 14746 15278 14780
rect 15244 14678 15278 14712
rect 15244 14610 15278 14644
rect 15244 14542 15278 14576
rect 15244 14474 15278 14508
rect 15244 14406 15278 14440
rect 15244 14338 15278 14372
rect 15244 14270 15278 14304
rect 15244 14202 15278 14236
rect 15244 14134 15278 14168
rect 15244 14066 15278 14100
rect 15244 13998 15278 14032
rect 15244 13930 15278 13964
rect 15244 13862 15278 13896
rect 15244 13794 15278 13828
rect 15244 13726 15278 13760
rect 15244 13658 15278 13692
rect 15244 13590 15278 13624
rect 15244 13522 15278 13556
rect 15244 13454 15278 13488
rect 15244 13386 15278 13420
rect 15244 13318 15278 13352
rect 15244 13250 15278 13284
rect 15244 13182 15278 13216
rect 15244 13114 15278 13148
rect 15244 13046 15278 13080
rect 15244 12978 15278 13012
rect 15244 12910 15278 12944
rect 15244 12842 15278 12876
rect 15244 12774 15278 12808
rect 15244 12706 15278 12740
rect 15244 12638 15278 12672
rect 15244 12570 15278 12604
rect 15244 12502 15278 12536
rect 15244 12434 15278 12468
rect 15244 12366 15278 12400
rect 15244 12298 15278 12332
rect 15244 12230 15278 12264
rect 15244 12162 15278 12196
rect 15244 12094 15278 12128
rect 15244 12026 15278 12060
rect 15244 11958 15278 11992
rect 15244 11890 15278 11924
rect 15244 11822 15278 11856
rect 15244 11754 15278 11788
rect 12860 11686 12894 11720
rect 13040 11686 13081 11720
rect 13125 11686 13149 11720
rect 13197 11686 13217 11720
rect 13269 11686 13285 11720
rect 13341 11686 13353 11720
rect 13413 11686 13421 11720
rect 13485 11686 13489 11720
rect 13591 11686 13595 11720
rect 13659 11686 13667 11720
rect 13727 11686 13739 11720
rect 13795 11686 13811 11720
rect 13863 11686 13883 11720
rect 13931 11686 13955 11720
rect 13999 11686 14139 11720
rect 14183 11686 14207 11720
rect 14255 11686 14275 11720
rect 14327 11686 14343 11720
rect 14399 11686 14411 11720
rect 14471 11686 14479 11720
rect 14543 11686 14547 11720
rect 14649 11686 14653 11720
rect 14717 11686 14725 11720
rect 14785 11686 14797 11720
rect 14853 11686 14869 11720
rect 14921 11686 14941 11720
rect 14989 11686 15013 11720
rect 15057 11686 15098 11720
rect 15244 11686 15278 11720
rect 13972 11670 14192 11686
rect -9108 11565 -3289 11595
rect -9108 11531 -8832 11565
rect -8798 11531 -8764 11565
rect -8730 11531 -8696 11565
rect -8662 11531 -8628 11565
rect -8594 11531 -8560 11565
rect -8526 11531 -8492 11565
rect -8458 11531 -8424 11565
rect -8390 11531 -8356 11565
rect -8322 11531 -8288 11565
rect -8254 11531 -8220 11565
rect -8186 11531 -8152 11565
rect -8118 11531 -8084 11565
rect -8050 11531 -8016 11565
rect -7982 11531 -7948 11565
rect -7914 11531 -7880 11565
rect -7846 11531 -7812 11565
rect -7778 11531 -7744 11565
rect -7710 11531 -7676 11565
rect -7642 11531 -7608 11565
rect -7574 11531 -7540 11565
rect -7506 11531 -7472 11565
rect -7438 11531 -7404 11565
rect -7370 11531 -7336 11565
rect -7302 11531 -7268 11565
rect -7234 11531 -7200 11565
rect -7166 11531 -7132 11565
rect -7098 11531 -7064 11565
rect -7030 11531 -6996 11565
rect -6962 11531 -6928 11565
rect -6894 11531 -6860 11565
rect -6826 11531 -6792 11565
rect -6758 11531 -6724 11565
rect -6690 11531 -6656 11565
rect -6622 11531 -6588 11565
rect -6554 11531 -6520 11565
rect -6486 11531 -6452 11565
rect -6418 11531 -6384 11565
rect -6350 11531 -6316 11565
rect -6282 11531 -6248 11565
rect -6214 11531 -6180 11565
rect -6146 11531 -6112 11565
rect -6078 11531 -6044 11565
rect -6010 11531 -5976 11565
rect -5942 11531 -5908 11565
rect -5874 11531 -5840 11565
rect -5806 11531 -5772 11565
rect -5738 11531 -5704 11565
rect -5670 11531 -5636 11565
rect -5602 11531 -5568 11565
rect -5534 11531 -5500 11565
rect -5466 11531 -5432 11565
rect -5398 11531 -5364 11565
rect -5330 11531 -5296 11565
rect -5262 11531 -5228 11565
rect -5194 11531 -5160 11565
rect -5126 11531 -5092 11565
rect -5058 11531 -5024 11565
rect -4990 11531 -4956 11565
rect -4922 11531 -4888 11565
rect -4854 11531 -4820 11565
rect -4786 11531 -4752 11565
rect -4718 11531 -4684 11565
rect -4650 11531 -4616 11565
rect -4582 11531 -4548 11565
rect -4514 11531 -4480 11565
rect -4446 11531 -4412 11565
rect -4378 11531 -4344 11565
rect -4310 11531 -4276 11565
rect -4242 11531 -4208 11565
rect -4174 11531 -4140 11565
rect -4106 11531 -4072 11565
rect -4038 11531 -4004 11565
rect -3970 11531 -3936 11565
rect -3902 11531 -3868 11565
rect -3834 11531 -3800 11565
rect -3766 11531 -3732 11565
rect -3698 11531 -3664 11565
rect -3630 11531 -3596 11565
rect -3562 11531 -3289 11565
rect 12860 11582 12894 11652
rect 15244 11582 15278 11652
rect 12860 11548 12964 11582
rect 12998 11548 13032 11582
rect 13066 11548 13100 11582
rect 13134 11548 13168 11582
rect 13202 11548 13236 11582
rect 13270 11548 13304 11582
rect 13338 11548 13372 11582
rect 13406 11548 13440 11582
rect 13474 11548 13508 11582
rect 13542 11548 13576 11582
rect 13610 11548 13644 11582
rect 13678 11548 13712 11582
rect 13746 11548 13780 11582
rect 13814 11548 13848 11582
rect 13882 11548 13916 11582
rect 13950 11548 13984 11582
rect 14018 11548 14052 11582
rect 14086 11548 14120 11582
rect 14154 11548 14188 11582
rect 14222 11548 14256 11582
rect 14290 11548 14324 11582
rect 14358 11548 14392 11582
rect 14426 11548 14460 11582
rect 14494 11548 14528 11582
rect 14562 11548 14596 11582
rect 14630 11548 14664 11582
rect 14698 11548 14732 11582
rect 14766 11548 14800 11582
rect 14834 11548 14868 11582
rect 14902 11548 14936 11582
rect 14970 11548 15004 11582
rect 15038 11548 15072 11582
rect 15106 11548 15140 11582
rect 15174 11548 15278 11582
rect 15430 14882 15464 14952
rect 16756 14882 16790 14952
rect 15430 14814 15464 14848
rect 15610 14814 15651 14848
rect 15695 14814 15719 14848
rect 15767 14814 15787 14848
rect 15839 14814 15855 14848
rect 15911 14814 15923 14848
rect 15983 14814 15991 14848
rect 16055 14814 16059 14848
rect 16161 14814 16165 14848
rect 16229 14814 16237 14848
rect 16297 14814 16309 14848
rect 16365 14814 16381 14848
rect 16433 14814 16453 14848
rect 16501 14814 16525 14848
rect 16569 14814 16610 14848
rect 16756 14814 16790 14848
rect 15430 14746 15464 14780
rect 15430 14678 15464 14712
rect 15430 14610 15464 14644
rect 15430 14542 15464 14576
rect 15430 14474 15464 14508
rect 15430 14406 15464 14440
rect 15430 14338 15464 14372
rect 15430 14270 15464 14304
rect 15430 14202 15464 14236
rect 15430 14134 15464 14168
rect 15430 14066 15464 14100
rect 15430 13998 15464 14032
rect 15430 13930 15464 13964
rect 15430 13862 15464 13896
rect 15430 13794 15464 13828
rect 15430 13726 15464 13760
rect 15430 13658 15464 13692
rect 15430 13590 15464 13624
rect 15430 13522 15464 13556
rect 15430 13454 15464 13488
rect 15430 13386 15464 13420
rect 15430 13318 15464 13352
rect 15430 13250 15464 13284
rect 15430 13182 15464 13216
rect 15430 13114 15464 13148
rect 15430 13046 15464 13080
rect 15430 12978 15464 13012
rect 15430 12910 15464 12944
rect 15430 12842 15464 12876
rect 15430 12774 15464 12808
rect 15430 12706 15464 12740
rect 15430 12638 15464 12672
rect 15430 12570 15464 12604
rect 15430 12502 15464 12536
rect 15430 12434 15464 12468
rect 15430 12366 15464 12400
rect 15430 12298 15464 12332
rect 15430 12230 15464 12264
rect 15430 12162 15464 12196
rect 15430 12094 15464 12128
rect 15430 12026 15464 12060
rect 15430 11958 15464 11992
rect 15430 11890 15464 11924
rect 15430 11822 15464 11856
rect 15430 11754 15464 11788
rect 15564 14746 15598 14771
rect 16622 14746 16656 14771
rect 15564 14678 15598 14690
rect 15564 14610 15598 14618
rect 15564 14542 15598 14546
rect 15564 14436 15598 14440
rect 16612 14690 16622 14710
rect 16756 14746 16790 14780
rect 16756 14710 16790 14712
rect 16656 14690 16790 14710
rect 16612 14678 16790 14690
rect 16612 14618 16622 14678
rect 16656 14644 16756 14678
rect 16656 14618 16790 14644
rect 16612 14610 16790 14618
rect 16612 14546 16622 14610
rect 16656 14576 16756 14610
rect 16656 14546 16790 14576
rect 16612 14542 16790 14546
rect 16612 14440 16622 14542
rect 16656 14508 16756 14542
rect 16656 14474 16790 14508
rect 16656 14440 16756 14474
rect 16612 14436 16790 14440
rect 16612 14420 16622 14436
rect 15564 14364 15598 14372
rect 15564 14292 15598 14304
rect 15564 14220 15598 14236
rect 15564 14148 15598 14168
rect 15564 14076 15598 14100
rect 15564 14004 15598 14032
rect 15564 13932 15598 13964
rect 15564 13862 15598 13896
rect 15564 13794 15598 13826
rect 15564 13726 15598 13754
rect 15564 13658 15598 13682
rect 15564 13590 15598 13610
rect 15564 13522 15598 13538
rect 15564 13454 15598 13466
rect 15564 13386 15598 13394
rect 15564 13318 15598 13322
rect 15564 13212 15598 13216
rect 15564 13140 15598 13148
rect 15564 13068 15598 13080
rect 15564 12996 15598 13012
rect 15564 12924 15598 12944
rect 15564 12852 15598 12876
rect 15564 12780 15598 12808
rect 15564 12708 15598 12740
rect 15564 12638 15598 12672
rect 15564 12570 15598 12602
rect 15564 12502 15598 12530
rect 15564 12434 15598 12458
rect 15564 12366 15598 12386
rect 15564 12298 15598 12314
rect 15564 12230 15598 12242
rect 15564 12162 15598 12170
rect 15564 12094 15598 12098
rect 15564 11988 15598 11992
rect 15564 11916 15598 11924
rect 15564 11844 15598 11856
rect 15564 11763 15598 11788
rect 16656 14420 16790 14436
rect 16622 14364 16656 14372
rect 16622 14292 16656 14304
rect 16622 14220 16656 14236
rect 16622 14148 16656 14168
rect 16622 14076 16656 14100
rect 16622 14004 16656 14032
rect 16622 13932 16656 13964
rect 16622 13862 16656 13896
rect 16622 13794 16656 13826
rect 16622 13726 16656 13754
rect 16622 13658 16656 13682
rect 16622 13590 16656 13610
rect 16622 13522 16656 13538
rect 16622 13454 16656 13466
rect 16622 13386 16656 13394
rect 16622 13318 16656 13322
rect 16622 13212 16656 13216
rect 16622 13140 16656 13148
rect 16622 13068 16656 13080
rect 16622 12996 16656 13012
rect 16622 12924 16656 12944
rect 16622 12852 16656 12876
rect 16622 12780 16656 12808
rect 16622 12708 16656 12740
rect 16622 12638 16656 12672
rect 16622 12570 16656 12602
rect 16622 12502 16656 12530
rect 16622 12434 16656 12458
rect 16622 12366 16656 12386
rect 16622 12298 16656 12314
rect 16622 12230 16656 12242
rect 16622 12162 16656 12170
rect 16622 12094 16656 12098
rect 16622 11988 16656 11992
rect 16622 11916 16656 11924
rect 16622 11844 16656 11856
rect 16622 11763 16656 11788
rect 16756 14406 16790 14420
rect 16756 14338 16790 14372
rect 16756 14270 16790 14304
rect 16756 14202 16790 14236
rect 16756 14134 16790 14168
rect 16756 14066 16790 14100
rect 16756 13998 16790 14032
rect 16756 13930 16790 13964
rect 16756 13862 16790 13896
rect 16756 13794 16790 13828
rect 16756 13726 16790 13760
rect 16756 13658 16790 13692
rect 16756 13590 16790 13624
rect 16756 13522 16790 13556
rect 16756 13454 16790 13488
rect 16756 13386 16790 13420
rect 16756 13318 16790 13352
rect 16756 13250 16790 13284
rect 16756 13182 16790 13216
rect 16756 13114 16790 13148
rect 16756 13046 16790 13080
rect 16756 12978 16790 13012
rect 16756 12910 16790 12944
rect 16756 12842 16790 12876
rect 16756 12774 16790 12808
rect 16756 12706 16790 12740
rect 16756 12638 16790 12672
rect 16756 12570 16790 12604
rect 16756 12502 16790 12536
rect 16756 12434 16790 12468
rect 16756 12366 16790 12400
rect 16756 12298 16790 12332
rect 16756 12230 16790 12264
rect 16756 12162 16790 12196
rect 16756 12094 16790 12128
rect 16756 12026 16790 12060
rect 16756 11958 16790 11992
rect 16756 11890 16790 11924
rect 16756 11822 16790 11856
rect 16756 11754 16790 11788
rect 15430 11686 15464 11720
rect 15610 11686 15651 11720
rect 15695 11686 15719 11720
rect 15767 11686 15787 11720
rect 15839 11686 15855 11720
rect 15911 11686 15923 11720
rect 15983 11686 15991 11720
rect 16055 11686 16059 11720
rect 16161 11686 16165 11720
rect 16229 11686 16237 11720
rect 16297 11686 16309 11720
rect 16365 11686 16381 11720
rect 16433 11686 16453 11720
rect 16501 11686 16525 11720
rect 16569 11686 16610 11720
rect 16756 11686 16790 11720
rect 15430 11582 15464 11652
rect 16756 11582 16790 11652
rect 15430 11548 15549 11582
rect 15583 11548 15617 11582
rect 15651 11548 15685 11582
rect 15719 11548 15753 11582
rect 15787 11548 15821 11582
rect 15855 11548 15889 11582
rect 15923 11548 15957 11582
rect 15991 11548 16025 11582
rect 16059 11548 16093 11582
rect 16127 11548 16161 11582
rect 16195 11548 16229 11582
rect 16263 11548 16297 11582
rect 16331 11548 16365 11582
rect 16399 11548 16433 11582
rect 16467 11548 16501 11582
rect 16535 11548 16569 11582
rect 16603 11548 16637 11582
rect 16671 11548 16790 11582
rect 16940 14892 16974 14952
rect 18266 14892 18300 14952
rect 16940 14824 16974 14858
rect 17120 14824 17161 14858
rect 17205 14824 17229 14858
rect 17277 14824 17297 14858
rect 17349 14824 17365 14858
rect 17421 14824 17433 14858
rect 17493 14824 17501 14858
rect 17565 14824 17569 14858
rect 17671 14824 17675 14858
rect 17739 14824 17747 14858
rect 17807 14824 17819 14858
rect 17875 14824 17891 14858
rect 17943 14824 17963 14858
rect 18011 14824 18035 14858
rect 18079 14824 18120 14858
rect 18266 14824 18300 14858
rect 16940 14756 16974 14790
rect 16940 14688 16974 14722
rect 16940 14620 16974 14654
rect 16940 14552 16974 14586
rect 16940 14484 16974 14518
rect 16940 14416 16974 14450
rect 16940 14348 16974 14382
rect 16940 14280 16974 14314
rect 16940 14212 16974 14246
rect 16940 14144 16974 14178
rect 16940 14076 16974 14110
rect 16940 14008 16974 14042
rect 16940 13940 16974 13974
rect 16940 13872 16974 13906
rect 16940 13804 16974 13838
rect 16940 13736 16974 13770
rect 16940 13668 16974 13702
rect 16940 13600 16974 13634
rect 16940 13532 16974 13566
rect 16940 13464 16974 13498
rect 16940 13396 16974 13430
rect 16940 13328 16974 13362
rect 16940 13260 16974 13294
rect 16940 13192 16974 13226
rect 16940 13124 16974 13158
rect 16940 13056 16974 13090
rect 16940 12988 16974 13022
rect 16940 12920 16974 12954
rect 16940 12852 16974 12886
rect 16940 12784 16974 12818
rect 16940 12716 16974 12750
rect 16940 12648 16974 12682
rect 16940 12580 16974 12614
rect 16940 12512 16974 12546
rect 16940 12444 16974 12478
rect 16940 12376 16974 12410
rect 16940 12308 16974 12342
rect 16940 12240 16974 12274
rect 16940 12172 16974 12206
rect 16940 12104 16974 12138
rect 16940 12036 16974 12070
rect 16940 11968 16974 12002
rect 16940 11900 16974 11934
rect 16940 11832 16974 11866
rect 16940 11764 16974 11798
rect 17074 14756 17108 14781
rect 18132 14770 18166 14781
rect 18266 14770 18300 14790
rect 18404 14946 18523 14952
rect 18557 14946 18591 14980
rect 18625 14946 18659 14980
rect 18693 14946 18727 14980
rect 18761 14946 18795 14980
rect 18829 14946 18863 14980
rect 18897 14946 18931 14980
rect 18965 14946 18999 14980
rect 19033 14946 19067 14980
rect 19101 14946 19135 14980
rect 19169 14946 19203 14980
rect 19237 14946 19271 14980
rect 19305 14946 19339 14980
rect 19373 14946 19407 14980
rect 19441 14946 19475 14980
rect 19509 14946 19543 14980
rect 19577 14946 19611 14980
rect 19645 14952 22482 14980
rect 19645 14946 19764 14952
rect 18404 14876 18438 14946
rect 19730 14876 19764 14946
rect 18404 14808 18438 14842
rect 18584 14808 18625 14842
rect 18669 14808 18693 14842
rect 18741 14808 18761 14842
rect 18813 14808 18829 14842
rect 18885 14808 18897 14842
rect 18957 14808 18965 14842
rect 19029 14808 19033 14842
rect 19135 14808 19139 14842
rect 19203 14808 19211 14842
rect 19271 14808 19283 14842
rect 19339 14808 19355 14842
rect 19407 14808 19427 14842
rect 19475 14808 19499 14842
rect 19543 14808 19584 14842
rect 19730 14808 19764 14842
rect 17074 14688 17108 14700
rect 17074 14620 17108 14628
rect 17074 14552 17108 14556
rect 17074 14446 17108 14450
rect 17074 14374 17108 14382
rect 17074 14302 17108 14314
rect 18122 14756 18302 14770
rect 18122 14700 18132 14756
rect 18166 14722 18266 14756
rect 18300 14722 18302 14756
rect 18166 14700 18302 14722
rect 18122 14688 18302 14700
rect 18122 14628 18132 14688
rect 18166 14654 18266 14688
rect 18300 14654 18302 14688
rect 18166 14628 18302 14654
rect 18122 14620 18302 14628
rect 18122 14556 18132 14620
rect 18166 14586 18266 14620
rect 18300 14586 18302 14620
rect 18166 14556 18302 14586
rect 18122 14552 18302 14556
rect 18122 14450 18132 14552
rect 18166 14518 18266 14552
rect 18300 14518 18302 14552
rect 18166 14484 18302 14518
rect 18166 14450 18266 14484
rect 18300 14450 18302 14484
rect 18122 14446 18302 14450
rect 18122 14382 18132 14446
rect 18166 14416 18302 14446
rect 18166 14382 18266 14416
rect 18300 14382 18302 14416
rect 18122 14374 18302 14382
rect 18122 14314 18132 14374
rect 18166 14348 18302 14374
rect 18166 14314 18266 14348
rect 18300 14314 18302 14348
rect 18122 14302 18302 14314
rect 18122 14250 18132 14302
rect 18166 14280 18302 14302
rect 17074 14230 17108 14246
rect 17074 14158 17108 14178
rect 17074 14086 17108 14110
rect 17074 14014 17108 14042
rect 17074 13942 17108 13974
rect 17074 13872 17108 13906
rect 17074 13804 17108 13836
rect 17074 13736 17108 13764
rect 17074 13668 17108 13692
rect 17074 13600 17108 13620
rect 17074 13532 17108 13548
rect 17074 13464 17108 13476
rect 17074 13396 17108 13404
rect 17074 13328 17108 13332
rect 17074 13222 17108 13226
rect 17074 13150 17108 13158
rect 17074 13078 17108 13090
rect 17074 13006 17108 13022
rect 17074 12934 17108 12954
rect 17074 12862 17108 12886
rect 17074 12790 17108 12818
rect 17074 12718 17108 12750
rect 17074 12648 17108 12682
rect 17074 12580 17108 12612
rect 17074 12512 17108 12540
rect 17074 12444 17108 12468
rect 17074 12376 17108 12396
rect 17074 12308 17108 12324
rect 17074 12240 17108 12252
rect 17074 12172 17108 12180
rect 17074 12104 17108 12108
rect 17074 11998 17108 12002
rect 17074 11926 17108 11934
rect 17074 11854 17108 11866
rect 17074 11773 17108 11798
rect 18166 14250 18266 14280
rect 18132 14230 18166 14246
rect 18132 14158 18166 14178
rect 18132 14086 18166 14110
rect 18132 14014 18166 14042
rect 18132 13942 18166 13974
rect 18132 13872 18166 13906
rect 18132 13804 18166 13836
rect 18132 13736 18166 13764
rect 18132 13668 18166 13692
rect 18132 13600 18166 13620
rect 18132 13532 18166 13548
rect 18132 13464 18166 13476
rect 18132 13396 18166 13404
rect 18132 13328 18166 13332
rect 18132 13222 18166 13226
rect 18132 13150 18166 13158
rect 18132 13078 18166 13090
rect 18132 13006 18166 13022
rect 18132 12934 18166 12954
rect 18132 12862 18166 12886
rect 18132 12790 18166 12818
rect 18132 12718 18166 12750
rect 18132 12648 18166 12682
rect 18132 12580 18166 12612
rect 18132 12512 18166 12540
rect 18132 12444 18166 12468
rect 18132 12376 18166 12396
rect 18132 12308 18166 12324
rect 18132 12240 18166 12252
rect 18132 12172 18166 12180
rect 18132 12104 18166 12108
rect 18132 11998 18166 12002
rect 18132 11926 18166 11934
rect 18132 11854 18166 11866
rect 18132 11773 18166 11798
rect 18300 14250 18302 14280
rect 18404 14740 18438 14774
rect 18404 14672 18438 14706
rect 18404 14604 18438 14638
rect 18404 14536 18438 14570
rect 18404 14468 18438 14502
rect 18404 14400 18438 14434
rect 18404 14332 18438 14366
rect 18404 14264 18438 14298
rect 18266 14212 18300 14246
rect 18266 14144 18300 14178
rect 18266 14076 18300 14110
rect 18266 14008 18300 14042
rect 18266 13940 18300 13974
rect 18266 13872 18300 13906
rect 18266 13804 18300 13838
rect 18266 13736 18300 13770
rect 18266 13668 18300 13702
rect 18266 13600 18300 13634
rect 18266 13532 18300 13566
rect 18266 13464 18300 13498
rect 18266 13396 18300 13430
rect 18266 13328 18300 13362
rect 18266 13260 18300 13294
rect 18266 13192 18300 13226
rect 18266 13124 18300 13158
rect 18266 13056 18300 13090
rect 18266 12988 18300 13022
rect 18266 12920 18300 12954
rect 18266 12852 18300 12886
rect 18266 12784 18300 12818
rect 18266 12716 18300 12750
rect 18266 12648 18300 12682
rect 18266 12580 18300 12614
rect 18266 12512 18300 12546
rect 18266 12444 18300 12478
rect 18266 12376 18300 12410
rect 18266 12308 18300 12342
rect 18266 12240 18300 12274
rect 18266 12172 18300 12206
rect 18266 12104 18300 12138
rect 18266 12036 18300 12070
rect 18266 11968 18300 12002
rect 18266 11900 18300 11934
rect 18266 11832 18300 11866
rect 18266 11764 18300 11798
rect 16940 11696 16974 11730
rect 17120 11696 17161 11730
rect 17205 11696 17229 11730
rect 17277 11696 17297 11730
rect 17349 11696 17365 11730
rect 17421 11696 17433 11730
rect 17493 11696 17501 11730
rect 17565 11696 17569 11730
rect 17671 11696 17675 11730
rect 17739 11696 17747 11730
rect 17807 11696 17819 11730
rect 17875 11696 17891 11730
rect 17943 11696 17963 11730
rect 18011 11696 18035 11730
rect 18079 11696 18120 11730
rect 18266 11696 18300 11730
rect 16940 11592 16974 11662
rect 18266 11592 18300 11662
rect 16940 11558 17059 11592
rect 17093 11558 17127 11592
rect 17161 11558 17195 11592
rect 17229 11558 17263 11592
rect 17297 11558 17331 11592
rect 17365 11558 17399 11592
rect 17433 11558 17467 11592
rect 17501 11558 17535 11592
rect 17569 11558 17603 11592
rect 17637 11558 17671 11592
rect 17705 11558 17739 11592
rect 17773 11558 17807 11592
rect 17841 11558 17875 11592
rect 17909 11558 17943 11592
rect 17977 11558 18011 11592
rect 18045 11558 18079 11592
rect 18113 11558 18147 11592
rect 18181 11558 18300 11592
rect 18404 14196 18438 14230
rect 18404 14128 18438 14162
rect 18404 14060 18438 14094
rect 18404 13992 18438 14026
rect 18404 13924 18438 13958
rect 18404 13856 18438 13890
rect 18404 13788 18438 13822
rect 18404 13720 18438 13754
rect 18404 13652 18438 13686
rect 18404 13584 18438 13618
rect 18404 13516 18438 13550
rect 18404 13448 18438 13482
rect 18404 13380 18438 13414
rect 18404 13312 18438 13346
rect 18404 13244 18438 13278
rect 18404 13176 18438 13210
rect 18404 13108 18438 13142
rect 18404 13040 18438 13074
rect 18404 12972 18438 13006
rect 18404 12904 18438 12938
rect 18404 12836 18438 12870
rect 18404 12768 18438 12802
rect 18404 12700 18438 12734
rect 18404 12632 18438 12666
rect 18404 12564 18438 12598
rect 18404 12496 18438 12530
rect 18404 12428 18438 12462
rect 18404 12360 18438 12394
rect 18404 12292 18438 12326
rect 18404 12224 18438 12258
rect 18404 12156 18438 12190
rect 18404 12088 18438 12122
rect 18404 12020 18438 12054
rect 18404 11952 18438 11986
rect 18404 11884 18438 11918
rect 18404 11816 18438 11850
rect 18404 11748 18438 11782
rect 18538 14740 18572 14765
rect 19596 14754 19630 14765
rect 19730 14754 19764 14774
rect 18538 14672 18572 14684
rect 18538 14604 18572 14612
rect 18538 14536 18572 14540
rect 18538 14430 18572 14434
rect 18538 14358 18572 14366
rect 18538 14286 18572 14298
rect 19586 14740 19766 14754
rect 19586 14684 19596 14740
rect 19630 14706 19730 14740
rect 19764 14706 19766 14740
rect 19630 14684 19766 14706
rect 19586 14672 19766 14684
rect 19586 14612 19596 14672
rect 19630 14638 19730 14672
rect 19764 14638 19766 14672
rect 19630 14612 19766 14638
rect 19586 14604 19766 14612
rect 19586 14540 19596 14604
rect 19630 14570 19730 14604
rect 19764 14570 19766 14604
rect 19630 14540 19766 14570
rect 19586 14536 19766 14540
rect 19586 14434 19596 14536
rect 19630 14502 19730 14536
rect 19764 14502 19766 14536
rect 19630 14468 19766 14502
rect 20382 14566 20497 14600
rect 20531 14566 20565 14600
rect 20599 14566 20633 14600
rect 20667 14566 20701 14600
rect 20735 14566 20769 14600
rect 20803 14566 20837 14600
rect 20871 14566 20905 14600
rect 20939 14566 20973 14600
rect 21007 14566 21041 14600
rect 21075 14566 21109 14600
rect 21143 14566 21177 14600
rect 21211 14566 21245 14600
rect 21279 14566 21313 14600
rect 21347 14566 21381 14600
rect 21415 14566 21449 14600
rect 21483 14566 21517 14600
rect 21551 14566 21666 14600
rect 20382 14474 20416 14566
rect 21632 14474 21666 14566
rect 19630 14434 19730 14468
rect 19764 14434 19766 14468
rect 19586 14430 19766 14434
rect 19586 14366 19596 14430
rect 19630 14400 19766 14430
rect 19630 14366 19730 14400
rect 19764 14366 19766 14400
rect 19586 14358 19766 14366
rect 19586 14298 19596 14358
rect 19630 14332 19766 14358
rect 19630 14298 19730 14332
rect 19764 14298 19766 14332
rect 19586 14286 19766 14298
rect 19586 14234 19596 14286
rect 19630 14264 19766 14286
rect 18538 14214 18572 14230
rect 18538 14142 18572 14162
rect 18538 14070 18572 14094
rect 18538 13998 18572 14026
rect 18538 13926 18572 13958
rect 18538 13856 18572 13890
rect 18538 13788 18572 13820
rect 18538 13720 18572 13748
rect 18538 13652 18572 13676
rect 18538 13584 18572 13604
rect 18538 13516 18572 13532
rect 18538 13448 18572 13460
rect 18538 13380 18572 13388
rect 18538 13312 18572 13316
rect 18538 13206 18572 13210
rect 18538 13134 18572 13142
rect 18538 13062 18572 13074
rect 18538 12990 18572 13006
rect 18538 12918 18572 12938
rect 18538 12846 18572 12870
rect 18538 12774 18572 12802
rect 18538 12702 18572 12734
rect 18538 12632 18572 12666
rect 18538 12564 18572 12596
rect 18538 12496 18572 12524
rect 18538 12428 18572 12452
rect 18538 12360 18572 12380
rect 18538 12292 18572 12308
rect 18538 12224 18572 12236
rect 18538 12156 18572 12164
rect 18538 12088 18572 12092
rect 18538 11982 18572 11986
rect 18538 11910 18572 11918
rect 18538 11838 18572 11850
rect 18538 11757 18572 11782
rect 19630 14234 19730 14264
rect 19596 14214 19630 14230
rect 19596 14142 19630 14162
rect 19596 14070 19630 14094
rect 19596 13998 19630 14026
rect 19596 13926 19630 13958
rect 19596 13856 19630 13890
rect 19596 13788 19630 13820
rect 19596 13720 19630 13748
rect 19596 13652 19630 13676
rect 19596 13584 19630 13604
rect 19596 13516 19630 13532
rect 19596 13448 19630 13460
rect 19596 13380 19630 13388
rect 19596 13312 19630 13316
rect 19596 13206 19630 13210
rect 19596 13134 19630 13142
rect 19596 13062 19630 13074
rect 19596 12990 19630 13006
rect 19596 12918 19630 12938
rect 19596 12846 19630 12870
rect 19596 12774 19630 12802
rect 19596 12702 19630 12734
rect 19596 12632 19630 12666
rect 19596 12564 19630 12596
rect 19596 12496 19630 12524
rect 19596 12428 19630 12452
rect 19596 12360 19630 12380
rect 19596 12292 19630 12308
rect 19596 12224 19630 12236
rect 19596 12156 19630 12164
rect 19596 12088 19630 12092
rect 19596 11982 19630 11986
rect 19596 11910 19630 11918
rect 19596 11838 19630 11850
rect 19596 11757 19630 11782
rect 19764 14234 19766 14264
rect 20376 14440 20382 14472
rect 20416 14470 20582 14472
rect 21464 14470 21632 14474
rect 20416 14440 20512 14470
rect 20376 14406 20512 14440
rect 20376 14372 20382 14406
rect 20416 14372 20512 14406
rect 20376 14338 20512 14372
rect 20376 14304 20382 14338
rect 20416 14304 20512 14338
rect 20376 14270 20512 14304
rect 20376 14236 20382 14270
rect 20416 14236 20512 14270
rect 19730 14196 19764 14230
rect 19730 14128 19764 14162
rect 19730 14060 19764 14094
rect 20376 14202 20512 14236
rect 20376 14168 20382 14202
rect 20416 14168 20512 14202
rect 20376 14134 20512 14168
rect 20376 14100 20382 14134
rect 20416 14100 20512 14134
rect 20376 14066 20512 14100
rect 20376 14036 20382 14066
rect 19730 13992 19764 14026
rect 19730 13924 19764 13958
rect 19730 13856 19764 13890
rect 19730 13788 19764 13822
rect 19730 13720 19764 13754
rect 19730 13652 19764 13686
rect 19730 13584 19764 13618
rect 19730 13516 19764 13550
rect 19730 13448 19764 13482
rect 19730 13380 19764 13414
rect 19730 13312 19764 13346
rect 19730 13244 19764 13278
rect 19730 13176 19764 13210
rect 19730 13108 19764 13142
rect 19730 13040 19764 13074
rect 19730 12972 19764 13006
rect 19730 12904 19764 12938
rect 19730 12836 19764 12870
rect 19730 12768 19764 12802
rect 19730 12700 19764 12734
rect 19730 12632 19764 12666
rect 19730 12564 19764 12598
rect 19730 12496 19764 12530
rect 19730 12428 19764 12462
rect 19730 12360 19764 12394
rect 19730 12292 19764 12326
rect 19730 12224 19764 12258
rect 19730 12156 19764 12190
rect 19730 12088 19764 12122
rect 19730 12020 19764 12054
rect 19730 11952 19764 11986
rect 19730 11884 19764 11918
rect 19730 11816 19764 11850
rect 19730 11748 19764 11782
rect 18404 11680 18438 11714
rect 18584 11680 18625 11714
rect 18669 11680 18693 11714
rect 18741 11680 18761 11714
rect 18813 11680 18829 11714
rect 18885 11680 18897 11714
rect 18957 11680 18965 11714
rect 19029 11680 19033 11714
rect 19135 11680 19139 11714
rect 19203 11680 19211 11714
rect 19271 11680 19283 11714
rect 19339 11680 19355 11714
rect 19407 11680 19427 11714
rect 19475 11680 19499 11714
rect 19543 11680 19584 11714
rect 19730 11680 19764 11714
rect 18404 11576 18438 11646
rect 19730 11576 19764 11646
rect 18404 11542 18523 11576
rect 18557 11542 18591 11576
rect 18625 11542 18659 11576
rect 18693 11542 18727 11576
rect 18761 11542 18795 11576
rect 18829 11542 18863 11576
rect 18897 11542 18931 11576
rect 18965 11542 18999 11576
rect 19033 11542 19067 11576
rect 19101 11542 19135 11576
rect 19169 11542 19203 11576
rect 19237 11542 19271 11576
rect 19305 11542 19339 11576
rect 19373 11542 19407 11576
rect 19441 11542 19475 11576
rect 19509 11542 19543 11576
rect 19577 11542 19611 11576
rect 19645 11542 19764 11576
rect 20416 14038 20512 14066
rect 21464 14038 21466 14470
rect 21536 14440 21632 14470
rect 21666 14440 21670 14474
rect 21536 14406 21670 14440
rect 21536 14372 21632 14406
rect 21666 14372 21670 14406
rect 21536 14338 21670 14372
rect 21536 14304 21632 14338
rect 21666 14304 21670 14338
rect 21536 14270 21670 14304
rect 21536 14236 21632 14270
rect 21666 14236 21670 14270
rect 21536 14202 21670 14236
rect 21536 14168 21632 14202
rect 21666 14168 21670 14202
rect 21536 14134 21670 14168
rect 21536 14100 21632 14134
rect 21666 14100 21670 14134
rect 21536 14066 21670 14100
rect 21536 14038 21632 14066
rect 20416 14036 20582 14038
rect 20382 13998 20416 14032
rect 20382 13930 20416 13964
rect 20382 13862 20416 13896
rect 20382 13794 20416 13828
rect 20382 13726 20416 13760
rect 20382 13658 20416 13692
rect 20382 13590 20416 13624
rect 20382 13522 20416 13556
rect 20382 13454 20416 13488
rect 20382 13386 20416 13420
rect 20382 13318 20416 13352
rect 20382 13250 20416 13284
rect 20382 13182 20416 13216
rect 20382 13114 20416 13148
rect 20382 13046 20416 13080
rect 20382 12978 20416 13012
rect 20382 12910 20416 12944
rect 20382 12842 20416 12876
rect 20382 12774 20416 12808
rect 20382 12706 20416 12740
rect 20382 12638 20416 12672
rect 20382 12570 20416 12604
rect 20382 12502 20416 12536
rect 20382 12434 20416 12468
rect 20382 12366 20416 12400
rect 20382 12298 20416 12332
rect 20382 12230 20416 12264
rect 20382 12162 20416 12196
rect 20382 12094 20416 12128
rect 20382 12026 20416 12060
rect 20382 11958 20416 11992
rect 20382 11890 20416 11924
rect 20382 11822 20416 11856
rect 20382 11754 20416 11788
rect 20382 11686 20416 11720
rect 20382 11618 20416 11652
rect 20382 11550 20416 11584
rect -9108 11501 -3289 11531
rect -9108 11375 -9016 11501
rect -9108 11341 -9081 11375
rect -9047 11341 -9016 11375
rect -9108 11307 -9016 11341
rect -9108 11273 -9081 11307
rect -9047 11273 -9016 11307
rect -9108 11239 -9016 11273
rect -9108 11205 -9081 11239
rect -9047 11205 -9016 11239
rect -3389 11335 -3289 11501
rect 20382 11482 20416 11516
rect 14820 11432 14924 11466
rect 14958 11432 14992 11466
rect 15026 11432 15060 11466
rect 15094 11432 15128 11466
rect 15162 11432 15196 11466
rect 15230 11432 15264 11466
rect 15298 11432 15332 11466
rect 15366 11432 15400 11466
rect 15434 11432 15468 11466
rect 15502 11432 15536 11466
rect 15570 11432 15604 11466
rect 15638 11432 15672 11466
rect 15706 11432 15740 11466
rect 15774 11432 15808 11466
rect 15842 11432 15876 11466
rect 15910 11432 15944 11466
rect 15978 11432 16012 11466
rect 16046 11432 16080 11466
rect 16114 11432 16148 11466
rect 16182 11432 16216 11466
rect 16250 11432 16284 11466
rect 16318 11432 16352 11466
rect 16386 11432 16420 11466
rect 16454 11432 16488 11466
rect 16522 11432 16556 11466
rect 16590 11432 16624 11466
rect 16658 11432 16692 11466
rect 16726 11432 16760 11466
rect 16794 11432 16828 11466
rect 16862 11432 16896 11466
rect 16930 11432 16964 11466
rect 16998 11432 17032 11466
rect 17066 11432 17100 11466
rect 17134 11432 17238 11466
rect 14820 11362 14854 11432
rect -3389 11301 -3355 11335
rect -3321 11301 -3289 11335
rect -3389 11267 -3289 11301
rect -9108 11171 -9016 11205
rect -8769 11202 -8722 11236
rect -8686 11202 -8652 11236
rect -8616 11202 -8569 11236
rect -8511 11202 -8464 11236
rect -8428 11202 -8394 11236
rect -8358 11202 -8311 11236
rect -8253 11202 -8206 11236
rect -8170 11202 -8136 11236
rect -8100 11202 -8053 11236
rect -7995 11202 -7948 11236
rect -7912 11202 -7878 11236
rect -7842 11202 -7795 11236
rect -7737 11202 -7690 11236
rect -7654 11202 -7620 11236
rect -7584 11202 -7537 11236
rect -7479 11202 -7432 11236
rect -7396 11202 -7362 11236
rect -7326 11202 -7279 11236
rect -7221 11202 -7174 11236
rect -7138 11202 -7104 11236
rect -7068 11202 -7021 11236
rect -6963 11202 -6916 11236
rect -6880 11202 -6846 11236
rect -6810 11202 -6763 11236
rect -6705 11202 -6658 11236
rect -6622 11202 -6588 11236
rect -6552 11202 -6505 11236
rect -6447 11202 -6400 11236
rect -6364 11202 -6330 11236
rect -6294 11202 -6247 11236
rect -6189 11202 -6142 11236
rect -6106 11202 -6072 11236
rect -6036 11202 -5989 11236
rect -5931 11202 -5884 11236
rect -5848 11202 -5814 11236
rect -5778 11202 -5731 11236
rect -5673 11202 -5626 11236
rect -5590 11202 -5556 11236
rect -5520 11202 -5473 11236
rect -5415 11202 -5368 11236
rect -5332 11202 -5298 11236
rect -5262 11202 -5215 11236
rect -5157 11202 -5110 11236
rect -5074 11202 -5040 11236
rect -5004 11202 -4957 11236
rect -4899 11202 -4852 11236
rect -4816 11202 -4782 11236
rect -4746 11202 -4699 11236
rect -4641 11202 -4594 11236
rect -4558 11202 -4524 11236
rect -4488 11202 -4441 11236
rect -4383 11202 -4336 11236
rect -4300 11202 -4266 11236
rect -4230 11202 -4183 11236
rect -4125 11202 -4078 11236
rect -4042 11202 -4008 11236
rect -3972 11202 -3925 11236
rect -3867 11202 -3820 11236
rect -3784 11202 -3750 11236
rect -3714 11202 -3667 11236
rect -3389 11233 -3355 11267
rect -3321 11233 -3289 11267
rect -9108 11137 -9081 11171
rect -9047 11137 -9016 11171
rect -3389 11199 -3289 11233
rect -9108 11103 -9016 11137
rect -9108 11069 -9081 11103
rect -9047 11069 -9016 11103
rect -9108 11035 -9016 11069
rect -9108 11001 -9081 11035
rect -9047 11001 -9016 11035
rect -9108 10967 -9016 11001
rect -9108 10933 -9081 10967
rect -9047 10933 -9016 10967
rect -9108 10899 -9016 10933
rect -9108 10865 -9081 10899
rect -9047 10865 -9016 10899
rect -9108 10831 -9016 10865
rect -9108 10797 -9081 10831
rect -9047 10797 -9016 10831
rect -9108 10763 -9016 10797
rect -9108 10729 -9081 10763
rect -9047 10729 -9016 10763
rect -9108 10695 -9016 10729
rect -9108 10661 -9081 10695
rect -9047 10661 -9016 10695
rect -9108 10627 -9016 10661
rect -9108 10593 -9081 10627
rect -9047 10593 -9016 10627
rect -9108 10559 -9016 10593
rect -9108 10525 -9081 10559
rect -9047 10525 -9016 10559
rect -9108 10491 -9016 10525
rect -9108 10457 -9081 10491
rect -9047 10457 -9016 10491
rect -9108 10423 -9016 10457
rect -9108 10389 -9081 10423
rect -9047 10389 -9016 10423
rect -9108 10355 -9016 10389
rect -9108 10321 -9081 10355
rect -9047 10321 -9016 10355
rect -9108 10287 -9016 10321
rect -9108 10253 -9081 10287
rect -9047 10253 -9016 10287
rect -9108 10219 -9016 10253
rect -9108 10185 -9081 10219
rect -9047 10185 -9016 10219
rect -9108 10151 -9016 10185
rect -8815 11149 -8781 11168
rect -8815 11077 -8781 11089
rect -8815 11005 -8781 11021
rect -8815 10933 -8781 10953
rect -8815 10861 -8781 10885
rect -8815 10789 -8781 10817
rect -8815 10717 -8781 10749
rect -8815 10647 -8781 10681
rect -8815 10579 -8781 10611
rect -8815 10511 -8781 10539
rect -8815 10443 -8781 10467
rect -8815 10375 -8781 10395
rect -8815 10307 -8781 10323
rect -8815 10239 -8781 10251
rect -8815 10160 -8781 10179
rect -8557 11149 -8523 11168
rect -8557 11077 -8523 11089
rect -8557 11005 -8523 11021
rect -8557 10933 -8523 10953
rect -8557 10861 -8523 10885
rect -8557 10789 -8523 10817
rect -8557 10717 -8523 10749
rect -8557 10647 -8523 10681
rect -8557 10579 -8523 10611
rect -8557 10511 -8523 10539
rect -8557 10443 -8523 10467
rect -8557 10375 -8523 10395
rect -8557 10307 -8523 10323
rect -8557 10239 -8523 10251
rect -8557 10160 -8523 10179
rect -8299 11149 -8265 11168
rect -8299 11077 -8265 11089
rect -8299 11005 -8265 11021
rect -8299 10933 -8265 10953
rect -8299 10861 -8265 10885
rect -8299 10789 -8265 10817
rect -8299 10717 -8265 10749
rect -8299 10647 -8265 10681
rect -8299 10579 -8265 10611
rect -8299 10511 -8265 10539
rect -8299 10443 -8265 10467
rect -8299 10375 -8265 10395
rect -8299 10307 -8265 10323
rect -8299 10239 -8265 10251
rect -8299 10160 -8265 10179
rect -8041 11149 -8007 11168
rect -8041 11077 -8007 11089
rect -8041 11005 -8007 11021
rect -8041 10933 -8007 10953
rect -8041 10861 -8007 10885
rect -8041 10789 -8007 10817
rect -8041 10717 -8007 10749
rect -8041 10647 -8007 10681
rect -8041 10579 -8007 10611
rect -8041 10511 -8007 10539
rect -8041 10443 -8007 10467
rect -8041 10375 -8007 10395
rect -8041 10307 -8007 10323
rect -8041 10239 -8007 10251
rect -8041 10160 -8007 10179
rect -7783 11149 -7749 11168
rect -7783 11077 -7749 11089
rect -7783 11005 -7749 11021
rect -7783 10933 -7749 10953
rect -7783 10861 -7749 10885
rect -7783 10789 -7749 10817
rect -7783 10717 -7749 10749
rect -7783 10647 -7749 10681
rect -7783 10579 -7749 10611
rect -7783 10511 -7749 10539
rect -7783 10443 -7749 10467
rect -7783 10375 -7749 10395
rect -7783 10307 -7749 10323
rect -7783 10239 -7749 10251
rect -7783 10160 -7749 10179
rect -7525 11149 -7491 11168
rect -7525 11077 -7491 11089
rect -7525 11005 -7491 11021
rect -7525 10933 -7491 10953
rect -7525 10861 -7491 10885
rect -7525 10789 -7491 10817
rect -7525 10717 -7491 10749
rect -7525 10647 -7491 10681
rect -7525 10579 -7491 10611
rect -7525 10511 -7491 10539
rect -7525 10443 -7491 10467
rect -7525 10375 -7491 10395
rect -7525 10307 -7491 10323
rect -7525 10239 -7491 10251
rect -7525 10160 -7491 10179
rect -7267 11149 -7233 11168
rect -7267 11077 -7233 11089
rect -7267 11005 -7233 11021
rect -7267 10933 -7233 10953
rect -7267 10861 -7233 10885
rect -7267 10789 -7233 10817
rect -7267 10717 -7233 10749
rect -7267 10647 -7233 10681
rect -7267 10579 -7233 10611
rect -7267 10511 -7233 10539
rect -7267 10443 -7233 10467
rect -7267 10375 -7233 10395
rect -7267 10307 -7233 10323
rect -7267 10239 -7233 10251
rect -7267 10160 -7233 10179
rect -7009 11149 -6975 11168
rect -7009 11077 -6975 11089
rect -7009 11005 -6975 11021
rect -7009 10933 -6975 10953
rect -7009 10861 -6975 10885
rect -7009 10789 -6975 10817
rect -7009 10717 -6975 10749
rect -7009 10647 -6975 10681
rect -7009 10579 -6975 10611
rect -7009 10511 -6975 10539
rect -7009 10443 -6975 10467
rect -7009 10375 -6975 10395
rect -7009 10307 -6975 10323
rect -7009 10239 -6975 10251
rect -7009 10160 -6975 10179
rect -6751 11149 -6717 11168
rect -6751 11077 -6717 11089
rect -6751 11005 -6717 11021
rect -6751 10933 -6717 10953
rect -6751 10861 -6717 10885
rect -6751 10789 -6717 10817
rect -6751 10717 -6717 10749
rect -6751 10647 -6717 10681
rect -6751 10579 -6717 10611
rect -6751 10511 -6717 10539
rect -6751 10443 -6717 10467
rect -6751 10375 -6717 10395
rect -6751 10307 -6717 10323
rect -6751 10239 -6717 10251
rect -6751 10160 -6717 10179
rect -6493 11149 -6459 11168
rect -6493 11077 -6459 11089
rect -6493 11005 -6459 11021
rect -6493 10933 -6459 10953
rect -6493 10861 -6459 10885
rect -6493 10789 -6459 10817
rect -6493 10717 -6459 10749
rect -6493 10647 -6459 10681
rect -6493 10579 -6459 10611
rect -6493 10511 -6459 10539
rect -6493 10443 -6459 10467
rect -6493 10375 -6459 10395
rect -6493 10307 -6459 10323
rect -6493 10239 -6459 10251
rect -6493 10160 -6459 10179
rect -6235 11149 -6201 11168
rect -6235 11077 -6201 11089
rect -6235 11005 -6201 11021
rect -6235 10933 -6201 10953
rect -6235 10861 -6201 10885
rect -6235 10789 -6201 10817
rect -6235 10717 -6201 10749
rect -6235 10647 -6201 10681
rect -6235 10579 -6201 10611
rect -6235 10511 -6201 10539
rect -6235 10443 -6201 10467
rect -6235 10375 -6201 10395
rect -6235 10307 -6201 10323
rect -6235 10239 -6201 10251
rect -6235 10160 -6201 10179
rect -5977 11149 -5943 11168
rect -5977 11077 -5943 11089
rect -5977 11005 -5943 11021
rect -5977 10933 -5943 10953
rect -5977 10861 -5943 10885
rect -5977 10789 -5943 10817
rect -5977 10717 -5943 10749
rect -5977 10647 -5943 10681
rect -5977 10579 -5943 10611
rect -5977 10511 -5943 10539
rect -5977 10443 -5943 10467
rect -5977 10375 -5943 10395
rect -5977 10307 -5943 10323
rect -5977 10239 -5943 10251
rect -5977 10160 -5943 10179
rect -5719 11149 -5685 11168
rect -5719 11077 -5685 11089
rect -5719 11005 -5685 11021
rect -5719 10933 -5685 10953
rect -5719 10861 -5685 10885
rect -5719 10789 -5685 10817
rect -5719 10717 -5685 10749
rect -5719 10647 -5685 10681
rect -5719 10579 -5685 10611
rect -5719 10511 -5685 10539
rect -5719 10443 -5685 10467
rect -5719 10375 -5685 10395
rect -5719 10307 -5685 10323
rect -5719 10239 -5685 10251
rect -5719 10160 -5685 10179
rect -5461 11149 -5427 11168
rect -5461 11077 -5427 11089
rect -5461 11005 -5427 11021
rect -5461 10933 -5427 10953
rect -5461 10861 -5427 10885
rect -5461 10789 -5427 10817
rect -5461 10717 -5427 10749
rect -5461 10647 -5427 10681
rect -5461 10579 -5427 10611
rect -5461 10511 -5427 10539
rect -5461 10443 -5427 10467
rect -5461 10375 -5427 10395
rect -5461 10307 -5427 10323
rect -5461 10239 -5427 10251
rect -5461 10160 -5427 10179
rect -5203 11149 -5169 11168
rect -5203 11077 -5169 11089
rect -5203 11005 -5169 11021
rect -5203 10933 -5169 10953
rect -5203 10861 -5169 10885
rect -5203 10789 -5169 10817
rect -5203 10717 -5169 10749
rect -5203 10647 -5169 10681
rect -5203 10579 -5169 10611
rect -5203 10511 -5169 10539
rect -5203 10443 -5169 10467
rect -5203 10375 -5169 10395
rect -5203 10307 -5169 10323
rect -5203 10239 -5169 10251
rect -5203 10160 -5169 10179
rect -4945 11149 -4911 11168
rect -4945 11077 -4911 11089
rect -4945 11005 -4911 11021
rect -4945 10933 -4911 10953
rect -4945 10861 -4911 10885
rect -4945 10789 -4911 10817
rect -4945 10717 -4911 10749
rect -4945 10647 -4911 10681
rect -4945 10579 -4911 10611
rect -4945 10511 -4911 10539
rect -4945 10443 -4911 10467
rect -4945 10375 -4911 10395
rect -4945 10307 -4911 10323
rect -4945 10239 -4911 10251
rect -4945 10160 -4911 10179
rect -4687 11149 -4653 11168
rect -4687 11077 -4653 11089
rect -4687 11005 -4653 11021
rect -4687 10933 -4653 10953
rect -4687 10861 -4653 10885
rect -4687 10789 -4653 10817
rect -4687 10717 -4653 10749
rect -4687 10647 -4653 10681
rect -4687 10579 -4653 10611
rect -4687 10511 -4653 10539
rect -4687 10443 -4653 10467
rect -4687 10375 -4653 10395
rect -4687 10307 -4653 10323
rect -4687 10239 -4653 10251
rect -4687 10160 -4653 10179
rect -4429 11149 -4395 11168
rect -4429 11077 -4395 11089
rect -4429 11005 -4395 11021
rect -4429 10933 -4395 10953
rect -4429 10861 -4395 10885
rect -4429 10789 -4395 10817
rect -4429 10717 -4395 10749
rect -4429 10647 -4395 10681
rect -4429 10579 -4395 10611
rect -4429 10511 -4395 10539
rect -4429 10443 -4395 10467
rect -4429 10375 -4395 10395
rect -4429 10307 -4395 10323
rect -4429 10239 -4395 10251
rect -4429 10160 -4395 10179
rect -4171 11149 -4137 11168
rect -4171 11077 -4137 11089
rect -4171 11005 -4137 11021
rect -4171 10933 -4137 10953
rect -4171 10861 -4137 10885
rect -4171 10789 -4137 10817
rect -4171 10717 -4137 10749
rect -4171 10647 -4137 10681
rect -4171 10579 -4137 10611
rect -4171 10511 -4137 10539
rect -4171 10443 -4137 10467
rect -4171 10375 -4137 10395
rect -4171 10307 -4137 10323
rect -4171 10239 -4137 10251
rect -4171 10160 -4137 10179
rect -3913 11149 -3879 11168
rect -3913 11077 -3879 11089
rect -3913 11005 -3879 11021
rect -3913 10933 -3879 10953
rect -3913 10861 -3879 10885
rect -3913 10789 -3879 10817
rect -3913 10717 -3879 10749
rect -3913 10647 -3879 10681
rect -3913 10579 -3879 10611
rect -3913 10511 -3879 10539
rect -3913 10443 -3879 10467
rect -3913 10375 -3879 10395
rect -3913 10307 -3879 10323
rect -3913 10239 -3879 10251
rect -3913 10160 -3879 10179
rect -3655 11149 -3621 11168
rect -3655 11077 -3621 11089
rect -3655 11005 -3621 11021
rect -3655 10933 -3621 10953
rect -3655 10861 -3621 10885
rect -3655 10789 -3621 10817
rect -3655 10717 -3621 10749
rect -3655 10647 -3621 10681
rect -3655 10579 -3621 10611
rect -3655 10511 -3621 10539
rect -3655 10443 -3621 10467
rect -3655 10375 -3621 10395
rect -3655 10307 -3621 10323
rect -3655 10239 -3621 10251
rect -3655 10160 -3621 10179
rect -3389 11165 -3355 11199
rect -3321 11165 -3289 11199
rect -3389 11131 -3289 11165
rect -3389 11097 -3355 11131
rect -3321 11097 -3289 11131
rect -3389 11063 -3289 11097
rect -3389 11029 -3355 11063
rect -3321 11029 -3289 11063
rect -3389 10995 -3289 11029
rect -3389 10961 -3355 10995
rect -3321 10961 -3289 10995
rect -3389 10927 -3289 10961
rect -3389 10893 -3355 10927
rect -3321 10893 -3289 10927
rect -3389 10859 -3289 10893
rect -3389 10825 -3355 10859
rect -3321 10825 -3289 10859
rect -3389 10791 -3289 10825
rect -3389 10757 -3355 10791
rect -3321 10757 -3289 10791
rect -3389 10723 -3289 10757
rect -3389 10689 -3355 10723
rect -3321 10689 -3289 10723
rect -3389 10655 -3289 10689
rect -3389 10621 -3355 10655
rect -3321 10621 -3289 10655
rect -3389 10587 -3289 10621
rect -3389 10553 -3355 10587
rect -3321 10553 -3289 10587
rect -3389 10519 -3289 10553
rect -3389 10485 -3355 10519
rect -3321 10485 -3289 10519
rect -3389 10451 -3289 10485
rect -3389 10417 -3355 10451
rect -3321 10417 -3289 10451
rect -3389 10383 -3289 10417
rect -3389 10349 -3355 10383
rect -3321 10349 -3289 10383
rect -3389 10315 -3289 10349
rect -3389 10281 -3355 10315
rect -3321 10281 -3289 10315
rect -3389 10247 -3289 10281
rect -3389 10213 -3355 10247
rect -3321 10213 -3289 10247
rect -3389 10179 -3289 10213
rect -9108 10117 -9081 10151
rect -9047 10117 -9016 10151
rect -3389 10145 -3355 10179
rect -3321 10145 -3289 10179
rect -9108 10083 -9016 10117
rect -8769 10092 -8722 10126
rect -8686 10092 -8652 10126
rect -8616 10092 -8569 10126
rect -8511 10092 -8464 10126
rect -8428 10092 -8394 10126
rect -8358 10092 -8311 10126
rect -8253 10092 -8206 10126
rect -8170 10092 -8136 10126
rect -8100 10092 -8053 10126
rect -7995 10092 -7948 10126
rect -7912 10092 -7878 10126
rect -7842 10092 -7795 10126
rect -7737 10092 -7690 10126
rect -7654 10092 -7620 10126
rect -7584 10092 -7537 10126
rect -7479 10092 -7432 10126
rect -7396 10092 -7362 10126
rect -7326 10092 -7279 10126
rect -7221 10092 -7174 10126
rect -7138 10092 -7104 10126
rect -7068 10092 -7021 10126
rect -6963 10092 -6916 10126
rect -6880 10092 -6846 10126
rect -6810 10092 -6763 10126
rect -6705 10092 -6658 10126
rect -6622 10092 -6588 10126
rect -6552 10092 -6505 10126
rect -6447 10092 -6400 10126
rect -6364 10092 -6330 10126
rect -6294 10092 -6247 10126
rect -6189 10092 -6142 10126
rect -6106 10092 -6072 10126
rect -6036 10092 -5989 10126
rect -5931 10092 -5884 10126
rect -5848 10092 -5814 10126
rect -5778 10092 -5731 10126
rect -5673 10092 -5626 10126
rect -5590 10092 -5556 10126
rect -5520 10092 -5473 10126
rect -5415 10092 -5368 10126
rect -5332 10092 -5298 10126
rect -5262 10092 -5215 10126
rect -5157 10092 -5110 10126
rect -5074 10092 -5040 10126
rect -5004 10092 -4957 10126
rect -4899 10092 -4852 10126
rect -4816 10092 -4782 10126
rect -4746 10092 -4699 10126
rect -4641 10092 -4594 10126
rect -4558 10092 -4524 10126
rect -4488 10092 -4441 10126
rect -4383 10092 -4336 10126
rect -4300 10092 -4266 10126
rect -4230 10092 -4183 10126
rect -4125 10092 -4078 10126
rect -4042 10092 -4008 10126
rect -3972 10092 -3925 10126
rect -3867 10092 -3820 10126
rect -3784 10092 -3750 10126
rect -3714 10092 -3667 10126
rect -3389 10111 -3289 10145
rect -9108 10049 -9081 10083
rect -9047 10049 -9016 10083
rect -9108 10015 -9016 10049
rect -9108 9981 -9081 10015
rect -9047 9981 -9016 10015
rect -9108 9947 -9016 9981
rect -9108 9913 -9081 9947
rect -9047 9913 -9016 9947
rect -9108 9879 -9016 9913
rect -9108 9845 -9081 9879
rect -9047 9845 -9016 9879
rect -3389 10077 -3355 10111
rect -3321 10077 -3289 10111
rect -3389 10043 -3289 10077
rect -3389 10009 -3355 10043
rect -3321 10009 -3289 10043
rect -3389 9975 -3289 10009
rect -3389 9941 -3355 9975
rect -3321 9941 -3289 9975
rect -3389 9907 -3289 9941
rect -3389 9873 -3355 9907
rect -3321 9873 -3289 9907
rect -9108 9811 -9016 9845
rect -7734 9837 -7687 9871
rect -7651 9837 -7617 9871
rect -7581 9837 -7534 9871
rect -7268 9837 -7221 9871
rect -7185 9837 -7151 9871
rect -7115 9837 -7068 9871
rect -7010 9837 -6963 9871
rect -6927 9837 -6893 9871
rect -6857 9837 -6810 9871
rect -6752 9837 -6705 9871
rect -6669 9837 -6635 9871
rect -6599 9837 -6552 9871
rect -6494 9837 -6447 9871
rect -6411 9837 -6377 9871
rect -6341 9837 -6294 9871
rect -6236 9837 -6189 9871
rect -6153 9837 -6119 9871
rect -6083 9837 -6036 9871
rect -5978 9837 -5931 9871
rect -5895 9837 -5861 9871
rect -5825 9837 -5778 9871
rect -5720 9837 -5673 9871
rect -5637 9837 -5603 9871
rect -5567 9837 -5520 9871
rect -5462 9837 -5415 9871
rect -5379 9837 -5345 9871
rect -5309 9837 -5262 9871
rect -5204 9837 -5157 9871
rect -5121 9837 -5087 9871
rect -5051 9837 -5004 9871
rect -4946 9837 -4899 9871
rect -4863 9837 -4829 9871
rect -4793 9837 -4746 9871
rect -3389 9839 -3289 9873
rect -9108 9777 -9081 9811
rect -9047 9777 -9016 9811
rect -3389 9805 -3355 9839
rect -3321 9805 -3289 9839
rect -9108 9743 -9016 9777
rect -9108 9709 -9081 9743
rect -9047 9709 -9016 9743
rect -9108 9675 -9016 9709
rect -9108 9641 -9081 9675
rect -9047 9641 -9016 9675
rect -9108 9607 -9016 9641
rect -9108 9573 -9081 9607
rect -9047 9573 -9016 9607
rect -9108 9539 -9016 9573
rect -9108 9505 -9081 9539
rect -9047 9505 -9016 9539
rect -9108 9471 -9016 9505
rect -9108 9437 -9081 9471
rect -9047 9437 -9016 9471
rect -9108 9403 -9016 9437
rect -9108 9369 -9081 9403
rect -9047 9369 -9016 9403
rect -9108 9335 -9016 9369
rect -9108 9301 -9081 9335
rect -9047 9301 -9016 9335
rect -9108 9267 -9016 9301
rect -9108 9233 -9081 9267
rect -9047 9233 -9016 9267
rect -9108 9199 -9016 9233
rect -9108 9165 -9081 9199
rect -9047 9165 -9016 9199
rect -9108 9131 -9016 9165
rect -9108 9097 -9081 9131
rect -9047 9097 -9016 9131
rect -9108 9063 -9016 9097
rect -9108 9029 -9081 9063
rect -9047 9029 -9016 9063
rect -9108 8995 -9016 9029
rect -9108 8961 -9081 8995
rect -9047 8961 -9016 8995
rect -9108 8927 -9016 8961
rect -9108 8893 -9081 8927
rect -9047 8893 -9016 8927
rect -9108 8859 -9016 8893
rect -9108 8825 -9081 8859
rect -9047 8825 -9016 8859
rect -9108 8791 -9016 8825
rect -7780 9784 -7746 9803
rect -7780 9712 -7746 9724
rect -7780 9640 -7746 9656
rect -7780 9568 -7746 9588
rect -7780 9496 -7746 9520
rect -7780 9424 -7746 9452
rect -7780 9352 -7746 9384
rect -7780 9282 -7746 9316
rect -7780 9214 -7746 9246
rect -7780 9146 -7746 9174
rect -7780 9078 -7746 9102
rect -7780 9010 -7746 9030
rect -7780 8942 -7746 8958
rect -7780 8874 -7746 8886
rect -7780 8795 -7746 8814
rect -7522 9784 -7488 9803
rect -7522 9712 -7488 9724
rect -7522 9640 -7488 9656
rect -7522 9568 -7488 9588
rect -7522 9496 -7488 9520
rect -7522 9424 -7488 9452
rect -7522 9352 -7488 9384
rect -7522 9282 -7488 9316
rect -7522 9214 -7488 9246
rect -7522 9146 -7488 9174
rect -7522 9078 -7488 9102
rect -7522 9010 -7488 9030
rect -7522 8942 -7488 8958
rect -7522 8874 -7488 8886
rect -7522 8795 -7488 8814
rect -7314 9784 -7280 9803
rect -7314 9712 -7280 9724
rect -7314 9640 -7280 9656
rect -7314 9568 -7280 9588
rect -7314 9496 -7280 9520
rect -7314 9424 -7280 9452
rect -7314 9352 -7280 9384
rect -7314 9282 -7280 9316
rect -7314 9214 -7280 9246
rect -7314 9146 -7280 9174
rect -7314 9078 -7280 9102
rect -7314 9010 -7280 9030
rect -7314 8942 -7280 8958
rect -7314 8874 -7280 8886
rect -7314 8795 -7280 8814
rect -7056 9784 -7022 9803
rect -7056 9712 -7022 9724
rect -7056 9640 -7022 9656
rect -7056 9568 -7022 9588
rect -7056 9496 -7022 9520
rect -7056 9424 -7022 9452
rect -7056 9352 -7022 9384
rect -7056 9282 -7022 9316
rect -7056 9214 -7022 9246
rect -7056 9146 -7022 9174
rect -7056 9078 -7022 9102
rect -7056 9010 -7022 9030
rect -7056 8942 -7022 8958
rect -7056 8874 -7022 8886
rect -7056 8795 -7022 8814
rect -6798 9784 -6764 9803
rect -6798 9712 -6764 9724
rect -6798 9640 -6764 9656
rect -6798 9568 -6764 9588
rect -6798 9496 -6764 9520
rect -6798 9424 -6764 9452
rect -6798 9352 -6764 9384
rect -6798 9282 -6764 9316
rect -6798 9214 -6764 9246
rect -6798 9146 -6764 9174
rect -6798 9078 -6764 9102
rect -6798 9010 -6764 9030
rect -6798 8942 -6764 8958
rect -6798 8874 -6764 8886
rect -6798 8795 -6764 8814
rect -6540 9784 -6506 9803
rect -6540 9712 -6506 9724
rect -6540 9640 -6506 9656
rect -6540 9568 -6506 9588
rect -6540 9496 -6506 9520
rect -6540 9424 -6506 9452
rect -6540 9352 -6506 9384
rect -6540 9282 -6506 9316
rect -6540 9214 -6506 9246
rect -6540 9146 -6506 9174
rect -6540 9078 -6506 9102
rect -6540 9010 -6506 9030
rect -6540 8942 -6506 8958
rect -6540 8874 -6506 8886
rect -6540 8795 -6506 8814
rect -6282 9784 -6248 9803
rect -6282 9712 -6248 9724
rect -6282 9640 -6248 9656
rect -6282 9568 -6248 9588
rect -6282 9496 -6248 9520
rect -6282 9424 -6248 9452
rect -6282 9352 -6248 9384
rect -6282 9282 -6248 9316
rect -6282 9214 -6248 9246
rect -6282 9146 -6248 9174
rect -6282 9078 -6248 9102
rect -6282 9010 -6248 9030
rect -6282 8942 -6248 8958
rect -6282 8874 -6248 8886
rect -6282 8795 -6248 8814
rect -6024 9784 -5990 9803
rect -6024 9712 -5990 9724
rect -6024 9640 -5990 9656
rect -6024 9568 -5990 9588
rect -6024 9496 -5990 9520
rect -6024 9424 -5990 9452
rect -6024 9352 -5990 9384
rect -6024 9282 -5990 9316
rect -6024 9214 -5990 9246
rect -6024 9146 -5990 9174
rect -6024 9078 -5990 9102
rect -6024 9010 -5990 9030
rect -6024 8942 -5990 8958
rect -6024 8874 -5990 8886
rect -6024 8795 -5990 8814
rect -5766 9784 -5732 9803
rect -5766 9712 -5732 9724
rect -5766 9640 -5732 9656
rect -5766 9568 -5732 9588
rect -5766 9496 -5732 9520
rect -5766 9424 -5732 9452
rect -5766 9352 -5732 9384
rect -5766 9282 -5732 9316
rect -5766 9214 -5732 9246
rect -5766 9146 -5732 9174
rect -5766 9078 -5732 9102
rect -5766 9010 -5732 9030
rect -5766 8942 -5732 8958
rect -5766 8874 -5732 8886
rect -5766 8795 -5732 8814
rect -5508 9784 -5474 9803
rect -5508 9712 -5474 9724
rect -5508 9640 -5474 9656
rect -5508 9568 -5474 9588
rect -5508 9496 -5474 9520
rect -5508 9424 -5474 9452
rect -5508 9352 -5474 9384
rect -5508 9282 -5474 9316
rect -5508 9214 -5474 9246
rect -5508 9146 -5474 9174
rect -5508 9078 -5474 9102
rect -5508 9010 -5474 9030
rect -5508 8942 -5474 8958
rect -5508 8874 -5474 8886
rect -5508 8795 -5474 8814
rect -5250 9784 -5216 9803
rect -5250 9712 -5216 9724
rect -5250 9640 -5216 9656
rect -5250 9568 -5216 9588
rect -5250 9496 -5216 9520
rect -5250 9424 -5216 9452
rect -5250 9352 -5216 9384
rect -5250 9282 -5216 9316
rect -5250 9214 -5216 9246
rect -5250 9146 -5216 9174
rect -5250 9078 -5216 9102
rect -5250 9010 -5216 9030
rect -5250 8942 -5216 8958
rect -5250 8874 -5216 8886
rect -5250 8795 -5216 8814
rect -4992 9784 -4958 9803
rect -4992 9712 -4958 9724
rect -4992 9640 -4958 9656
rect -4992 9568 -4958 9588
rect -4992 9496 -4958 9520
rect -4992 9424 -4958 9452
rect -4992 9352 -4958 9384
rect -4992 9282 -4958 9316
rect -4992 9214 -4958 9246
rect -4992 9146 -4958 9174
rect -4992 9078 -4958 9102
rect -4992 9010 -4958 9030
rect -4992 8942 -4958 8958
rect -4992 8874 -4958 8886
rect -4992 8795 -4958 8814
rect -4734 9784 -4700 9803
rect -4734 9712 -4700 9724
rect -4734 9640 -4700 9656
rect -4734 9568 -4700 9588
rect -4734 9496 -4700 9520
rect -4734 9424 -4700 9452
rect -4734 9352 -4700 9384
rect -4734 9282 -4700 9316
rect -4734 9214 -4700 9246
rect -4734 9146 -4700 9174
rect -4734 9078 -4700 9102
rect -4734 9010 -4700 9030
rect -4734 8942 -4700 8958
rect -4734 8874 -4700 8886
rect -4734 8795 -4700 8814
rect -3389 9771 -3289 9805
rect -3389 9737 -3355 9771
rect -3321 9737 -3289 9771
rect -3389 9703 -3289 9737
rect -3389 9669 -3355 9703
rect -3321 9669 -3289 9703
rect -3389 9635 -3289 9669
rect -3389 9601 -3355 9635
rect -3321 9601 -3289 9635
rect -3389 9567 -3289 9601
rect -3389 9533 -3355 9567
rect -3321 9533 -3289 9567
rect -3389 9499 -3289 9533
rect -3389 9465 -3355 9499
rect -3321 9465 -3289 9499
rect -3389 9431 -3289 9465
rect -3389 9397 -3355 9431
rect -3321 9397 -3289 9431
rect -3389 9363 -3289 9397
rect -3389 9329 -3355 9363
rect -3321 9329 -3289 9363
rect -3389 9295 -3289 9329
rect -3389 9261 -3355 9295
rect -3321 9261 -3289 9295
rect -3389 9227 -3289 9261
rect -3389 9193 -3355 9227
rect -3321 9193 -3289 9227
rect -3389 9159 -3289 9193
rect -3389 9125 -3355 9159
rect -3321 9125 -3289 9159
rect -3389 9091 -3289 9125
rect -3389 9057 -3355 9091
rect -3321 9057 -3289 9091
rect -3389 9023 -3289 9057
rect -3389 8989 -3355 9023
rect -3321 8989 -3289 9023
rect -3389 8955 -3289 8989
rect -3389 8921 -3355 8955
rect -3321 8921 -3289 8955
rect -3389 8887 -3289 8921
rect -3389 8853 -3355 8887
rect -3321 8853 -3289 8887
rect -3389 8819 -3289 8853
rect -9108 8757 -9081 8791
rect -9047 8757 -9016 8791
rect -3389 8785 -3355 8819
rect -3321 8785 -3289 8819
rect -9108 8723 -9016 8757
rect -7734 8727 -7687 8761
rect -7651 8727 -7617 8761
rect -7581 8727 -7534 8761
rect -7268 8727 -7221 8761
rect -7185 8727 -7151 8761
rect -7115 8727 -7068 8761
rect -7010 8727 -6963 8761
rect -6927 8727 -6893 8761
rect -6857 8727 -6810 8761
rect -6752 8727 -6705 8761
rect -6669 8727 -6635 8761
rect -6599 8727 -6552 8761
rect -6494 8727 -6447 8761
rect -6411 8727 -6377 8761
rect -6341 8727 -6294 8761
rect -6236 8727 -6189 8761
rect -6153 8727 -6119 8761
rect -6083 8727 -6036 8761
rect -5978 8727 -5931 8761
rect -5895 8727 -5861 8761
rect -5825 8727 -5778 8761
rect -5720 8727 -5673 8761
rect -5637 8727 -5603 8761
rect -5567 8727 -5520 8761
rect -5462 8727 -5415 8761
rect -5379 8727 -5345 8761
rect -5309 8727 -5262 8761
rect -5204 8727 -5157 8761
rect -5121 8727 -5087 8761
rect -5051 8727 -5004 8761
rect -4946 8727 -4899 8761
rect -4863 8727 -4829 8761
rect -4793 8727 -4746 8761
rect -3389 8751 -3289 8785
rect -9108 8689 -9081 8723
rect -9047 8689 -9016 8723
rect -9108 8655 -9016 8689
rect -9108 8621 -9081 8655
rect -9047 8621 -9016 8655
rect -9108 8429 -9016 8621
rect -3389 8717 -3355 8751
rect -3321 8717 -3289 8751
rect -3389 8683 -3289 8717
rect -3389 8649 -3355 8683
rect -3321 8649 -3289 8683
rect -3389 8615 -3289 8649
rect -3389 8581 -3355 8615
rect -3321 8581 -3289 8615
rect -3389 8429 -3289 8581
rect -9108 8399 -3289 8429
rect -9108 8365 -8813 8399
rect -8779 8365 -8745 8399
rect -8711 8365 -8677 8399
rect -8643 8365 -8609 8399
rect -8575 8365 -8541 8399
rect -8507 8365 -8473 8399
rect -8439 8365 -8405 8399
rect -8371 8365 -8337 8399
rect -8303 8365 -8269 8399
rect -8235 8365 -8201 8399
rect -8167 8365 -8133 8399
rect -8099 8365 -8065 8399
rect -8031 8365 -7997 8399
rect -7963 8365 -7929 8399
rect -7895 8365 -7861 8399
rect -7827 8365 -7793 8399
rect -7759 8365 -7725 8399
rect -7691 8365 -7657 8399
rect -7623 8365 -7589 8399
rect -7555 8365 -7521 8399
rect -7487 8365 -7453 8399
rect -7419 8365 -7385 8399
rect -7351 8365 -7317 8399
rect -7283 8365 -7249 8399
rect -7215 8365 -7181 8399
rect -7147 8365 -7113 8399
rect -7079 8365 -7045 8399
rect -7011 8365 -6977 8399
rect -6943 8365 -6909 8399
rect -6875 8365 -6841 8399
rect -6807 8365 -6773 8399
rect -6739 8365 -6705 8399
rect -6671 8365 -6637 8399
rect -6603 8365 -6569 8399
rect -6535 8365 -6501 8399
rect -6467 8365 -6433 8399
rect -6399 8365 -6365 8399
rect -6331 8365 -6297 8399
rect -6263 8365 -6229 8399
rect -6195 8365 -6161 8399
rect -6127 8365 -6093 8399
rect -6059 8365 -6025 8399
rect -5991 8365 -5957 8399
rect -5923 8365 -5889 8399
rect -5855 8365 -5821 8399
rect -5787 8365 -5753 8399
rect -5719 8365 -5685 8399
rect -5651 8365 -5617 8399
rect -5583 8365 -5549 8399
rect -5515 8365 -5481 8399
rect -5447 8365 -5413 8399
rect -5379 8365 -5345 8399
rect -5311 8365 -5277 8399
rect -5243 8365 -5209 8399
rect -5175 8365 -5141 8399
rect -5107 8365 -5073 8399
rect -5039 8365 -5005 8399
rect -4971 8365 -4937 8399
rect -4903 8365 -4869 8399
rect -4835 8365 -4801 8399
rect -4767 8365 -4733 8399
rect -4699 8365 -4665 8399
rect -4631 8365 -4597 8399
rect -4563 8365 -4529 8399
rect -4495 8365 -4461 8399
rect -4427 8365 -4393 8399
rect -4359 8365 -4325 8399
rect -4291 8365 -4257 8399
rect -4223 8365 -4189 8399
rect -4155 8365 -4121 8399
rect -4087 8365 -4053 8399
rect -4019 8365 -3985 8399
rect -3951 8365 -3917 8399
rect -3883 8365 -3849 8399
rect -3815 8365 -3781 8399
rect -3747 8365 -3713 8399
rect -3679 8365 -3645 8399
rect -3611 8365 -3577 8399
rect -3543 8365 -3289 8399
rect -9108 8337 -3289 8365
rect 12756 11334 12871 11357
rect 12756 11299 14070 11334
rect 12756 11276 12912 11299
rect 12756 11242 12816 11276
rect 12850 11265 12912 11276
rect 12946 11265 13002 11299
rect 13036 11265 13092 11299
rect 13126 11265 13182 11299
rect 13216 11265 13272 11299
rect 13306 11265 13362 11299
rect 13396 11265 13452 11299
rect 13486 11265 13542 11299
rect 13576 11265 13632 11299
rect 13666 11265 13722 11299
rect 13756 11265 13812 11299
rect 13846 11265 13902 11299
rect 13936 11276 14070 11299
rect 13936 11265 14003 11276
rect 12850 11242 14003 11265
rect 14037 11242 14070 11276
rect 12756 11235 14070 11242
rect 12756 11186 12881 11235
rect 12756 11152 12816 11186
rect 12850 11152 12881 11186
rect 13971 11186 14070 11235
rect 12756 11096 12881 11152
rect 12756 11062 12816 11096
rect 12850 11062 12881 11096
rect 12756 11006 12881 11062
rect 12756 10972 12816 11006
rect 12850 10972 12881 11006
rect 12756 10916 12881 10972
rect 12756 10882 12816 10916
rect 12850 10882 12881 10916
rect 12756 10826 12881 10882
rect 12756 10792 12816 10826
rect 12850 10792 12881 10826
rect 12756 10736 12881 10792
rect 12756 10702 12816 10736
rect 12850 10702 12881 10736
rect 12756 10646 12881 10702
rect 12756 10612 12816 10646
rect 12850 10612 12881 10646
rect 12756 10556 12881 10612
rect 12756 10522 12816 10556
rect 12850 10522 12881 10556
rect 12756 10466 12881 10522
rect 12756 10432 12816 10466
rect 12850 10432 12881 10466
rect 12756 10376 12881 10432
rect 12756 10342 12816 10376
rect 12850 10342 12881 10376
rect 12756 10286 12881 10342
rect 12756 10252 12816 10286
rect 12850 10252 12881 10286
rect 12756 10196 12881 10252
rect 12945 11152 13907 11171
rect 12945 11118 13076 11152
rect 13110 11118 13166 11152
rect 13200 11118 13256 11152
rect 13290 11118 13346 11152
rect 13380 11118 13436 11152
rect 13470 11118 13526 11152
rect 13560 11118 13616 11152
rect 13650 11118 13706 11152
rect 13740 11118 13796 11152
rect 13830 11118 13907 11152
rect 12945 11099 13907 11118
rect 12945 11095 13017 11099
rect 12945 11061 12964 11095
rect 12998 11061 13017 11095
rect 12945 11005 13017 11061
rect 13835 11076 13907 11099
rect 13835 11042 13854 11076
rect 13888 11042 13907 11076
rect 12945 10971 12964 11005
rect 12998 10971 13017 11005
rect 12945 10915 13017 10971
rect 12945 10881 12964 10915
rect 12998 10881 13017 10915
rect 12945 10825 13017 10881
rect 12945 10791 12964 10825
rect 12998 10791 13017 10825
rect 12945 10735 13017 10791
rect 12945 10701 12964 10735
rect 12998 10701 13017 10735
rect 12945 10645 13017 10701
rect 12945 10611 12964 10645
rect 12998 10611 13017 10645
rect 12945 10555 13017 10611
rect 12945 10521 12964 10555
rect 12998 10521 13017 10555
rect 12945 10465 13017 10521
rect 12945 10431 12964 10465
rect 12998 10431 13017 10465
rect 12945 10375 13017 10431
rect 12945 10341 12964 10375
rect 12998 10341 13017 10375
rect 13079 10978 13773 11037
rect 13079 10944 13140 10978
rect 13174 10950 13230 10978
rect 13264 10950 13320 10978
rect 13354 10950 13410 10978
rect 13186 10944 13230 10950
rect 13286 10944 13320 10950
rect 13386 10944 13410 10950
rect 13444 10950 13500 10978
rect 13444 10944 13452 10950
rect 13079 10916 13152 10944
rect 13186 10916 13252 10944
rect 13286 10916 13352 10944
rect 13386 10916 13452 10944
rect 13486 10944 13500 10950
rect 13534 10950 13590 10978
rect 13534 10944 13552 10950
rect 13486 10916 13552 10944
rect 13586 10944 13590 10950
rect 13624 10950 13680 10978
rect 13624 10944 13652 10950
rect 13714 10944 13773 10978
rect 13586 10916 13652 10944
rect 13686 10916 13773 10944
rect 13079 10888 13773 10916
rect 13079 10854 13140 10888
rect 13174 10854 13230 10888
rect 13264 10854 13320 10888
rect 13354 10854 13410 10888
rect 13444 10854 13500 10888
rect 13534 10854 13590 10888
rect 13624 10854 13680 10888
rect 13714 10854 13773 10888
rect 13079 10850 13773 10854
rect 13079 10816 13152 10850
rect 13186 10816 13252 10850
rect 13286 10816 13352 10850
rect 13386 10816 13452 10850
rect 13486 10816 13552 10850
rect 13586 10816 13652 10850
rect 13686 10816 13773 10850
rect 13079 10798 13773 10816
rect 13079 10764 13140 10798
rect 13174 10764 13230 10798
rect 13264 10764 13320 10798
rect 13354 10764 13410 10798
rect 13444 10764 13500 10798
rect 13534 10764 13590 10798
rect 13624 10764 13680 10798
rect 13714 10764 13773 10798
rect 13079 10750 13773 10764
rect 13079 10716 13152 10750
rect 13186 10716 13252 10750
rect 13286 10716 13352 10750
rect 13386 10716 13452 10750
rect 13486 10716 13552 10750
rect 13586 10716 13652 10750
rect 13686 10716 13773 10750
rect 13079 10708 13773 10716
rect 13079 10674 13140 10708
rect 13174 10674 13230 10708
rect 13264 10674 13320 10708
rect 13354 10674 13410 10708
rect 13444 10674 13500 10708
rect 13534 10674 13590 10708
rect 13624 10674 13680 10708
rect 13714 10674 13773 10708
rect 13079 10650 13773 10674
rect 13079 10618 13152 10650
rect 13186 10618 13252 10650
rect 13286 10618 13352 10650
rect 13386 10618 13452 10650
rect 13079 10584 13140 10618
rect 13186 10616 13230 10618
rect 13286 10616 13320 10618
rect 13386 10616 13410 10618
rect 13174 10584 13230 10616
rect 13264 10584 13320 10616
rect 13354 10584 13410 10616
rect 13444 10616 13452 10618
rect 13486 10618 13552 10650
rect 13486 10616 13500 10618
rect 13444 10584 13500 10616
rect 13534 10616 13552 10618
rect 13586 10618 13652 10650
rect 13686 10618 13773 10650
rect 13586 10616 13590 10618
rect 13534 10584 13590 10616
rect 13624 10616 13652 10618
rect 13624 10584 13680 10616
rect 13714 10584 13773 10618
rect 13079 10550 13773 10584
rect 13079 10528 13152 10550
rect 13186 10528 13252 10550
rect 13286 10528 13352 10550
rect 13386 10528 13452 10550
rect 13079 10494 13140 10528
rect 13186 10516 13230 10528
rect 13286 10516 13320 10528
rect 13386 10516 13410 10528
rect 13174 10494 13230 10516
rect 13264 10494 13320 10516
rect 13354 10494 13410 10516
rect 13444 10516 13452 10528
rect 13486 10528 13552 10550
rect 13486 10516 13500 10528
rect 13444 10494 13500 10516
rect 13534 10516 13552 10528
rect 13586 10528 13652 10550
rect 13686 10528 13773 10550
rect 13586 10516 13590 10528
rect 13534 10494 13590 10516
rect 13624 10516 13652 10528
rect 13624 10494 13680 10516
rect 13714 10494 13773 10528
rect 13079 10450 13773 10494
rect 13079 10438 13152 10450
rect 13186 10438 13252 10450
rect 13286 10438 13352 10450
rect 13386 10438 13452 10450
rect 13079 10404 13140 10438
rect 13186 10416 13230 10438
rect 13286 10416 13320 10438
rect 13386 10416 13410 10438
rect 13174 10404 13230 10416
rect 13264 10404 13320 10416
rect 13354 10404 13410 10416
rect 13444 10416 13452 10438
rect 13486 10438 13552 10450
rect 13486 10416 13500 10438
rect 13444 10404 13500 10416
rect 13534 10416 13552 10438
rect 13586 10438 13652 10450
rect 13686 10438 13773 10450
rect 13586 10416 13590 10438
rect 13534 10404 13590 10416
rect 13624 10416 13652 10438
rect 13624 10404 13680 10416
rect 13714 10404 13773 10438
rect 13079 10343 13773 10404
rect 13835 10986 13907 11042
rect 13835 10952 13854 10986
rect 13888 10952 13907 10986
rect 13835 10896 13907 10952
rect 13835 10862 13854 10896
rect 13888 10862 13907 10896
rect 13835 10806 13907 10862
rect 13835 10772 13854 10806
rect 13888 10772 13907 10806
rect 13835 10716 13907 10772
rect 13835 10682 13854 10716
rect 13888 10682 13907 10716
rect 13835 10626 13907 10682
rect 13835 10592 13854 10626
rect 13888 10592 13907 10626
rect 13835 10536 13907 10592
rect 13835 10502 13854 10536
rect 13888 10502 13907 10536
rect 13835 10446 13907 10502
rect 13835 10412 13854 10446
rect 13888 10412 13907 10446
rect 13835 10356 13907 10412
rect 12945 10290 13017 10341
rect 13835 10322 13854 10356
rect 13888 10322 13907 10356
rect 13835 10290 13907 10322
rect 12945 10262 13907 10290
rect 12945 10228 13042 10262
rect 13076 10228 13132 10262
rect 13166 10228 13222 10262
rect 13256 10228 13312 10262
rect 13346 10228 13402 10262
rect 13436 10228 13492 10262
rect 13526 10228 13582 10262
rect 13616 10228 13672 10262
rect 13706 10228 13762 10262
rect 13796 10228 13907 10262
rect 12945 10209 13907 10228
rect 13971 11152 14003 11186
rect 14037 11152 14070 11186
rect 13971 11096 14070 11152
rect 13971 11062 14003 11096
rect 14037 11062 14070 11096
rect 13971 11006 14070 11062
rect 13971 10972 14003 11006
rect 14037 10972 14070 11006
rect 13971 10916 14070 10972
rect 13971 10882 14003 10916
rect 14037 10882 14070 10916
rect 13971 10826 14070 10882
rect 13971 10792 14003 10826
rect 14037 10792 14070 10826
rect 13971 10736 14070 10792
rect 13971 10702 14003 10736
rect 14037 10702 14070 10736
rect 13971 10646 14070 10702
rect 13971 10612 14003 10646
rect 14037 10612 14070 10646
rect 13971 10556 14070 10612
rect 13971 10522 14003 10556
rect 14037 10522 14070 10556
rect 13971 10466 14070 10522
rect 13971 10432 14003 10466
rect 14037 10432 14070 10466
rect 13971 10376 14070 10432
rect 13971 10342 14003 10376
rect 14037 10342 14070 10376
rect 13971 10286 14070 10342
rect 13971 10252 14003 10286
rect 14037 10252 14070 10286
rect 12756 10162 12816 10196
rect 12850 10162 12881 10196
rect 12756 10145 12881 10162
rect 12946 10145 13906 10209
rect 13971 10196 14070 10252
rect 13971 10162 14003 10196
rect 14037 10162 14070 10196
rect 13971 10145 14070 10162
rect 12756 10112 14070 10145
rect 12756 10078 12912 10112
rect 12946 10078 13002 10112
rect 13036 10078 13092 10112
rect 13126 10078 13182 10112
rect 13216 10078 13272 10112
rect 13306 10078 13362 10112
rect 13396 10078 13452 10112
rect 13486 10078 13542 10112
rect 13576 10078 13632 10112
rect 13666 10078 13722 10112
rect 13756 10078 13812 10112
rect 13846 10078 13902 10112
rect 13936 10078 14070 10112
rect 12756 10046 14070 10078
rect 17204 11362 17238 11432
rect 14820 11294 14854 11328
rect 15000 11294 15041 11328
rect 15085 11294 15109 11328
rect 15157 11294 15177 11328
rect 15229 11294 15245 11328
rect 15301 11294 15313 11328
rect 15373 11294 15381 11328
rect 15445 11294 15449 11328
rect 15551 11294 15555 11328
rect 15619 11294 15627 11328
rect 15687 11294 15699 11328
rect 15755 11294 15771 11328
rect 15823 11294 15843 11328
rect 15891 11294 15915 11328
rect 15959 11294 16000 11328
rect 16058 11294 16099 11328
rect 16143 11294 16167 11328
rect 16215 11294 16235 11328
rect 16287 11294 16303 11328
rect 16359 11294 16371 11328
rect 16431 11294 16439 11328
rect 16503 11294 16507 11328
rect 16609 11294 16613 11328
rect 16677 11294 16685 11328
rect 16745 11294 16757 11328
rect 16813 11294 16829 11328
rect 16881 11294 16901 11328
rect 16949 11294 16973 11328
rect 17017 11294 17058 11328
rect 17204 11294 17238 11328
rect 14820 11226 14854 11260
rect 14820 11158 14854 11192
rect 14820 11090 14854 11124
rect 14820 11022 14854 11056
rect 14820 10954 14854 10988
rect 14820 10886 14854 10920
rect 14820 10818 14854 10852
rect 14820 10750 14854 10784
rect 14820 10682 14854 10716
rect 14820 10614 14854 10648
rect 14820 10546 14854 10580
rect 14820 10478 14854 10512
rect 14820 10410 14854 10444
rect 14820 10342 14854 10376
rect 14820 10274 14854 10308
rect 14820 10206 14854 10240
rect 14820 10138 14854 10172
rect 14820 10070 14854 10104
rect 12756 9844 12871 10046
rect 12946 10040 13906 10046
rect 14820 10002 14854 10036
rect 14820 9934 14854 9968
rect 14820 9866 14854 9900
rect 12756 9809 14070 9844
rect 12756 9786 12912 9809
rect 12756 9752 12816 9786
rect 12850 9775 12912 9786
rect 12946 9775 13002 9809
rect 13036 9775 13092 9809
rect 13126 9775 13182 9809
rect 13216 9775 13272 9809
rect 13306 9775 13362 9809
rect 13396 9775 13452 9809
rect 13486 9775 13542 9809
rect 13576 9775 13632 9809
rect 13666 9775 13722 9809
rect 13756 9775 13812 9809
rect 13846 9775 13902 9809
rect 13936 9786 14070 9809
rect 13936 9775 14003 9786
rect 12850 9752 14003 9775
rect 14037 9752 14070 9786
rect 12756 9745 14070 9752
rect 12756 9696 12881 9745
rect 12756 9662 12816 9696
rect 12850 9662 12881 9696
rect 13971 9696 14070 9745
rect 12756 9606 12881 9662
rect 12756 9572 12816 9606
rect 12850 9572 12881 9606
rect 12756 9516 12881 9572
rect 12756 9482 12816 9516
rect 12850 9482 12881 9516
rect 12756 9426 12881 9482
rect 12756 9392 12816 9426
rect 12850 9392 12881 9426
rect 12756 9336 12881 9392
rect 12756 9302 12816 9336
rect 12850 9302 12881 9336
rect 12756 9246 12881 9302
rect 12756 9212 12816 9246
rect 12850 9212 12881 9246
rect 12756 9156 12881 9212
rect 12756 9122 12816 9156
rect 12850 9122 12881 9156
rect 12756 9066 12881 9122
rect 12756 9032 12816 9066
rect 12850 9032 12881 9066
rect 12756 8976 12881 9032
rect 12756 8942 12816 8976
rect 12850 8942 12881 8976
rect 12756 8886 12881 8942
rect 12756 8852 12816 8886
rect 12850 8852 12881 8886
rect 12756 8796 12881 8852
rect 12756 8762 12816 8796
rect 12850 8762 12881 8796
rect 12756 8706 12881 8762
rect 12945 9662 13907 9681
rect 12945 9628 13076 9662
rect 13110 9628 13166 9662
rect 13200 9628 13256 9662
rect 13290 9628 13346 9662
rect 13380 9628 13436 9662
rect 13470 9628 13526 9662
rect 13560 9628 13616 9662
rect 13650 9628 13706 9662
rect 13740 9628 13796 9662
rect 13830 9628 13907 9662
rect 12945 9609 13907 9628
rect 12945 9605 13017 9609
rect 12945 9571 12964 9605
rect 12998 9571 13017 9605
rect 12945 9515 13017 9571
rect 13835 9586 13907 9609
rect 13835 9552 13854 9586
rect 13888 9552 13907 9586
rect 12945 9481 12964 9515
rect 12998 9481 13017 9515
rect 12945 9425 13017 9481
rect 12945 9391 12964 9425
rect 12998 9391 13017 9425
rect 12945 9335 13017 9391
rect 12945 9301 12964 9335
rect 12998 9301 13017 9335
rect 12945 9245 13017 9301
rect 12945 9211 12964 9245
rect 12998 9211 13017 9245
rect 12945 9155 13017 9211
rect 12945 9121 12964 9155
rect 12998 9121 13017 9155
rect 12945 9065 13017 9121
rect 12945 9031 12964 9065
rect 12998 9031 13017 9065
rect 12945 8975 13017 9031
rect 12945 8941 12964 8975
rect 12998 8941 13017 8975
rect 12945 8885 13017 8941
rect 12945 8851 12964 8885
rect 12998 8851 13017 8885
rect 13079 9488 13773 9547
rect 13079 9454 13140 9488
rect 13174 9460 13230 9488
rect 13264 9460 13320 9488
rect 13354 9460 13410 9488
rect 13186 9454 13230 9460
rect 13286 9454 13320 9460
rect 13386 9454 13410 9460
rect 13444 9460 13500 9488
rect 13444 9454 13452 9460
rect 13079 9426 13152 9454
rect 13186 9426 13252 9454
rect 13286 9426 13352 9454
rect 13386 9426 13452 9454
rect 13486 9454 13500 9460
rect 13534 9460 13590 9488
rect 13534 9454 13552 9460
rect 13486 9426 13552 9454
rect 13586 9454 13590 9460
rect 13624 9460 13680 9488
rect 13624 9454 13652 9460
rect 13714 9454 13773 9488
rect 13586 9426 13652 9454
rect 13686 9426 13773 9454
rect 13079 9398 13773 9426
rect 13079 9364 13140 9398
rect 13174 9364 13230 9398
rect 13264 9364 13320 9398
rect 13354 9364 13410 9398
rect 13444 9364 13500 9398
rect 13534 9364 13590 9398
rect 13624 9364 13680 9398
rect 13714 9364 13773 9398
rect 13079 9360 13773 9364
rect 13079 9326 13152 9360
rect 13186 9326 13252 9360
rect 13286 9326 13352 9360
rect 13386 9326 13452 9360
rect 13486 9326 13552 9360
rect 13586 9326 13652 9360
rect 13686 9326 13773 9360
rect 13079 9308 13773 9326
rect 13079 9274 13140 9308
rect 13174 9274 13230 9308
rect 13264 9274 13320 9308
rect 13354 9274 13410 9308
rect 13444 9274 13500 9308
rect 13534 9274 13590 9308
rect 13624 9274 13680 9308
rect 13714 9274 13773 9308
rect 13079 9260 13773 9274
rect 13079 9226 13152 9260
rect 13186 9226 13252 9260
rect 13286 9226 13352 9260
rect 13386 9226 13452 9260
rect 13486 9226 13552 9260
rect 13586 9226 13652 9260
rect 13686 9226 13773 9260
rect 13079 9218 13773 9226
rect 13079 9184 13140 9218
rect 13174 9184 13230 9218
rect 13264 9184 13320 9218
rect 13354 9184 13410 9218
rect 13444 9184 13500 9218
rect 13534 9184 13590 9218
rect 13624 9184 13680 9218
rect 13714 9184 13773 9218
rect 13079 9160 13773 9184
rect 13079 9128 13152 9160
rect 13186 9128 13252 9160
rect 13286 9128 13352 9160
rect 13386 9128 13452 9160
rect 13079 9094 13140 9128
rect 13186 9126 13230 9128
rect 13286 9126 13320 9128
rect 13386 9126 13410 9128
rect 13174 9094 13230 9126
rect 13264 9094 13320 9126
rect 13354 9094 13410 9126
rect 13444 9126 13452 9128
rect 13486 9128 13552 9160
rect 13486 9126 13500 9128
rect 13444 9094 13500 9126
rect 13534 9126 13552 9128
rect 13586 9128 13652 9160
rect 13686 9128 13773 9160
rect 13586 9126 13590 9128
rect 13534 9094 13590 9126
rect 13624 9126 13652 9128
rect 13624 9094 13680 9126
rect 13714 9094 13773 9128
rect 13079 9060 13773 9094
rect 13079 9038 13152 9060
rect 13186 9038 13252 9060
rect 13286 9038 13352 9060
rect 13386 9038 13452 9060
rect 13079 9004 13140 9038
rect 13186 9026 13230 9038
rect 13286 9026 13320 9038
rect 13386 9026 13410 9038
rect 13174 9004 13230 9026
rect 13264 9004 13320 9026
rect 13354 9004 13410 9026
rect 13444 9026 13452 9038
rect 13486 9038 13552 9060
rect 13486 9026 13500 9038
rect 13444 9004 13500 9026
rect 13534 9026 13552 9038
rect 13586 9038 13652 9060
rect 13686 9038 13773 9060
rect 13586 9026 13590 9038
rect 13534 9004 13590 9026
rect 13624 9026 13652 9038
rect 13624 9004 13680 9026
rect 13714 9004 13773 9038
rect 13079 8960 13773 9004
rect 13079 8948 13152 8960
rect 13186 8948 13252 8960
rect 13286 8948 13352 8960
rect 13386 8948 13452 8960
rect 13079 8914 13140 8948
rect 13186 8926 13230 8948
rect 13286 8926 13320 8948
rect 13386 8926 13410 8948
rect 13174 8914 13230 8926
rect 13264 8914 13320 8926
rect 13354 8914 13410 8926
rect 13444 8926 13452 8948
rect 13486 8948 13552 8960
rect 13486 8926 13500 8948
rect 13444 8914 13500 8926
rect 13534 8926 13552 8948
rect 13586 8948 13652 8960
rect 13686 8948 13773 8960
rect 13586 8926 13590 8948
rect 13534 8914 13590 8926
rect 13624 8926 13652 8948
rect 13624 8914 13680 8926
rect 13714 8914 13773 8948
rect 13079 8853 13773 8914
rect 13835 9496 13907 9552
rect 13835 9462 13854 9496
rect 13888 9462 13907 9496
rect 13835 9406 13907 9462
rect 13835 9372 13854 9406
rect 13888 9372 13907 9406
rect 13835 9316 13907 9372
rect 13835 9282 13854 9316
rect 13888 9282 13907 9316
rect 13835 9226 13907 9282
rect 13835 9192 13854 9226
rect 13888 9192 13907 9226
rect 13835 9136 13907 9192
rect 13835 9102 13854 9136
rect 13888 9102 13907 9136
rect 13835 9046 13907 9102
rect 13835 9012 13854 9046
rect 13888 9012 13907 9046
rect 13835 8956 13907 9012
rect 13835 8922 13854 8956
rect 13888 8922 13907 8956
rect 13835 8866 13907 8922
rect 12945 8800 13017 8851
rect 13835 8832 13854 8866
rect 13888 8832 13907 8866
rect 13835 8800 13907 8832
rect 12945 8772 13907 8800
rect 12945 8738 13042 8772
rect 13076 8738 13132 8772
rect 13166 8738 13222 8772
rect 13256 8738 13312 8772
rect 13346 8738 13402 8772
rect 13436 8738 13492 8772
rect 13526 8738 13582 8772
rect 13616 8738 13672 8772
rect 13706 8738 13762 8772
rect 13796 8738 13907 8772
rect 12945 8719 13907 8738
rect 13971 9662 14003 9696
rect 14037 9662 14070 9696
rect 13971 9606 14070 9662
rect 13971 9572 14003 9606
rect 14037 9572 14070 9606
rect 13971 9516 14070 9572
rect 13971 9482 14003 9516
rect 14037 9482 14070 9516
rect 13971 9426 14070 9482
rect 13971 9392 14003 9426
rect 14037 9392 14070 9426
rect 13971 9336 14070 9392
rect 13971 9302 14003 9336
rect 14037 9302 14070 9336
rect 13971 9246 14070 9302
rect 13971 9212 14003 9246
rect 14037 9212 14070 9246
rect 13971 9156 14070 9212
rect 13971 9122 14003 9156
rect 14037 9122 14070 9156
rect 13971 9066 14070 9122
rect 13971 9032 14003 9066
rect 14037 9032 14070 9066
rect 13971 8976 14070 9032
rect 13971 8942 14003 8976
rect 14037 8942 14070 8976
rect 13971 8886 14070 8942
rect 13971 8852 14003 8886
rect 14037 8852 14070 8886
rect 13971 8796 14070 8852
rect 13971 8762 14003 8796
rect 14037 8762 14070 8796
rect 12756 8672 12816 8706
rect 12850 8672 12881 8706
rect 12756 8655 12881 8672
rect 12946 8655 13906 8719
rect 13971 8706 14070 8762
rect 13971 8672 14003 8706
rect 14037 8672 14070 8706
rect 13971 8655 14070 8672
rect 12756 8622 14070 8655
rect 12756 8588 12912 8622
rect 12946 8588 13002 8622
rect 13036 8588 13092 8622
rect 13126 8588 13182 8622
rect 13216 8588 13272 8622
rect 13306 8588 13362 8622
rect 13396 8588 13452 8622
rect 13486 8588 13542 8622
rect 13576 8588 13632 8622
rect 13666 8588 13722 8622
rect 13756 8588 13812 8622
rect 13846 8588 13902 8622
rect 13936 8588 14070 8622
rect 12756 8556 14070 8588
rect 14820 9798 14854 9832
rect 14820 9730 14854 9764
rect 14820 9662 14854 9696
rect 14820 9594 14854 9628
rect 14820 9526 14854 9560
rect 14820 9458 14854 9492
rect 14820 9390 14854 9424
rect 14820 9322 14854 9356
rect 14820 9254 14854 9288
rect 14820 9186 14854 9220
rect 14820 9118 14854 9152
rect 14820 9050 14854 9084
rect 14820 8982 14854 9016
rect 14820 8914 14854 8948
rect 14820 8846 14854 8880
rect 14820 8778 14854 8812
rect 14820 8710 14854 8744
rect 14820 8642 14854 8676
rect 14820 8574 14854 8608
rect 12756 8434 12871 8556
rect 12946 8550 13906 8556
rect 14820 8506 14854 8540
rect 14820 8438 14854 8472
rect 12756 8399 14060 8434
rect 12756 8376 12902 8399
rect 12756 8342 12806 8376
rect 12840 8365 12902 8376
rect 12936 8365 12992 8399
rect 13026 8365 13082 8399
rect 13116 8365 13172 8399
rect 13206 8365 13262 8399
rect 13296 8365 13352 8399
rect 13386 8365 13442 8399
rect 13476 8365 13532 8399
rect 13566 8365 13622 8399
rect 13656 8365 13712 8399
rect 13746 8365 13802 8399
rect 13836 8365 13892 8399
rect 13926 8376 14060 8399
rect 13926 8365 13993 8376
rect 12840 8342 13993 8365
rect 14027 8342 14060 8376
rect -9108 8336 -9016 8337
rect -7984 7859 -3408 8337
rect -7984 7825 -7749 7859
rect -7715 7825 -7681 7859
rect -7647 7825 -7613 7859
rect -7579 7825 -7545 7859
rect -7511 7825 -7477 7859
rect -7443 7825 -7409 7859
rect -7375 7825 -7341 7859
rect -7307 7825 -7273 7859
rect -7239 7825 -7205 7859
rect -7171 7825 -7137 7859
rect -7103 7825 -7069 7859
rect -7035 7825 -7001 7859
rect -6967 7825 -6933 7859
rect -6899 7825 -6865 7859
rect -6831 7825 -6797 7859
rect -6763 7825 -6729 7859
rect -6695 7825 -6661 7859
rect -6627 7825 -6593 7859
rect -6559 7825 -6525 7859
rect -6491 7825 -6457 7859
rect -6423 7825 -6389 7859
rect -6355 7825 -6321 7859
rect -6287 7825 -6253 7859
rect -6219 7825 -6185 7859
rect -6151 7825 -6117 7859
rect -6083 7825 -6049 7859
rect -6015 7825 -5981 7859
rect -5947 7825 -5913 7859
rect -5879 7825 -5845 7859
rect -5811 7825 -5777 7859
rect -5743 7825 -5709 7859
rect -5675 7825 -5641 7859
rect -5607 7825 -5573 7859
rect -5539 7825 -5505 7859
rect -5471 7825 -5437 7859
rect -5403 7825 -5369 7859
rect -5335 7825 -5301 7859
rect -5267 7825 -5233 7859
rect -5199 7825 -5165 7859
rect -5131 7825 -5097 7859
rect -5063 7825 -5029 7859
rect -4995 7825 -4961 7859
rect -4927 7825 -4893 7859
rect -4859 7825 -4825 7859
rect -4791 7825 -4757 7859
rect -4723 7825 -4689 7859
rect -4655 7825 -4621 7859
rect -4587 7825 -4553 7859
rect -4519 7825 -4485 7859
rect -4451 7825 -4417 7859
rect -4383 7825 -4349 7859
rect -4315 7825 -4281 7859
rect -4247 7825 -4213 7859
rect -4179 7825 -4145 7859
rect -4111 7825 -4077 7859
rect -4043 7825 -4009 7859
rect -3975 7825 -3941 7859
rect -3907 7825 -3873 7859
rect -3839 7825 -3805 7859
rect -3771 7825 -3737 7859
rect -3703 7825 -3669 7859
rect -3635 7825 -3601 7859
rect -3567 7825 -3408 7859
rect -7984 7814 -3408 7825
rect -7984 7682 -7918 7814
rect -7984 7648 -7968 7682
rect -7934 7648 -7918 7682
rect -7984 7614 -7918 7648
rect -7984 7580 -7968 7614
rect -7934 7580 -7918 7614
rect -3470 7694 -3408 7814
rect -3470 7660 -3456 7694
rect -3422 7660 -3408 7694
rect -3470 7626 -3408 7660
rect -7984 7546 -7918 7580
rect -7734 7576 -7687 7610
rect -7651 7576 -7617 7610
rect -7581 7576 -7534 7610
rect -7476 7576 -7429 7610
rect -7393 7576 -7359 7610
rect -7323 7576 -7276 7610
rect -7218 7576 -7171 7610
rect -7135 7576 -7101 7610
rect -7065 7576 -7018 7610
rect -6960 7576 -6913 7610
rect -6877 7576 -6843 7610
rect -6807 7576 -6760 7610
rect -6702 7576 -6655 7610
rect -6619 7576 -6585 7610
rect -6549 7576 -6502 7610
rect -6444 7576 -6397 7610
rect -6361 7576 -6327 7610
rect -6291 7576 -6244 7610
rect -6186 7576 -6139 7610
rect -6103 7576 -6069 7610
rect -6033 7576 -5986 7610
rect -5928 7576 -5881 7610
rect -5845 7576 -5811 7610
rect -5775 7576 -5728 7610
rect -5670 7576 -5623 7610
rect -5587 7576 -5553 7610
rect -5517 7576 -5470 7610
rect -5412 7576 -5365 7610
rect -5329 7576 -5295 7610
rect -5259 7576 -5212 7610
rect -5154 7576 -5107 7610
rect -5071 7576 -5037 7610
rect -5001 7576 -4954 7610
rect -4896 7576 -4849 7610
rect -4813 7576 -4779 7610
rect -4743 7576 -4696 7610
rect -4638 7576 -4591 7610
rect -4555 7576 -4521 7610
rect -4485 7576 -4438 7610
rect -4380 7576 -4333 7610
rect -4297 7576 -4263 7610
rect -4227 7576 -4180 7610
rect -4122 7576 -4075 7610
rect -4039 7576 -4005 7610
rect -3969 7576 -3922 7610
rect -3864 7576 -3817 7610
rect -3781 7576 -3747 7610
rect -3711 7576 -3664 7610
rect -3470 7592 -3456 7626
rect -3422 7592 -3408 7626
rect -7984 7512 -7968 7546
rect -7934 7512 -7918 7546
rect -3470 7558 -3408 7592
rect -7984 7478 -7918 7512
rect -7984 7444 -7968 7478
rect -7934 7444 -7918 7478
rect -7984 7410 -7918 7444
rect -7984 7376 -7968 7410
rect -7934 7376 -7918 7410
rect -7984 7342 -7918 7376
rect -7984 7308 -7968 7342
rect -7934 7308 -7918 7342
rect -7984 7274 -7918 7308
rect -7984 7240 -7968 7274
rect -7934 7240 -7918 7274
rect -7984 7206 -7918 7240
rect -7984 7172 -7968 7206
rect -7934 7172 -7918 7206
rect -7984 7138 -7918 7172
rect -7984 7104 -7968 7138
rect -7934 7104 -7918 7138
rect -7984 7070 -7918 7104
rect -7984 7036 -7968 7070
rect -7934 7036 -7918 7070
rect -7984 7002 -7918 7036
rect -7984 6968 -7968 7002
rect -7934 6968 -7918 7002
rect -7984 6934 -7918 6968
rect -7984 6900 -7968 6934
rect -7934 6900 -7918 6934
rect -7984 6866 -7918 6900
rect -7984 6832 -7968 6866
rect -7934 6832 -7918 6866
rect -7984 6798 -7918 6832
rect -7984 6764 -7968 6798
rect -7934 6764 -7918 6798
rect -7984 6730 -7918 6764
rect -7984 6696 -7968 6730
rect -7934 6696 -7918 6730
rect -7984 6662 -7918 6696
rect -7984 6628 -7968 6662
rect -7934 6628 -7918 6662
rect -7984 6594 -7918 6628
rect -7984 6560 -7968 6594
rect -7934 6560 -7918 6594
rect -7984 6526 -7918 6560
rect -7984 6492 -7968 6526
rect -7934 6492 -7918 6526
rect -7984 6458 -7918 6492
rect -7984 6424 -7968 6458
rect -7934 6424 -7918 6458
rect -7984 6390 -7918 6424
rect -7984 6356 -7968 6390
rect -7934 6356 -7918 6390
rect -7984 6322 -7918 6356
rect -7984 6288 -7968 6322
rect -7934 6288 -7918 6322
rect -7984 6254 -7918 6288
rect -7984 6220 -7968 6254
rect -7934 6220 -7918 6254
rect -7984 6186 -7918 6220
rect -7984 6152 -7968 6186
rect -7934 6152 -7918 6186
rect -7984 6118 -7918 6152
rect -7984 6084 -7968 6118
rect -7934 6084 -7918 6118
rect -7984 6050 -7918 6084
rect -7984 6016 -7968 6050
rect -7934 6016 -7918 6050
rect -7984 5982 -7918 6016
rect -7984 5948 -7968 5982
rect -7934 5948 -7918 5982
rect -7984 5914 -7918 5948
rect -7984 5886 -7968 5914
rect -7984 5852 -7969 5886
rect -7934 5880 -7918 5914
rect -7935 5852 -7918 5880
rect -7984 5846 -7918 5852
rect -7984 5814 -7968 5846
rect -7984 5780 -7969 5814
rect -7934 5812 -7918 5846
rect -7935 5780 -7918 5812
rect -7984 5778 -7918 5780
rect -7984 5744 -7968 5778
rect -7934 5744 -7918 5778
rect -7984 5742 -7918 5744
rect -7984 5708 -7969 5742
rect -7935 5710 -7918 5742
rect -7984 5676 -7968 5708
rect -7934 5676 -7918 5710
rect -7984 5642 -7918 5676
rect -7984 5608 -7968 5642
rect -7934 5608 -7918 5642
rect -7984 5574 -7918 5608
rect -7984 5540 -7968 5574
rect -7934 5540 -7918 5574
rect -7984 5506 -7918 5540
rect -7780 7507 -7746 7542
rect -7780 7439 -7746 7457
rect -7780 7371 -7746 7385
rect -7780 7303 -7746 7313
rect -7780 7235 -7746 7241
rect -7780 7167 -7746 7169
rect -7780 7131 -7746 7133
rect -7780 7059 -7746 7065
rect -7780 6987 -7746 6997
rect -7780 6915 -7746 6929
rect -7780 6843 -7746 6861
rect -7780 6771 -7746 6793
rect -7780 6699 -7746 6725
rect -7780 6627 -7746 6657
rect -7780 6555 -7746 6589
rect -7780 6487 -7746 6521
rect -7780 6419 -7746 6449
rect -7780 6351 -7746 6377
rect -7780 6283 -7746 6305
rect -7780 6215 -7746 6233
rect -7780 6147 -7746 6161
rect -7780 6079 -7746 6089
rect -7780 6011 -7746 6017
rect -7780 5943 -7746 5945
rect -7780 5907 -7746 5909
rect -7780 5835 -7746 5841
rect -7780 5763 -7746 5773
rect -7780 5691 -7746 5705
rect -7780 5619 -7746 5637
rect -7780 5534 -7746 5569
rect -7522 7507 -7488 7542
rect -7522 7439 -7488 7457
rect -7522 7371 -7488 7385
rect -7522 7303 -7488 7313
rect -7522 7235 -7488 7241
rect -7522 7167 -7488 7169
rect -7522 7131 -7488 7133
rect -7522 7059 -7488 7065
rect -7522 6987 -7488 6997
rect -7522 6915 -7488 6929
rect -7522 6843 -7488 6861
rect -7522 6771 -7488 6793
rect -7522 6699 -7488 6725
rect -7522 6627 -7488 6657
rect -7522 6555 -7488 6589
rect -7522 6487 -7488 6521
rect -7522 6419 -7488 6449
rect -7522 6351 -7488 6377
rect -7522 6283 -7488 6305
rect -7522 6215 -7488 6233
rect -7522 6147 -7488 6161
rect -7522 6079 -7488 6089
rect -7522 6011 -7488 6017
rect -7522 5943 -7488 5945
rect -7522 5907 -7488 5909
rect -7522 5835 -7488 5841
rect -7522 5763 -7488 5773
rect -7522 5691 -7488 5705
rect -7522 5619 -7488 5637
rect -7522 5534 -7488 5569
rect -7264 7507 -7230 7542
rect -7264 7439 -7230 7457
rect -7264 7371 -7230 7385
rect -7264 7303 -7230 7313
rect -7264 7235 -7230 7241
rect -7264 7167 -7230 7169
rect -7264 7131 -7230 7133
rect -7264 7059 -7230 7065
rect -7264 6987 -7230 6997
rect -7264 6915 -7230 6929
rect -7264 6843 -7230 6861
rect -7264 6771 -7230 6793
rect -7264 6699 -7230 6725
rect -7264 6627 -7230 6657
rect -7264 6555 -7230 6589
rect -7264 6487 -7230 6521
rect -7264 6419 -7230 6449
rect -7264 6351 -7230 6377
rect -7264 6283 -7230 6305
rect -7264 6215 -7230 6233
rect -7264 6147 -7230 6161
rect -7264 6079 -7230 6089
rect -7264 6011 -7230 6017
rect -7264 5943 -7230 5945
rect -7264 5907 -7230 5909
rect -7264 5835 -7230 5841
rect -7264 5763 -7230 5773
rect -7264 5691 -7230 5705
rect -7264 5619 -7230 5637
rect -7264 5534 -7230 5569
rect -7006 7507 -6972 7542
rect -7006 7439 -6972 7457
rect -7006 7371 -6972 7385
rect -7006 7303 -6972 7313
rect -7006 7235 -6972 7241
rect -7006 7167 -6972 7169
rect -7006 7131 -6972 7133
rect -7006 7059 -6972 7065
rect -7006 6987 -6972 6997
rect -7006 6915 -6972 6929
rect -7006 6843 -6972 6861
rect -7006 6771 -6972 6793
rect -7006 6699 -6972 6725
rect -7006 6627 -6972 6657
rect -7006 6555 -6972 6589
rect -7006 6487 -6972 6521
rect -7006 6419 -6972 6449
rect -7006 6351 -6972 6377
rect -7006 6283 -6972 6305
rect -7006 6215 -6972 6233
rect -7006 6147 -6972 6161
rect -7006 6079 -6972 6089
rect -7006 6011 -6972 6017
rect -7006 5943 -6972 5945
rect -7006 5907 -6972 5909
rect -7006 5835 -6972 5841
rect -7006 5763 -6972 5773
rect -7006 5691 -6972 5705
rect -7006 5619 -6972 5637
rect -7006 5534 -6972 5569
rect -6748 7507 -6714 7542
rect -6748 7439 -6714 7457
rect -6748 7371 -6714 7385
rect -6748 7303 -6714 7313
rect -6748 7235 -6714 7241
rect -6748 7167 -6714 7169
rect -6748 7131 -6714 7133
rect -6748 7059 -6714 7065
rect -6748 6987 -6714 6997
rect -6748 6915 -6714 6929
rect -6748 6843 -6714 6861
rect -6748 6771 -6714 6793
rect -6748 6699 -6714 6725
rect -6748 6627 -6714 6657
rect -6748 6555 -6714 6589
rect -6748 6487 -6714 6521
rect -6748 6419 -6714 6449
rect -6748 6351 -6714 6377
rect -6748 6283 -6714 6305
rect -6748 6215 -6714 6233
rect -6748 6147 -6714 6161
rect -6748 6079 -6714 6089
rect -6748 6011 -6714 6017
rect -6748 5943 -6714 5945
rect -6748 5907 -6714 5909
rect -6748 5835 -6714 5841
rect -6748 5763 -6714 5773
rect -6748 5691 -6714 5705
rect -6748 5619 -6714 5637
rect -6748 5534 -6714 5569
rect -6490 7507 -6456 7542
rect -6490 7439 -6456 7457
rect -6490 7371 -6456 7385
rect -6490 7303 -6456 7313
rect -6490 7235 -6456 7241
rect -6490 7167 -6456 7169
rect -6490 7131 -6456 7133
rect -6490 7059 -6456 7065
rect -6490 6987 -6456 6997
rect -6490 6915 -6456 6929
rect -6490 6843 -6456 6861
rect -6490 6771 -6456 6793
rect -6490 6699 -6456 6725
rect -6490 6627 -6456 6657
rect -6490 6555 -6456 6589
rect -6490 6487 -6456 6521
rect -6490 6419 -6456 6449
rect -6490 6351 -6456 6377
rect -6490 6283 -6456 6305
rect -6490 6215 -6456 6233
rect -6490 6147 -6456 6161
rect -6490 6079 -6456 6089
rect -6490 6011 -6456 6017
rect -6490 5943 -6456 5945
rect -6490 5907 -6456 5909
rect -6490 5835 -6456 5841
rect -6490 5763 -6456 5773
rect -6490 5691 -6456 5705
rect -6490 5619 -6456 5637
rect -6490 5534 -6456 5569
rect -6232 7507 -6198 7542
rect -6232 7439 -6198 7457
rect -6232 7371 -6198 7385
rect -6232 7303 -6198 7313
rect -6232 7235 -6198 7241
rect -6232 7167 -6198 7169
rect -6232 7131 -6198 7133
rect -6232 7059 -6198 7065
rect -6232 6987 -6198 6997
rect -6232 6915 -6198 6929
rect -6232 6843 -6198 6861
rect -6232 6771 -6198 6793
rect -6232 6699 -6198 6725
rect -6232 6627 -6198 6657
rect -6232 6555 -6198 6589
rect -6232 6487 -6198 6521
rect -6232 6419 -6198 6449
rect -6232 6351 -6198 6377
rect -6232 6283 -6198 6305
rect -6232 6215 -6198 6233
rect -6232 6147 -6198 6161
rect -6232 6079 -6198 6089
rect -6232 6011 -6198 6017
rect -6232 5943 -6198 5945
rect -6232 5907 -6198 5909
rect -6232 5835 -6198 5841
rect -6232 5763 -6198 5773
rect -6232 5691 -6198 5705
rect -6232 5619 -6198 5637
rect -6232 5534 -6198 5569
rect -5974 7507 -5940 7542
rect -5974 7439 -5940 7457
rect -5974 7371 -5940 7385
rect -5974 7303 -5940 7313
rect -5974 7235 -5940 7241
rect -5974 7167 -5940 7169
rect -5974 7131 -5940 7133
rect -5974 7059 -5940 7065
rect -5974 6987 -5940 6997
rect -5974 6915 -5940 6929
rect -5974 6843 -5940 6861
rect -5974 6771 -5940 6793
rect -5974 6699 -5940 6725
rect -5974 6627 -5940 6657
rect -5974 6555 -5940 6589
rect -5974 6487 -5940 6521
rect -5974 6419 -5940 6449
rect -5974 6351 -5940 6377
rect -5974 6283 -5940 6305
rect -5974 6215 -5940 6233
rect -5974 6147 -5940 6161
rect -5974 6079 -5940 6089
rect -5974 6011 -5940 6017
rect -5974 5943 -5940 5945
rect -5974 5907 -5940 5909
rect -5974 5835 -5940 5841
rect -5974 5763 -5940 5773
rect -5974 5691 -5940 5705
rect -5974 5619 -5940 5637
rect -5974 5534 -5940 5569
rect -5716 7507 -5682 7542
rect -5716 7439 -5682 7457
rect -5716 7371 -5682 7385
rect -5716 7303 -5682 7313
rect -5716 7235 -5682 7241
rect -5716 7167 -5682 7169
rect -5716 7131 -5682 7133
rect -5716 7059 -5682 7065
rect -5716 6987 -5682 6997
rect -5716 6915 -5682 6929
rect -5716 6843 -5682 6861
rect -5716 6771 -5682 6793
rect -5716 6699 -5682 6725
rect -5716 6627 -5682 6657
rect -5716 6555 -5682 6589
rect -5716 6487 -5682 6521
rect -5716 6419 -5682 6449
rect -5716 6351 -5682 6377
rect -5716 6283 -5682 6305
rect -5716 6215 -5682 6233
rect -5716 6147 -5682 6161
rect -5716 6079 -5682 6089
rect -5716 6011 -5682 6017
rect -5716 5943 -5682 5945
rect -5716 5907 -5682 5909
rect -5716 5835 -5682 5841
rect -5716 5763 -5682 5773
rect -5716 5691 -5682 5705
rect -5716 5619 -5682 5637
rect -5716 5534 -5682 5569
rect -5458 7507 -5424 7542
rect -5458 7439 -5424 7457
rect -5458 7371 -5424 7385
rect -5458 7303 -5424 7313
rect -5458 7235 -5424 7241
rect -5458 7167 -5424 7169
rect -5458 7131 -5424 7133
rect -5458 7059 -5424 7065
rect -5458 6987 -5424 6997
rect -5458 6915 -5424 6929
rect -5458 6843 -5424 6861
rect -5458 6771 -5424 6793
rect -5458 6699 -5424 6725
rect -5458 6627 -5424 6657
rect -5458 6555 -5424 6589
rect -5458 6487 -5424 6521
rect -5458 6419 -5424 6449
rect -5458 6351 -5424 6377
rect -5458 6283 -5424 6305
rect -5458 6215 -5424 6233
rect -5458 6147 -5424 6161
rect -5458 6079 -5424 6089
rect -5458 6011 -5424 6017
rect -5458 5943 -5424 5945
rect -5458 5907 -5424 5909
rect -5458 5835 -5424 5841
rect -5458 5763 -5424 5773
rect -5458 5691 -5424 5705
rect -5458 5619 -5424 5637
rect -5458 5534 -5424 5569
rect -5200 7507 -5166 7542
rect -5200 7439 -5166 7457
rect -5200 7371 -5166 7385
rect -5200 7303 -5166 7313
rect -5200 7235 -5166 7241
rect -5200 7167 -5166 7169
rect -5200 7131 -5166 7133
rect -5200 7059 -5166 7065
rect -5200 6987 -5166 6997
rect -5200 6915 -5166 6929
rect -5200 6843 -5166 6861
rect -5200 6771 -5166 6793
rect -5200 6699 -5166 6725
rect -5200 6627 -5166 6657
rect -5200 6555 -5166 6589
rect -5200 6487 -5166 6521
rect -5200 6419 -5166 6449
rect -5200 6351 -5166 6377
rect -5200 6283 -5166 6305
rect -5200 6215 -5166 6233
rect -5200 6147 -5166 6161
rect -5200 6079 -5166 6089
rect -5200 6011 -5166 6017
rect -5200 5943 -5166 5945
rect -5200 5907 -5166 5909
rect -5200 5835 -5166 5841
rect -5200 5763 -5166 5773
rect -5200 5691 -5166 5705
rect -5200 5619 -5166 5637
rect -5200 5534 -5166 5569
rect -4942 7507 -4908 7542
rect -4942 7439 -4908 7457
rect -4942 7371 -4908 7385
rect -4942 7303 -4908 7313
rect -4942 7235 -4908 7241
rect -4942 7167 -4908 7169
rect -4942 7131 -4908 7133
rect -4942 7059 -4908 7065
rect -4942 6987 -4908 6997
rect -4942 6915 -4908 6929
rect -4942 6843 -4908 6861
rect -4942 6771 -4908 6793
rect -4942 6699 -4908 6725
rect -4942 6627 -4908 6657
rect -4942 6555 -4908 6589
rect -4942 6487 -4908 6521
rect -4942 6419 -4908 6449
rect -4942 6351 -4908 6377
rect -4942 6283 -4908 6305
rect -4942 6215 -4908 6233
rect -4942 6147 -4908 6161
rect -4942 6079 -4908 6089
rect -4942 6011 -4908 6017
rect -4942 5943 -4908 5945
rect -4942 5907 -4908 5909
rect -4942 5835 -4908 5841
rect -4942 5763 -4908 5773
rect -4942 5691 -4908 5705
rect -4942 5619 -4908 5637
rect -4942 5534 -4908 5569
rect -4684 7507 -4650 7542
rect -4684 7439 -4650 7457
rect -4684 7371 -4650 7385
rect -4684 7303 -4650 7313
rect -4684 7235 -4650 7241
rect -4684 7167 -4650 7169
rect -4684 7131 -4650 7133
rect -4684 7059 -4650 7065
rect -4684 6987 -4650 6997
rect -4684 6915 -4650 6929
rect -4684 6843 -4650 6861
rect -4684 6771 -4650 6793
rect -4684 6699 -4650 6725
rect -4684 6627 -4650 6657
rect -4684 6555 -4650 6589
rect -4684 6487 -4650 6521
rect -4684 6419 -4650 6449
rect -4684 6351 -4650 6377
rect -4684 6283 -4650 6305
rect -4684 6215 -4650 6233
rect -4684 6147 -4650 6161
rect -4684 6079 -4650 6089
rect -4684 6011 -4650 6017
rect -4684 5943 -4650 5945
rect -4684 5907 -4650 5909
rect -4684 5835 -4650 5841
rect -4684 5763 -4650 5773
rect -4684 5691 -4650 5705
rect -4684 5619 -4650 5637
rect -4684 5534 -4650 5569
rect -4426 7507 -4392 7542
rect -4426 7439 -4392 7457
rect -4426 7371 -4392 7385
rect -4426 7303 -4392 7313
rect -4426 7235 -4392 7241
rect -4426 7167 -4392 7169
rect -4426 7131 -4392 7133
rect -4426 7059 -4392 7065
rect -4426 6987 -4392 6997
rect -4426 6915 -4392 6929
rect -4426 6843 -4392 6861
rect -4426 6771 -4392 6793
rect -4426 6699 -4392 6725
rect -4426 6627 -4392 6657
rect -4426 6555 -4392 6589
rect -4426 6487 -4392 6521
rect -4426 6419 -4392 6449
rect -4426 6351 -4392 6377
rect -4426 6283 -4392 6305
rect -4426 6215 -4392 6233
rect -4426 6147 -4392 6161
rect -4426 6079 -4392 6089
rect -4426 6011 -4392 6017
rect -4426 5943 -4392 5945
rect -4426 5907 -4392 5909
rect -4426 5835 -4392 5841
rect -4426 5763 -4392 5773
rect -4426 5691 -4392 5705
rect -4426 5619 -4392 5637
rect -4426 5534 -4392 5569
rect -4168 7507 -4134 7542
rect -4168 7439 -4134 7457
rect -4168 7371 -4134 7385
rect -4168 7303 -4134 7313
rect -4168 7235 -4134 7241
rect -4168 7167 -4134 7169
rect -4168 7131 -4134 7133
rect -4168 7059 -4134 7065
rect -4168 6987 -4134 6997
rect -4168 6915 -4134 6929
rect -4168 6843 -4134 6861
rect -4168 6771 -4134 6793
rect -4168 6699 -4134 6725
rect -4168 6627 -4134 6657
rect -4168 6555 -4134 6589
rect -4168 6487 -4134 6521
rect -4168 6419 -4134 6449
rect -4168 6351 -4134 6377
rect -4168 6283 -4134 6305
rect -4168 6215 -4134 6233
rect -4168 6147 -4134 6161
rect -4168 6079 -4134 6089
rect -4168 6011 -4134 6017
rect -4168 5943 -4134 5945
rect -4168 5907 -4134 5909
rect -4168 5835 -4134 5841
rect -4168 5763 -4134 5773
rect -4168 5691 -4134 5705
rect -4168 5619 -4134 5637
rect -4168 5534 -4134 5569
rect -3910 7507 -3876 7542
rect -3910 7439 -3876 7457
rect -3910 7371 -3876 7385
rect -3910 7303 -3876 7313
rect -3910 7235 -3876 7241
rect -3910 7167 -3876 7169
rect -3910 7131 -3876 7133
rect -3910 7059 -3876 7065
rect -3910 6987 -3876 6997
rect -3910 6915 -3876 6929
rect -3910 6843 -3876 6861
rect -3910 6771 -3876 6793
rect -3910 6699 -3876 6725
rect -3910 6627 -3876 6657
rect -3910 6555 -3876 6589
rect -3910 6487 -3876 6521
rect -3910 6419 -3876 6449
rect -3910 6351 -3876 6377
rect -3910 6283 -3876 6305
rect -3910 6215 -3876 6233
rect -3910 6147 -3876 6161
rect -3910 6079 -3876 6089
rect -3910 6011 -3876 6017
rect -3910 5943 -3876 5945
rect -3910 5907 -3876 5909
rect -3910 5835 -3876 5841
rect -3910 5763 -3876 5773
rect -3910 5691 -3876 5705
rect -3910 5619 -3876 5637
rect -3910 5534 -3876 5569
rect -3652 7507 -3618 7542
rect -3652 7439 -3618 7457
rect -3652 7371 -3618 7385
rect -3652 7303 -3618 7313
rect -3652 7235 -3618 7241
rect -3652 7167 -3618 7169
rect -3652 7131 -3618 7133
rect -3652 7059 -3618 7065
rect -3652 6987 -3618 6997
rect -3652 6915 -3618 6929
rect -3652 6843 -3618 6861
rect -3652 6771 -3618 6793
rect -3652 6699 -3618 6725
rect -3652 6627 -3618 6657
rect -3652 6555 -3618 6589
rect -3652 6487 -3618 6521
rect -3652 6419 -3618 6449
rect -3652 6351 -3618 6377
rect -3652 6283 -3618 6305
rect -3652 6215 -3618 6233
rect -3652 6147 -3618 6161
rect -3652 6079 -3618 6089
rect -3652 6011 -3618 6017
rect -3652 5943 -3618 5945
rect -3652 5907 -3618 5909
rect -3652 5835 -3618 5841
rect -3652 5763 -3618 5773
rect -3652 5691 -3618 5705
rect -3652 5619 -3618 5637
rect -3652 5534 -3618 5569
rect -3470 7524 -3456 7558
rect -3422 7524 -3408 7558
rect -3470 7490 -3408 7524
rect -3470 7456 -3456 7490
rect -3422 7456 -3408 7490
rect -3470 7422 -3408 7456
rect -3470 7388 -3456 7422
rect -3422 7388 -3408 7422
rect -3470 7354 -3408 7388
rect -3470 7320 -3456 7354
rect -3422 7320 -3408 7354
rect -3470 7286 -3408 7320
rect -3470 7252 -3456 7286
rect -3422 7252 -3408 7286
rect -3470 7218 -3408 7252
rect -3470 7184 -3456 7218
rect -3422 7184 -3408 7218
rect -3470 7150 -3408 7184
rect -3470 7116 -3456 7150
rect -3422 7116 -3408 7150
rect -3470 7082 -3408 7116
rect -3470 7048 -3456 7082
rect -3422 7048 -3408 7082
rect -3470 7014 -3408 7048
rect -3470 6980 -3456 7014
rect -3422 6980 -3408 7014
rect -3470 6946 -3408 6980
rect -3470 6912 -3456 6946
rect -3422 6912 -3408 6946
rect -3470 6878 -3408 6912
rect -3470 6844 -3456 6878
rect -3422 6844 -3408 6878
rect -3470 6810 -3408 6844
rect -3470 6776 -3456 6810
rect -3422 6776 -3408 6810
rect -3470 6742 -3408 6776
rect -3470 6708 -3456 6742
rect -3422 6708 -3408 6742
rect -3470 6674 -3408 6708
rect -3470 6640 -3456 6674
rect -3422 6640 -3408 6674
rect -3470 6606 -3408 6640
rect -3470 6572 -3456 6606
rect -3422 6572 -3408 6606
rect -3470 6538 -3408 6572
rect -3470 6504 -3456 6538
rect -3422 6504 -3408 6538
rect -3470 6470 -3408 6504
rect -3470 6436 -3456 6470
rect -3422 6436 -3408 6470
rect -3470 6402 -3408 6436
rect -3470 6368 -3456 6402
rect -3422 6368 -3408 6402
rect -3470 6334 -3408 6368
rect -3470 6300 -3456 6334
rect -3422 6300 -3408 6334
rect -3470 6266 -3408 6300
rect -3470 6232 -3456 6266
rect -3422 6232 -3408 6266
rect -3470 6198 -3408 6232
rect -3470 6164 -3456 6198
rect -3422 6164 -3408 6198
rect -3470 6130 -3408 6164
rect -3470 6096 -3456 6130
rect -3422 6096 -3408 6130
rect -3470 6062 -3408 6096
rect -3470 6028 -3456 6062
rect -3422 6028 -3408 6062
rect -3470 5994 -3408 6028
rect -3470 5960 -3456 5994
rect -3422 5960 -3408 5994
rect -3470 5926 -3408 5960
rect -3470 5892 -3456 5926
rect -3422 5892 -3408 5926
rect -3470 5885 -3408 5892
rect -3470 5824 -3456 5885
rect -3422 5824 -3408 5885
rect -3470 5813 -3408 5824
rect -3470 5756 -3456 5813
rect -3422 5756 -3408 5813
rect -3470 5741 -3408 5756
rect -3470 5688 -3456 5741
rect -3422 5688 -3408 5741
rect -3470 5654 -3408 5688
rect -3470 5620 -3456 5654
rect -3422 5620 -3408 5654
rect -3470 5586 -3408 5620
rect -3470 5552 -3456 5586
rect -3422 5552 -3408 5586
rect -7984 5472 -7968 5506
rect -7934 5472 -7918 5506
rect -3470 5518 -3408 5552
rect -7984 5438 -7918 5472
rect -7734 5466 -7687 5500
rect -7651 5466 -7617 5500
rect -7581 5466 -7534 5500
rect -7476 5466 -7429 5500
rect -7393 5466 -7359 5500
rect -7323 5466 -7276 5500
rect -7218 5466 -7171 5500
rect -7135 5466 -7101 5500
rect -7065 5466 -7018 5500
rect -6960 5466 -6913 5500
rect -6877 5466 -6843 5500
rect -6807 5466 -6760 5500
rect -6702 5466 -6655 5500
rect -6619 5466 -6585 5500
rect -6549 5466 -6502 5500
rect -6444 5466 -6397 5500
rect -6361 5466 -6327 5500
rect -6291 5466 -6244 5500
rect -6186 5466 -6139 5500
rect -6103 5466 -6069 5500
rect -6033 5466 -5986 5500
rect -5928 5466 -5881 5500
rect -5845 5466 -5811 5500
rect -5775 5466 -5728 5500
rect -5670 5466 -5623 5500
rect -5587 5466 -5553 5500
rect -5517 5466 -5470 5500
rect -5412 5466 -5365 5500
rect -5329 5466 -5295 5500
rect -5259 5466 -5212 5500
rect -5154 5466 -5107 5500
rect -5071 5466 -5037 5500
rect -5001 5466 -4954 5500
rect -4896 5466 -4849 5500
rect -4813 5466 -4779 5500
rect -4743 5466 -4696 5500
rect -4638 5466 -4591 5500
rect -4555 5466 -4521 5500
rect -4485 5466 -4438 5500
rect -4380 5466 -4333 5500
rect -4297 5466 -4263 5500
rect -4227 5466 -4180 5500
rect -4122 5466 -4075 5500
rect -4039 5466 -4005 5500
rect -3969 5466 -3922 5500
rect -3864 5466 -3817 5500
rect -3781 5466 -3747 5500
rect -3711 5466 -3664 5500
rect -3470 5484 -3456 5518
rect -3422 5484 -3408 5518
rect -7984 5404 -7968 5438
rect -7934 5404 -7918 5438
rect -7984 5292 -7918 5404
rect -3470 5450 -3408 5484
rect -3470 5416 -3456 5450
rect -3422 5416 -3408 5450
rect -3470 5292 -3408 5416
rect -7984 5289 -3408 5292
rect 12756 8335 14060 8342
rect 12756 8286 12871 8335
rect 12756 8252 12806 8286
rect 12840 8252 12871 8286
rect 13961 8286 14060 8335
rect 12756 8196 12871 8252
rect 12756 8162 12806 8196
rect 12840 8162 12871 8196
rect 12756 8106 12871 8162
rect 12756 8072 12806 8106
rect 12840 8072 12871 8106
rect 12756 8016 12871 8072
rect 12756 7982 12806 8016
rect 12840 7982 12871 8016
rect 12756 7926 12871 7982
rect 12756 7892 12806 7926
rect 12840 7892 12871 7926
rect 12756 7836 12871 7892
rect 12756 7802 12806 7836
rect 12840 7802 12871 7836
rect 12756 7746 12871 7802
rect 12756 7712 12806 7746
rect 12840 7712 12871 7746
rect 12756 7656 12871 7712
rect 12756 7622 12806 7656
rect 12840 7622 12871 7656
rect 12756 7566 12871 7622
rect 12756 7532 12806 7566
rect 12840 7532 12871 7566
rect 12756 7476 12871 7532
rect 12756 7442 12806 7476
rect 12840 7442 12871 7476
rect 12756 7386 12871 7442
rect 12935 8252 13897 8271
rect 12935 8218 13066 8252
rect 13100 8218 13156 8252
rect 13190 8218 13246 8252
rect 13280 8218 13336 8252
rect 13370 8218 13426 8252
rect 13460 8218 13516 8252
rect 13550 8218 13606 8252
rect 13640 8218 13696 8252
rect 13730 8218 13786 8252
rect 13820 8218 13897 8252
rect 12935 8199 13897 8218
rect 12935 8195 13007 8199
rect 12935 8161 12954 8195
rect 12988 8161 13007 8195
rect 12935 8105 13007 8161
rect 13825 8176 13897 8199
rect 13825 8142 13844 8176
rect 13878 8142 13897 8176
rect 12935 8071 12954 8105
rect 12988 8071 13007 8105
rect 12935 8015 13007 8071
rect 12935 7981 12954 8015
rect 12988 7981 13007 8015
rect 12935 7925 13007 7981
rect 12935 7891 12954 7925
rect 12988 7891 13007 7925
rect 12935 7835 13007 7891
rect 12935 7801 12954 7835
rect 12988 7801 13007 7835
rect 12935 7745 13007 7801
rect 12935 7711 12954 7745
rect 12988 7711 13007 7745
rect 12935 7655 13007 7711
rect 12935 7621 12954 7655
rect 12988 7621 13007 7655
rect 12935 7565 13007 7621
rect 12935 7531 12954 7565
rect 12988 7531 13007 7565
rect 12935 7475 13007 7531
rect 12935 7441 12954 7475
rect 12988 7441 13007 7475
rect 13069 8078 13763 8137
rect 13069 8044 13130 8078
rect 13164 8050 13220 8078
rect 13254 8050 13310 8078
rect 13344 8050 13400 8078
rect 13176 8044 13220 8050
rect 13276 8044 13310 8050
rect 13376 8044 13400 8050
rect 13434 8050 13490 8078
rect 13434 8044 13442 8050
rect 13069 8016 13142 8044
rect 13176 8016 13242 8044
rect 13276 8016 13342 8044
rect 13376 8016 13442 8044
rect 13476 8044 13490 8050
rect 13524 8050 13580 8078
rect 13524 8044 13542 8050
rect 13476 8016 13542 8044
rect 13576 8044 13580 8050
rect 13614 8050 13670 8078
rect 13614 8044 13642 8050
rect 13704 8044 13763 8078
rect 13576 8016 13642 8044
rect 13676 8016 13763 8044
rect 13069 7988 13763 8016
rect 13069 7954 13130 7988
rect 13164 7954 13220 7988
rect 13254 7954 13310 7988
rect 13344 7954 13400 7988
rect 13434 7954 13490 7988
rect 13524 7954 13580 7988
rect 13614 7954 13670 7988
rect 13704 7954 13763 7988
rect 13069 7950 13763 7954
rect 13069 7916 13142 7950
rect 13176 7916 13242 7950
rect 13276 7916 13342 7950
rect 13376 7916 13442 7950
rect 13476 7916 13542 7950
rect 13576 7916 13642 7950
rect 13676 7916 13763 7950
rect 13069 7898 13763 7916
rect 13069 7864 13130 7898
rect 13164 7864 13220 7898
rect 13254 7864 13310 7898
rect 13344 7864 13400 7898
rect 13434 7864 13490 7898
rect 13524 7864 13580 7898
rect 13614 7864 13670 7898
rect 13704 7864 13763 7898
rect 13069 7850 13763 7864
rect 13069 7816 13142 7850
rect 13176 7816 13242 7850
rect 13276 7816 13342 7850
rect 13376 7816 13442 7850
rect 13476 7816 13542 7850
rect 13576 7816 13642 7850
rect 13676 7816 13763 7850
rect 13069 7808 13763 7816
rect 13069 7774 13130 7808
rect 13164 7774 13220 7808
rect 13254 7774 13310 7808
rect 13344 7774 13400 7808
rect 13434 7774 13490 7808
rect 13524 7774 13580 7808
rect 13614 7774 13670 7808
rect 13704 7774 13763 7808
rect 13069 7750 13763 7774
rect 13069 7718 13142 7750
rect 13176 7718 13242 7750
rect 13276 7718 13342 7750
rect 13376 7718 13442 7750
rect 13069 7684 13130 7718
rect 13176 7716 13220 7718
rect 13276 7716 13310 7718
rect 13376 7716 13400 7718
rect 13164 7684 13220 7716
rect 13254 7684 13310 7716
rect 13344 7684 13400 7716
rect 13434 7716 13442 7718
rect 13476 7718 13542 7750
rect 13476 7716 13490 7718
rect 13434 7684 13490 7716
rect 13524 7716 13542 7718
rect 13576 7718 13642 7750
rect 13676 7718 13763 7750
rect 13576 7716 13580 7718
rect 13524 7684 13580 7716
rect 13614 7716 13642 7718
rect 13614 7684 13670 7716
rect 13704 7684 13763 7718
rect 13069 7650 13763 7684
rect 13069 7628 13142 7650
rect 13176 7628 13242 7650
rect 13276 7628 13342 7650
rect 13376 7628 13442 7650
rect 13069 7594 13130 7628
rect 13176 7616 13220 7628
rect 13276 7616 13310 7628
rect 13376 7616 13400 7628
rect 13164 7594 13220 7616
rect 13254 7594 13310 7616
rect 13344 7594 13400 7616
rect 13434 7616 13442 7628
rect 13476 7628 13542 7650
rect 13476 7616 13490 7628
rect 13434 7594 13490 7616
rect 13524 7616 13542 7628
rect 13576 7628 13642 7650
rect 13676 7628 13763 7650
rect 13576 7616 13580 7628
rect 13524 7594 13580 7616
rect 13614 7616 13642 7628
rect 13614 7594 13670 7616
rect 13704 7594 13763 7628
rect 13069 7550 13763 7594
rect 13069 7538 13142 7550
rect 13176 7538 13242 7550
rect 13276 7538 13342 7550
rect 13376 7538 13442 7550
rect 13069 7504 13130 7538
rect 13176 7516 13220 7538
rect 13276 7516 13310 7538
rect 13376 7516 13400 7538
rect 13164 7504 13220 7516
rect 13254 7504 13310 7516
rect 13344 7504 13400 7516
rect 13434 7516 13442 7538
rect 13476 7538 13542 7550
rect 13476 7516 13490 7538
rect 13434 7504 13490 7516
rect 13524 7516 13542 7538
rect 13576 7538 13642 7550
rect 13676 7538 13763 7550
rect 13576 7516 13580 7538
rect 13524 7504 13580 7516
rect 13614 7516 13642 7538
rect 13614 7504 13670 7516
rect 13704 7504 13763 7538
rect 13069 7443 13763 7504
rect 13825 8086 13897 8142
rect 13825 8052 13844 8086
rect 13878 8052 13897 8086
rect 13825 7996 13897 8052
rect 13825 7962 13844 7996
rect 13878 7962 13897 7996
rect 13825 7906 13897 7962
rect 13825 7872 13844 7906
rect 13878 7872 13897 7906
rect 13825 7816 13897 7872
rect 13825 7782 13844 7816
rect 13878 7782 13897 7816
rect 13825 7726 13897 7782
rect 13825 7692 13844 7726
rect 13878 7692 13897 7726
rect 13825 7636 13897 7692
rect 13825 7602 13844 7636
rect 13878 7602 13897 7636
rect 13825 7546 13897 7602
rect 13825 7512 13844 7546
rect 13878 7512 13897 7546
rect 13825 7456 13897 7512
rect 12935 7390 13007 7441
rect 13825 7422 13844 7456
rect 13878 7422 13897 7456
rect 13825 7390 13897 7422
rect 12756 7352 12806 7386
rect 12840 7352 12871 7386
rect 12756 7296 12871 7352
rect 12756 7262 12806 7296
rect 12840 7262 12871 7296
rect 12756 7245 12871 7262
rect 12916 7362 13897 7390
rect 12916 7328 13032 7362
rect 13066 7328 13122 7362
rect 13156 7328 13212 7362
rect 13246 7328 13302 7362
rect 13336 7328 13392 7362
rect 13426 7328 13482 7362
rect 13516 7328 13572 7362
rect 13606 7328 13662 7362
rect 13696 7328 13752 7362
rect 13786 7328 13897 7362
rect 12916 7309 13897 7328
rect 13961 8252 13993 8286
rect 14027 8252 14060 8286
rect 13961 8196 14060 8252
rect 13961 8162 13993 8196
rect 14027 8162 14060 8196
rect 13961 8106 14060 8162
rect 13961 8072 13993 8106
rect 14027 8072 14060 8106
rect 13961 8016 14060 8072
rect 14820 8370 14854 8404
rect 14820 8302 14854 8336
rect 14820 8234 14854 8268
rect 14954 11226 14988 11251
rect 14954 11158 14988 11170
rect 14954 11090 14988 11098
rect 14954 11022 14988 11026
rect 14954 10916 14988 10920
rect 14954 10844 14988 10852
rect 14954 10772 14988 10784
rect 14954 10700 14988 10716
rect 14954 10628 14988 10648
rect 14954 10556 14988 10580
rect 14954 10484 14988 10512
rect 14954 10412 14988 10444
rect 14954 10342 14988 10376
rect 14954 10274 14988 10306
rect 14954 10206 14988 10234
rect 14954 10138 14988 10162
rect 14954 10070 14988 10090
rect 14954 10002 14988 10018
rect 14954 9934 14988 9946
rect 14954 9866 14988 9874
rect 14954 9798 14988 9802
rect 14954 9692 14988 9696
rect 14954 9620 14988 9628
rect 14954 9548 14988 9560
rect 14954 9476 14988 9492
rect 14954 9404 14988 9424
rect 14954 9332 14988 9356
rect 14954 9260 14988 9288
rect 14954 9188 14988 9220
rect 14954 9118 14988 9152
rect 14954 9050 14988 9082
rect 14954 8982 14988 9010
rect 14954 8914 14988 8938
rect 14954 8846 14988 8866
rect 14954 8778 14988 8794
rect 14954 8710 14988 8722
rect 14954 8642 14988 8650
rect 14954 8574 14988 8578
rect 14954 8468 14988 8472
rect 14954 8396 14988 8404
rect 14954 8324 14988 8336
rect 14954 8243 14988 8268
rect 16012 11226 16046 11251
rect 16012 11158 16046 11170
rect 16012 11090 16046 11098
rect 16012 11022 16046 11026
rect 16012 10916 16046 10920
rect 16012 10844 16046 10852
rect 16012 10772 16046 10784
rect 16012 10700 16046 10716
rect 16012 10628 16046 10648
rect 16012 10556 16046 10580
rect 16012 10484 16046 10512
rect 16012 10412 16046 10444
rect 16012 10342 16046 10376
rect 16012 10274 16046 10306
rect 16012 10206 16046 10234
rect 16012 10138 16046 10162
rect 16012 10070 16046 10090
rect 16012 10002 16046 10018
rect 16012 9934 16046 9946
rect 16012 9866 16046 9874
rect 16012 9798 16046 9802
rect 16012 9692 16046 9696
rect 16012 9620 16046 9628
rect 16012 9548 16046 9560
rect 16012 9476 16046 9492
rect 16012 9404 16046 9424
rect 16012 9332 16046 9356
rect 16012 9260 16046 9288
rect 16012 9188 16046 9220
rect 16012 9118 16046 9152
rect 16012 9050 16046 9082
rect 16012 8982 16046 9010
rect 16012 8914 16046 8938
rect 16012 8846 16046 8866
rect 16012 8778 16046 8794
rect 16012 8710 16046 8722
rect 16012 8642 16046 8650
rect 16012 8574 16046 8578
rect 16012 8468 16046 8472
rect 16012 8396 16046 8404
rect 16012 8324 16046 8336
rect 16012 8243 16046 8268
rect 17070 11226 17104 11251
rect 17070 11158 17104 11170
rect 17070 11090 17104 11098
rect 17070 11022 17104 11026
rect 17070 10916 17104 10920
rect 17070 10844 17104 10852
rect 17070 10772 17104 10784
rect 17070 10700 17104 10716
rect 17070 10628 17104 10648
rect 17070 10556 17104 10580
rect 17070 10484 17104 10512
rect 17070 10412 17104 10444
rect 17070 10342 17104 10376
rect 17070 10274 17104 10306
rect 17070 10206 17104 10234
rect 17070 10138 17104 10162
rect 17070 10070 17104 10090
rect 17070 10002 17104 10018
rect 17070 9934 17104 9946
rect 17070 9866 17104 9874
rect 17070 9798 17104 9802
rect 17070 9692 17104 9696
rect 17070 9620 17104 9628
rect 17070 9548 17104 9560
rect 17070 9476 17104 9492
rect 17070 9404 17104 9424
rect 17070 9332 17104 9356
rect 17070 9260 17104 9288
rect 17070 9188 17104 9220
rect 17070 9118 17104 9152
rect 17070 9050 17104 9082
rect 17070 8982 17104 9010
rect 17070 8914 17104 8938
rect 17070 8846 17104 8866
rect 17070 8778 17104 8794
rect 17070 8710 17104 8722
rect 17070 8642 17104 8650
rect 17070 8574 17104 8578
rect 17070 8468 17104 8472
rect 17070 8396 17104 8404
rect 17070 8324 17104 8336
rect 17070 8243 17104 8268
rect 17204 11226 17238 11260
rect 17204 11158 17238 11192
rect 17204 11090 17238 11124
rect 17204 11022 17238 11056
rect 17204 10954 17238 10988
rect 17204 10886 17238 10920
rect 17204 10818 17238 10852
rect 17204 10750 17238 10784
rect 17204 10682 17238 10716
rect 17204 10614 17238 10648
rect 17204 10546 17238 10580
rect 17204 10478 17238 10512
rect 17204 10410 17238 10444
rect 17204 10342 17238 10376
rect 17204 10274 17238 10308
rect 17204 10206 17238 10240
rect 17204 10138 17238 10172
rect 17204 10070 17238 10104
rect 17204 10002 17238 10036
rect 17204 9934 17238 9968
rect 17204 9866 17238 9900
rect 17204 9798 17238 9832
rect 17204 9730 17238 9764
rect 17204 9662 17238 9696
rect 17204 9594 17238 9628
rect 17204 9526 17238 9560
rect 17204 9458 17238 9492
rect 17204 9390 17238 9424
rect 17204 9322 17238 9356
rect 17204 9254 17238 9288
rect 17204 9186 17238 9220
rect 17204 9118 17238 9152
rect 17204 9050 17238 9084
rect 17204 8982 17238 9016
rect 17204 8914 17238 8948
rect 17204 8846 17238 8880
rect 17204 8778 17238 8812
rect 17204 8710 17238 8744
rect 17204 8642 17238 8676
rect 17204 8574 17238 8608
rect 17204 8506 17238 8540
rect 17204 8438 17238 8472
rect 17204 8370 17238 8404
rect 17204 8302 17238 8336
rect 17204 8234 17238 8268
rect 14820 8166 14854 8200
rect 15000 8166 15041 8200
rect 15085 8166 15109 8200
rect 15157 8166 15177 8200
rect 15229 8166 15245 8200
rect 15301 8166 15313 8200
rect 15373 8166 15381 8200
rect 15445 8166 15449 8200
rect 15551 8166 15555 8200
rect 15619 8166 15627 8200
rect 15687 8166 15699 8200
rect 15755 8166 15771 8200
rect 15823 8166 15843 8200
rect 15891 8166 15915 8200
rect 15959 8166 16000 8200
rect 16058 8166 16099 8200
rect 16143 8166 16167 8200
rect 16215 8166 16235 8200
rect 16287 8166 16303 8200
rect 16359 8166 16371 8200
rect 16431 8166 16439 8200
rect 16503 8166 16507 8200
rect 16609 8166 16613 8200
rect 16677 8166 16685 8200
rect 16745 8166 16757 8200
rect 16813 8166 16829 8200
rect 16881 8166 16901 8200
rect 16949 8166 16973 8200
rect 17017 8166 17058 8200
rect 17204 8166 17238 8200
rect 14820 8062 14854 8132
rect 17204 8062 17238 8132
rect 14820 8028 14924 8062
rect 14958 8028 14992 8062
rect 15026 8028 15060 8062
rect 15094 8028 15128 8062
rect 15162 8028 15196 8062
rect 15230 8028 15264 8062
rect 15298 8028 15332 8062
rect 15366 8028 15400 8062
rect 15434 8028 15468 8062
rect 15502 8028 15536 8062
rect 15570 8028 15604 8062
rect 15638 8028 15672 8062
rect 15706 8028 15740 8062
rect 15774 8028 15808 8062
rect 15842 8028 15876 8062
rect 15910 8028 15944 8062
rect 15978 8028 16012 8062
rect 16046 8028 16080 8062
rect 16114 8028 16148 8062
rect 16182 8028 16216 8062
rect 16250 8028 16284 8062
rect 16318 8028 16352 8062
rect 16386 8028 16420 8062
rect 16454 8028 16488 8062
rect 16522 8028 16556 8062
rect 16590 8028 16624 8062
rect 16658 8028 16692 8062
rect 16726 8028 16760 8062
rect 16794 8028 16828 8062
rect 16862 8028 16896 8062
rect 16930 8028 16964 8062
rect 16998 8028 17032 8062
rect 17066 8028 17100 8062
rect 17134 8028 17238 8062
rect 17344 11406 17448 11440
rect 17482 11406 17516 11440
rect 17550 11406 17584 11440
rect 17618 11406 17652 11440
rect 17686 11406 17720 11440
rect 17754 11406 17788 11440
rect 17822 11406 17856 11440
rect 17890 11406 17924 11440
rect 17958 11406 17992 11440
rect 18026 11406 18060 11440
rect 18094 11406 18128 11440
rect 18162 11406 18196 11440
rect 18230 11406 18264 11440
rect 18298 11406 18332 11440
rect 18366 11406 18400 11440
rect 18434 11406 18468 11440
rect 18502 11406 18536 11440
rect 18570 11406 18604 11440
rect 18638 11406 18672 11440
rect 18706 11406 18740 11440
rect 18774 11406 18808 11440
rect 18842 11406 18876 11440
rect 18910 11406 18944 11440
rect 18978 11406 19012 11440
rect 19046 11406 19080 11440
rect 19114 11406 19148 11440
rect 19182 11406 19216 11440
rect 19250 11406 19284 11440
rect 19318 11406 19352 11440
rect 19386 11406 19420 11440
rect 19454 11406 19488 11440
rect 19522 11406 19556 11440
rect 19590 11406 19624 11440
rect 19658 11406 19762 11440
rect 17344 11336 17378 11406
rect 19728 11336 19762 11406
rect 17344 11268 17378 11302
rect 17524 11268 17565 11302
rect 17609 11268 17633 11302
rect 17681 11268 17701 11302
rect 17753 11268 17769 11302
rect 17825 11268 17837 11302
rect 17897 11268 17905 11302
rect 17969 11268 17973 11302
rect 18075 11268 18079 11302
rect 18143 11268 18151 11302
rect 18211 11268 18223 11302
rect 18279 11268 18295 11302
rect 18347 11268 18367 11302
rect 18415 11268 18439 11302
rect 18483 11268 18524 11302
rect 18582 11268 18623 11302
rect 18667 11268 18691 11302
rect 18739 11268 18759 11302
rect 18811 11268 18827 11302
rect 18883 11268 18895 11302
rect 18955 11268 18963 11302
rect 19027 11268 19031 11302
rect 19133 11268 19137 11302
rect 19201 11268 19209 11302
rect 19269 11268 19281 11302
rect 19337 11268 19353 11302
rect 19405 11268 19425 11302
rect 19473 11268 19497 11302
rect 19541 11268 19582 11302
rect 19728 11268 19762 11302
rect 17344 11200 17378 11234
rect 17344 11132 17378 11166
rect 17344 11064 17378 11098
rect 17344 10996 17378 11030
rect 17344 10928 17378 10962
rect 17344 10860 17378 10894
rect 17344 10792 17378 10826
rect 17344 10724 17378 10758
rect 17344 10656 17378 10690
rect 17344 10588 17378 10622
rect 17344 10520 17378 10554
rect 17344 10452 17378 10486
rect 17344 10384 17378 10418
rect 17344 10316 17378 10350
rect 17344 10248 17378 10282
rect 17344 10180 17378 10214
rect 17344 10112 17378 10146
rect 17344 10044 17378 10078
rect 17344 9976 17378 10010
rect 17344 9908 17378 9942
rect 17344 9840 17378 9874
rect 17344 9772 17378 9806
rect 17344 9704 17378 9738
rect 17344 9636 17378 9670
rect 17344 9568 17378 9602
rect 17344 9500 17378 9534
rect 17344 9432 17378 9466
rect 17344 9364 17378 9398
rect 17344 9296 17378 9330
rect 17344 9228 17378 9262
rect 17344 9160 17378 9194
rect 17344 9092 17378 9126
rect 17344 9024 17378 9058
rect 17344 8956 17378 8990
rect 17344 8888 17378 8922
rect 17344 8820 17378 8854
rect 17344 8752 17378 8786
rect 17344 8684 17378 8718
rect 17344 8616 17378 8650
rect 17344 8548 17378 8582
rect 17344 8480 17378 8514
rect 17344 8412 17378 8446
rect 17344 8344 17378 8378
rect 17344 8276 17378 8310
rect 17344 8208 17378 8242
rect 17478 11200 17512 11225
rect 17478 11132 17512 11144
rect 17478 11064 17512 11072
rect 17478 10996 17512 11000
rect 17478 10890 17512 10894
rect 17478 10818 17512 10826
rect 17478 10746 17512 10758
rect 17478 10674 17512 10690
rect 17478 10602 17512 10622
rect 17478 10530 17512 10554
rect 17478 10458 17512 10486
rect 17478 10386 17512 10418
rect 17478 10316 17512 10350
rect 17478 10248 17512 10280
rect 17478 10180 17512 10208
rect 17478 10112 17512 10136
rect 17478 10044 17512 10064
rect 17478 9976 17512 9992
rect 17478 9908 17512 9920
rect 17478 9840 17512 9848
rect 17478 9772 17512 9776
rect 17478 9666 17512 9670
rect 17478 9594 17512 9602
rect 17478 9522 17512 9534
rect 17478 9450 17512 9466
rect 17478 9378 17512 9398
rect 17478 9306 17512 9330
rect 17478 9234 17512 9262
rect 17478 9162 17512 9194
rect 17478 9092 17512 9126
rect 17478 9024 17512 9056
rect 17478 8956 17512 8984
rect 17478 8888 17512 8912
rect 17478 8820 17512 8840
rect 17478 8752 17512 8768
rect 17478 8684 17512 8696
rect 17478 8616 17512 8624
rect 17478 8548 17512 8552
rect 17478 8442 17512 8446
rect 17478 8370 17512 8378
rect 17478 8298 17512 8310
rect 17478 8217 17512 8242
rect 18536 11200 18570 11225
rect 18536 11132 18570 11144
rect 18536 11064 18570 11072
rect 18536 10996 18570 11000
rect 18536 10890 18570 10894
rect 18536 10818 18570 10826
rect 18536 10746 18570 10758
rect 18536 10674 18570 10690
rect 18536 10602 18570 10622
rect 18536 10530 18570 10554
rect 18536 10458 18570 10486
rect 18536 10386 18570 10418
rect 18536 10316 18570 10350
rect 18536 10248 18570 10280
rect 18536 10180 18570 10208
rect 18536 10112 18570 10136
rect 18536 10044 18570 10064
rect 18536 9976 18570 9992
rect 18536 9908 18570 9920
rect 18536 9840 18570 9848
rect 18536 9772 18570 9776
rect 18536 9666 18570 9670
rect 18536 9594 18570 9602
rect 18536 9522 18570 9534
rect 18536 9450 18570 9466
rect 18536 9378 18570 9398
rect 18536 9306 18570 9330
rect 18536 9234 18570 9262
rect 18536 9162 18570 9194
rect 18536 9092 18570 9126
rect 18536 9024 18570 9056
rect 18536 8956 18570 8984
rect 18536 8888 18570 8912
rect 18536 8820 18570 8840
rect 18536 8752 18570 8768
rect 18536 8684 18570 8696
rect 18536 8616 18570 8624
rect 18536 8548 18570 8552
rect 18536 8442 18570 8446
rect 18536 8370 18570 8378
rect 18536 8298 18570 8310
rect 18536 8217 18570 8242
rect 19594 11200 19628 11225
rect 19594 11132 19628 11144
rect 19594 11064 19628 11072
rect 19594 10996 19628 11000
rect 19594 10890 19628 10894
rect 19594 10818 19628 10826
rect 19594 10746 19628 10758
rect 19594 10674 19628 10690
rect 19594 10602 19628 10622
rect 19594 10530 19628 10554
rect 19594 10458 19628 10486
rect 19594 10386 19628 10418
rect 19594 10316 19628 10350
rect 19594 10248 19628 10280
rect 19594 10180 19628 10208
rect 19594 10112 19628 10136
rect 19594 10044 19628 10064
rect 19594 9976 19628 9992
rect 19594 9908 19628 9920
rect 19594 9840 19628 9848
rect 19594 9772 19628 9776
rect 19594 9666 19628 9670
rect 19594 9594 19628 9602
rect 19594 9522 19628 9534
rect 19594 9450 19628 9466
rect 19594 9378 19628 9398
rect 19594 9306 19628 9330
rect 19594 9234 19628 9262
rect 19594 9162 19628 9194
rect 19594 9092 19628 9126
rect 19594 9024 19628 9056
rect 19594 8956 19628 8984
rect 19594 8888 19628 8912
rect 19594 8820 19628 8840
rect 19594 8752 19628 8768
rect 19594 8684 19628 8696
rect 19594 8616 19628 8624
rect 19594 8548 19628 8552
rect 19594 8442 19628 8446
rect 19594 8370 19628 8378
rect 19594 8298 19628 8310
rect 19594 8217 19628 8242
rect 19728 11200 19762 11234
rect 19728 11132 19762 11166
rect 19728 11064 19762 11098
rect 19728 10996 19762 11030
rect 19728 10928 19762 10962
rect 19728 10860 19762 10894
rect 19728 10792 19762 10826
rect 19728 10724 19762 10758
rect 19728 10656 19762 10690
rect 19728 10588 19762 10622
rect 19728 10520 19762 10554
rect 19728 10452 19762 10486
rect 19728 10384 19762 10418
rect 19728 10316 19762 10350
rect 19728 10248 19762 10282
rect 19728 10180 19762 10214
rect 19728 10112 19762 10146
rect 19728 10044 19762 10078
rect 19728 9976 19762 10010
rect 19728 9908 19762 9942
rect 19728 9840 19762 9874
rect 19728 9772 19762 9806
rect 19728 9704 19762 9738
rect 19728 9636 19762 9670
rect 19728 9568 19762 9602
rect 19728 9500 19762 9534
rect 19728 9432 19762 9466
rect 19728 9364 19762 9398
rect 19728 9296 19762 9330
rect 19728 9228 19762 9262
rect 19728 9160 19762 9194
rect 19728 9092 19762 9126
rect 19728 9024 19762 9058
rect 19728 8956 19762 8990
rect 19728 8888 19762 8922
rect 19728 8820 19762 8854
rect 19728 8752 19762 8786
rect 19728 8684 19762 8718
rect 19728 8616 19762 8650
rect 19728 8548 19762 8582
rect 19728 8480 19762 8514
rect 19728 8412 19762 8446
rect 19728 8344 19762 8378
rect 19728 8276 19762 8310
rect 19728 8208 19762 8242
rect 17344 8140 17378 8174
rect 17524 8140 17565 8174
rect 17609 8140 17633 8174
rect 17681 8140 17701 8174
rect 17753 8140 17769 8174
rect 17825 8140 17837 8174
rect 17897 8140 17905 8174
rect 17969 8140 17973 8174
rect 18075 8140 18079 8174
rect 18143 8140 18151 8174
rect 18211 8140 18223 8174
rect 18279 8140 18295 8174
rect 18347 8140 18367 8174
rect 18415 8140 18439 8174
rect 18483 8140 18524 8174
rect 18582 8140 18623 8174
rect 18667 8140 18691 8174
rect 18739 8140 18759 8174
rect 18811 8140 18827 8174
rect 18883 8140 18895 8174
rect 18955 8140 18963 8174
rect 19027 8140 19031 8174
rect 19133 8140 19137 8174
rect 19201 8140 19209 8174
rect 19269 8140 19281 8174
rect 19337 8140 19353 8174
rect 19405 8140 19425 8174
rect 19473 8140 19497 8174
rect 19541 8140 19582 8174
rect 19728 8140 19762 8174
rect 17344 8036 17378 8106
rect 19728 8036 19762 8106
rect 13961 7982 13993 8016
rect 14027 7982 14060 8016
rect 17344 8002 17448 8036
rect 17482 8002 17516 8036
rect 17550 8002 17584 8036
rect 17618 8002 17652 8036
rect 17686 8002 17720 8036
rect 17754 8002 17788 8036
rect 17822 8002 17856 8036
rect 17890 8002 17924 8036
rect 17958 8002 17992 8036
rect 18026 8002 18060 8036
rect 18094 8002 18128 8036
rect 18162 8002 18196 8036
rect 18230 8002 18264 8036
rect 18298 8002 18332 8036
rect 18366 8002 18400 8036
rect 18434 8002 18468 8036
rect 18502 8002 18536 8036
rect 18570 8002 18604 8036
rect 18638 8002 18672 8036
rect 18706 8002 18740 8036
rect 18774 8002 18808 8036
rect 18842 8002 18876 8036
rect 18910 8002 18944 8036
rect 18978 8002 19012 8036
rect 19046 8002 19080 8036
rect 19114 8002 19148 8036
rect 19182 8002 19216 8036
rect 19250 8002 19284 8036
rect 19318 8002 19352 8036
rect 19386 8002 19420 8036
rect 19454 8002 19488 8036
rect 19522 8002 19556 8036
rect 19590 8002 19624 8036
rect 19658 8002 19762 8036
rect 20382 11414 20416 11448
rect 20382 11346 20416 11380
rect 20382 11278 20416 11312
rect 20382 11210 20416 11244
rect 20382 11142 20416 11176
rect 20382 11074 20416 11108
rect 20382 11006 20416 11040
rect 20382 10938 20416 10972
rect 20382 10870 20416 10904
rect 20382 10802 20416 10836
rect 20382 10734 20416 10768
rect 20382 10666 20416 10700
rect 20382 10598 20416 10632
rect 20382 10530 20416 10564
rect 20382 10462 20416 10496
rect 20382 10394 20416 10428
rect 20382 10326 20416 10360
rect 20382 10258 20416 10292
rect 20382 10190 20416 10224
rect 20382 10122 20416 10156
rect 20382 10054 20416 10088
rect 20382 9986 20416 10020
rect 20382 9918 20416 9952
rect 20382 9850 20416 9884
rect 20382 9782 20416 9816
rect 20382 9714 20416 9748
rect 20382 9646 20416 9680
rect 20382 9578 20416 9612
rect 20382 9510 20416 9544
rect 20382 9442 20416 9476
rect 20382 9374 20416 9408
rect 20382 9306 20416 9340
rect 20382 9238 20416 9272
rect 20382 9170 20416 9204
rect 20382 9102 20416 9136
rect 20382 9034 20416 9068
rect 20382 8966 20416 9000
rect 20382 8898 20416 8932
rect 20382 8830 20416 8864
rect 20382 8762 20416 8796
rect 20382 8694 20416 8728
rect 20382 8626 20416 8660
rect 20382 8558 20416 8592
rect 20382 8490 20416 8524
rect 20382 8422 20416 8456
rect 20382 8354 20416 8388
rect 20382 8286 20416 8320
rect 20382 8218 20416 8252
rect 20382 8150 20416 8184
rect 20382 8082 20416 8116
rect 20382 8014 20416 8048
rect 13961 7926 14060 7982
rect 13961 7892 13993 7926
rect 14027 7892 14060 7926
rect 13961 7836 14060 7892
rect 13961 7802 13993 7836
rect 14027 7802 14060 7836
rect 13961 7746 14060 7802
rect 20382 7946 20416 7980
rect 20382 7878 20416 7912
rect 20382 7810 20416 7844
rect 13961 7712 13993 7746
rect 14027 7712 14060 7746
rect 13961 7656 14060 7712
rect 13961 7622 13993 7656
rect 14027 7622 14060 7656
rect 13961 7566 14060 7622
rect 13961 7532 13993 7566
rect 14027 7532 14060 7566
rect 13961 7476 14060 7532
rect 13961 7442 13993 7476
rect 14027 7442 14060 7476
rect 13961 7386 14060 7442
rect 13961 7352 13993 7386
rect 14027 7352 14060 7386
rect 12916 7245 13876 7309
rect 13961 7296 14060 7352
rect 13961 7262 13993 7296
rect 14027 7262 14060 7296
rect 13961 7245 14060 7262
rect 12756 7212 14060 7245
rect 17300 7724 17419 7758
rect 17453 7724 17487 7758
rect 17521 7724 17555 7758
rect 17589 7724 17623 7758
rect 17657 7724 17691 7758
rect 17725 7724 17759 7758
rect 17793 7724 17827 7758
rect 17861 7724 17895 7758
rect 17929 7724 17963 7758
rect 17997 7724 18031 7758
rect 18065 7724 18099 7758
rect 18133 7724 18167 7758
rect 18201 7724 18235 7758
rect 18269 7724 18303 7758
rect 18337 7724 18371 7758
rect 18405 7724 18439 7758
rect 18473 7724 18507 7758
rect 18541 7724 18660 7758
rect 17300 7629 17334 7724
rect 18626 7629 18660 7724
rect 17300 7561 17334 7595
rect 17480 7586 17521 7620
rect 17565 7586 17589 7620
rect 17637 7586 17657 7620
rect 17709 7586 17725 7620
rect 17781 7586 17793 7620
rect 17853 7586 17861 7620
rect 17925 7586 17929 7620
rect 18031 7586 18035 7620
rect 18099 7586 18107 7620
rect 18167 7586 18179 7620
rect 18235 7586 18251 7620
rect 18303 7586 18323 7620
rect 18371 7586 18395 7620
rect 18439 7586 18480 7620
rect 18626 7561 18660 7595
rect 17300 7493 17334 7527
rect 17300 7425 17334 7459
rect 17300 7357 17334 7391
rect 17300 7289 17334 7323
rect 12756 7178 12902 7212
rect 12936 7178 12992 7212
rect 13026 7178 13082 7212
rect 13116 7178 13172 7212
rect 13206 7178 13262 7212
rect 13296 7178 13352 7212
rect 13386 7178 13442 7212
rect 13476 7178 13532 7212
rect 13566 7178 13622 7212
rect 13656 7178 13712 7212
rect 13746 7178 13802 7212
rect 13836 7178 13892 7212
rect 13926 7178 14060 7212
rect 12756 7146 14060 7178
rect 16080 7206 16206 7240
rect 16240 7206 16274 7240
rect 16308 7206 16342 7240
rect 16376 7206 16410 7240
rect 16444 7206 16478 7240
rect 16512 7206 16546 7240
rect 16580 7206 16614 7240
rect 16648 7206 16682 7240
rect 16716 7206 16750 7240
rect 16784 7206 16818 7240
rect 16852 7206 16886 7240
rect 16920 7206 17046 7240
rect 12756 7084 12856 7146
rect 12916 7140 13876 7146
rect 16080 7119 16114 7206
rect 14422 7110 15710 7114
rect 12756 7049 14060 7084
rect 12756 7026 12902 7049
rect 12756 6992 12806 7026
rect 12840 7015 12902 7026
rect 12936 7015 12992 7049
rect 13026 7015 13082 7049
rect 13116 7015 13172 7049
rect 13206 7015 13262 7049
rect 13296 7015 13352 7049
rect 13386 7015 13442 7049
rect 13476 7015 13532 7049
rect 13566 7015 13622 7049
rect 13656 7015 13712 7049
rect 13746 7015 13802 7049
rect 13836 7015 13892 7049
rect 13926 7026 14060 7049
rect 13926 7015 13993 7026
rect 12840 6992 13993 7015
rect 14027 6992 14060 7026
rect 12756 6985 14060 6992
rect 12756 6936 12871 6985
rect 12756 6902 12806 6936
rect 12840 6902 12871 6936
rect 13961 6936 14060 6985
rect 12756 6846 12871 6902
rect 12756 6812 12806 6846
rect 12840 6812 12871 6846
rect 12756 6756 12871 6812
rect 12756 6722 12806 6756
rect 12840 6722 12871 6756
rect 12756 6666 12871 6722
rect 12756 6632 12806 6666
rect 12840 6632 12871 6666
rect 12756 6576 12871 6632
rect 12756 6542 12806 6576
rect 12840 6542 12871 6576
rect 12756 6486 12871 6542
rect 12756 6452 12806 6486
rect 12840 6452 12871 6486
rect 12756 6396 12871 6452
rect 12756 6362 12806 6396
rect 12840 6362 12871 6396
rect 12756 6306 12871 6362
rect 12756 6272 12806 6306
rect 12840 6272 12871 6306
rect 12756 6216 12871 6272
rect 12756 6182 12806 6216
rect 12840 6182 12871 6216
rect 12756 6126 12871 6182
rect 12756 6092 12806 6126
rect 12840 6092 12871 6126
rect 12756 6036 12871 6092
rect 12756 6002 12806 6036
rect 12840 6002 12871 6036
rect 12935 6902 13897 6921
rect 12935 6868 13066 6902
rect 13100 6868 13156 6902
rect 13190 6868 13246 6902
rect 13280 6868 13336 6902
rect 13370 6868 13426 6902
rect 13460 6868 13516 6902
rect 13550 6868 13606 6902
rect 13640 6868 13696 6902
rect 13730 6868 13786 6902
rect 13820 6868 13897 6902
rect 12935 6849 13897 6868
rect 12935 6845 13007 6849
rect 12935 6811 12954 6845
rect 12988 6811 13007 6845
rect 12935 6755 13007 6811
rect 13825 6826 13897 6849
rect 13825 6792 13844 6826
rect 13878 6792 13897 6826
rect 12935 6721 12954 6755
rect 12988 6721 13007 6755
rect 12935 6665 13007 6721
rect 12935 6631 12954 6665
rect 12988 6631 13007 6665
rect 12935 6575 13007 6631
rect 12935 6541 12954 6575
rect 12988 6541 13007 6575
rect 12935 6485 13007 6541
rect 12935 6451 12954 6485
rect 12988 6451 13007 6485
rect 12935 6395 13007 6451
rect 12935 6361 12954 6395
rect 12988 6361 13007 6395
rect 12935 6305 13007 6361
rect 12935 6271 12954 6305
rect 12988 6271 13007 6305
rect 12935 6215 13007 6271
rect 12935 6181 12954 6215
rect 12988 6181 13007 6215
rect 12935 6125 13007 6181
rect 12935 6091 12954 6125
rect 12988 6091 13007 6125
rect 13069 6728 13763 6787
rect 13069 6694 13130 6728
rect 13164 6700 13220 6728
rect 13254 6700 13310 6728
rect 13344 6700 13400 6728
rect 13176 6694 13220 6700
rect 13276 6694 13310 6700
rect 13376 6694 13400 6700
rect 13434 6700 13490 6728
rect 13434 6694 13442 6700
rect 13069 6666 13142 6694
rect 13176 6666 13242 6694
rect 13276 6666 13342 6694
rect 13376 6666 13442 6694
rect 13476 6694 13490 6700
rect 13524 6700 13580 6728
rect 13524 6694 13542 6700
rect 13476 6666 13542 6694
rect 13576 6694 13580 6700
rect 13614 6700 13670 6728
rect 13614 6694 13642 6700
rect 13704 6694 13763 6728
rect 13576 6666 13642 6694
rect 13676 6666 13763 6694
rect 13069 6638 13763 6666
rect 13069 6604 13130 6638
rect 13164 6604 13220 6638
rect 13254 6604 13310 6638
rect 13344 6604 13400 6638
rect 13434 6604 13490 6638
rect 13524 6604 13580 6638
rect 13614 6604 13670 6638
rect 13704 6604 13763 6638
rect 13069 6600 13763 6604
rect 13069 6566 13142 6600
rect 13176 6566 13242 6600
rect 13276 6566 13342 6600
rect 13376 6566 13442 6600
rect 13476 6566 13542 6600
rect 13576 6566 13642 6600
rect 13676 6566 13763 6600
rect 13069 6548 13763 6566
rect 13069 6514 13130 6548
rect 13164 6514 13220 6548
rect 13254 6514 13310 6548
rect 13344 6514 13400 6548
rect 13434 6514 13490 6548
rect 13524 6514 13580 6548
rect 13614 6514 13670 6548
rect 13704 6514 13763 6548
rect 13069 6500 13763 6514
rect 13069 6466 13142 6500
rect 13176 6466 13242 6500
rect 13276 6466 13342 6500
rect 13376 6466 13442 6500
rect 13476 6466 13542 6500
rect 13576 6466 13642 6500
rect 13676 6466 13763 6500
rect 13069 6458 13763 6466
rect 13069 6424 13130 6458
rect 13164 6424 13220 6458
rect 13254 6424 13310 6458
rect 13344 6424 13400 6458
rect 13434 6424 13490 6458
rect 13524 6424 13580 6458
rect 13614 6424 13670 6458
rect 13704 6424 13763 6458
rect 13069 6400 13763 6424
rect 13069 6368 13142 6400
rect 13176 6368 13242 6400
rect 13276 6368 13342 6400
rect 13376 6368 13442 6400
rect 13069 6334 13130 6368
rect 13176 6366 13220 6368
rect 13276 6366 13310 6368
rect 13376 6366 13400 6368
rect 13164 6334 13220 6366
rect 13254 6334 13310 6366
rect 13344 6334 13400 6366
rect 13434 6366 13442 6368
rect 13476 6368 13542 6400
rect 13476 6366 13490 6368
rect 13434 6334 13490 6366
rect 13524 6366 13542 6368
rect 13576 6368 13642 6400
rect 13676 6368 13763 6400
rect 13576 6366 13580 6368
rect 13524 6334 13580 6366
rect 13614 6366 13642 6368
rect 13614 6334 13670 6366
rect 13704 6334 13763 6368
rect 13069 6300 13763 6334
rect 13069 6278 13142 6300
rect 13176 6278 13242 6300
rect 13276 6278 13342 6300
rect 13376 6278 13442 6300
rect 13069 6244 13130 6278
rect 13176 6266 13220 6278
rect 13276 6266 13310 6278
rect 13376 6266 13400 6278
rect 13164 6244 13220 6266
rect 13254 6244 13310 6266
rect 13344 6244 13400 6266
rect 13434 6266 13442 6278
rect 13476 6278 13542 6300
rect 13476 6266 13490 6278
rect 13434 6244 13490 6266
rect 13524 6266 13542 6278
rect 13576 6278 13642 6300
rect 13676 6278 13763 6300
rect 13576 6266 13580 6278
rect 13524 6244 13580 6266
rect 13614 6266 13642 6278
rect 13614 6244 13670 6266
rect 13704 6244 13763 6278
rect 13069 6200 13763 6244
rect 13069 6188 13142 6200
rect 13176 6188 13242 6200
rect 13276 6188 13342 6200
rect 13376 6188 13442 6200
rect 13069 6154 13130 6188
rect 13176 6166 13220 6188
rect 13276 6166 13310 6188
rect 13376 6166 13400 6188
rect 13164 6154 13220 6166
rect 13254 6154 13310 6166
rect 13344 6154 13400 6166
rect 13434 6166 13442 6188
rect 13476 6188 13542 6200
rect 13476 6166 13490 6188
rect 13434 6154 13490 6166
rect 13524 6166 13542 6188
rect 13576 6188 13642 6200
rect 13676 6188 13763 6200
rect 13576 6166 13580 6188
rect 13524 6154 13580 6166
rect 13614 6166 13642 6188
rect 13614 6154 13670 6166
rect 13704 6154 13763 6188
rect 13069 6093 13763 6154
rect 13825 6736 13897 6792
rect 13825 6702 13844 6736
rect 13878 6702 13897 6736
rect 13825 6646 13897 6702
rect 13825 6612 13844 6646
rect 13878 6612 13897 6646
rect 13825 6556 13897 6612
rect 13825 6522 13844 6556
rect 13878 6522 13897 6556
rect 13825 6466 13897 6522
rect 13825 6432 13844 6466
rect 13878 6432 13897 6466
rect 13825 6376 13897 6432
rect 13825 6342 13844 6376
rect 13878 6342 13897 6376
rect 13825 6286 13897 6342
rect 13825 6252 13844 6286
rect 13878 6252 13897 6286
rect 13825 6196 13897 6252
rect 13825 6162 13844 6196
rect 13878 6162 13897 6196
rect 13825 6106 13897 6162
rect 12935 6031 13007 6091
rect 13825 6072 13844 6106
rect 13878 6072 13897 6106
rect 13825 6031 13897 6072
rect 12935 6030 13897 6031
rect 12756 5946 12871 6002
rect 12756 5912 12806 5946
rect 12840 5912 12871 5946
rect 12756 5895 12871 5912
rect 12916 6012 13897 6030
rect 12916 5978 13032 6012
rect 13066 5978 13122 6012
rect 13156 5978 13212 6012
rect 13246 5978 13302 6012
rect 13336 5978 13392 6012
rect 13426 5978 13482 6012
rect 13516 5978 13572 6012
rect 13606 5978 13662 6012
rect 13696 5978 13752 6012
rect 13786 5978 13897 6012
rect 12916 5959 13897 5978
rect 13961 6902 13993 6936
rect 14027 6902 14060 6936
rect 13961 6846 14060 6902
rect 13961 6812 13993 6846
rect 14027 6812 14060 6846
rect 13961 6756 14060 6812
rect 13961 6722 13993 6756
rect 14027 6722 14060 6756
rect 13961 6666 14060 6722
rect 13961 6632 13993 6666
rect 14027 6632 14060 6666
rect 13961 6576 14060 6632
rect 13961 6542 13993 6576
rect 14027 6542 14060 6576
rect 13961 6486 14060 6542
rect 13961 6452 13993 6486
rect 14027 6452 14060 6486
rect 13961 6396 14060 6452
rect 13961 6362 13993 6396
rect 14027 6362 14060 6396
rect 13961 6306 14060 6362
rect 13961 6272 13993 6306
rect 14027 6272 14060 6306
rect 13961 6216 14060 6272
rect 13961 6182 13993 6216
rect 14027 6182 14060 6216
rect 13961 6126 14060 6182
rect 13961 6092 13993 6126
rect 14027 6092 14060 6126
rect 13961 6036 14060 6092
rect 13961 6002 13993 6036
rect 14027 6002 14060 6036
rect 12916 5895 13876 5959
rect 13961 5946 14060 6002
rect 13961 5912 13993 5946
rect 14027 5912 14060 5946
rect 13961 5895 14060 5912
rect 12756 5862 14060 5895
rect 12756 5828 12902 5862
rect 12936 5828 12992 5862
rect 13026 5828 13082 5862
rect 13116 5828 13172 5862
rect 13206 5828 13262 5862
rect 13296 5828 13352 5862
rect 13386 5828 13442 5862
rect 13476 5828 13532 5862
rect 13566 5828 13622 5862
rect 13656 5828 13712 5862
rect 13746 5828 13802 5862
rect 13836 5828 13892 5862
rect 13926 5828 14060 5862
rect 12756 5796 14060 5828
rect 14406 7079 15710 7110
rect 14406 7056 14552 7079
rect 14406 7022 14456 7056
rect 14490 7045 14552 7056
rect 14586 7045 14642 7079
rect 14676 7045 14732 7079
rect 14766 7045 14822 7079
rect 14856 7045 14912 7079
rect 14946 7045 15002 7079
rect 15036 7045 15092 7079
rect 15126 7045 15182 7079
rect 15216 7045 15272 7079
rect 15306 7045 15362 7079
rect 15396 7045 15452 7079
rect 15486 7045 15542 7079
rect 15576 7056 15710 7079
rect 15576 7045 15643 7056
rect 14490 7022 15643 7045
rect 15677 7022 15710 7056
rect 14406 7015 15710 7022
rect 14406 6966 14521 7015
rect 14406 6932 14456 6966
rect 14490 6932 14521 6966
rect 15611 6966 15710 7015
rect 14406 6876 14521 6932
rect 14406 6842 14456 6876
rect 14490 6842 14521 6876
rect 14406 6786 14521 6842
rect 14406 6752 14456 6786
rect 14490 6752 14521 6786
rect 14406 6696 14521 6752
rect 14406 6662 14456 6696
rect 14490 6662 14521 6696
rect 14406 6606 14521 6662
rect 14406 6572 14456 6606
rect 14490 6572 14521 6606
rect 14406 6516 14521 6572
rect 14406 6482 14456 6516
rect 14490 6482 14521 6516
rect 14406 6426 14521 6482
rect 14406 6392 14456 6426
rect 14490 6392 14521 6426
rect 14406 6336 14521 6392
rect 14406 6302 14456 6336
rect 14490 6302 14521 6336
rect 14406 6246 14521 6302
rect 14406 6212 14456 6246
rect 14490 6212 14521 6246
rect 14406 6156 14521 6212
rect 14406 6122 14456 6156
rect 14490 6122 14521 6156
rect 14406 6066 14521 6122
rect 14406 6032 14456 6066
rect 14490 6032 14521 6066
rect 14585 6932 15547 6951
rect 14585 6898 14716 6932
rect 14750 6898 14806 6932
rect 14840 6898 14896 6932
rect 14930 6898 14986 6932
rect 15020 6898 15076 6932
rect 15110 6898 15166 6932
rect 15200 6898 15256 6932
rect 15290 6898 15346 6932
rect 15380 6898 15436 6932
rect 15470 6898 15547 6932
rect 14585 6879 15547 6898
rect 14585 6875 14657 6879
rect 14585 6841 14604 6875
rect 14638 6841 14657 6875
rect 14585 6785 14657 6841
rect 15475 6856 15547 6879
rect 15475 6822 15494 6856
rect 15528 6822 15547 6856
rect 14585 6751 14604 6785
rect 14638 6751 14657 6785
rect 14585 6695 14657 6751
rect 14585 6661 14604 6695
rect 14638 6661 14657 6695
rect 14585 6605 14657 6661
rect 14585 6571 14604 6605
rect 14638 6571 14657 6605
rect 14585 6515 14657 6571
rect 14585 6481 14604 6515
rect 14638 6481 14657 6515
rect 14585 6425 14657 6481
rect 14585 6391 14604 6425
rect 14638 6391 14657 6425
rect 14585 6335 14657 6391
rect 14585 6301 14604 6335
rect 14638 6301 14657 6335
rect 14585 6245 14657 6301
rect 14585 6211 14604 6245
rect 14638 6211 14657 6245
rect 14585 6155 14657 6211
rect 14585 6121 14604 6155
rect 14638 6121 14657 6155
rect 14719 6758 15413 6817
rect 14719 6724 14780 6758
rect 14814 6730 14870 6758
rect 14904 6730 14960 6758
rect 14994 6730 15050 6758
rect 14826 6724 14870 6730
rect 14926 6724 14960 6730
rect 15026 6724 15050 6730
rect 15084 6730 15140 6758
rect 15084 6724 15092 6730
rect 14719 6696 14792 6724
rect 14826 6696 14892 6724
rect 14926 6696 14992 6724
rect 15026 6696 15092 6724
rect 15126 6724 15140 6730
rect 15174 6730 15230 6758
rect 15174 6724 15192 6730
rect 15126 6696 15192 6724
rect 15226 6724 15230 6730
rect 15264 6730 15320 6758
rect 15264 6724 15292 6730
rect 15354 6724 15413 6758
rect 15226 6696 15292 6724
rect 15326 6696 15413 6724
rect 14719 6668 15413 6696
rect 14719 6634 14780 6668
rect 14814 6634 14870 6668
rect 14904 6634 14960 6668
rect 14994 6634 15050 6668
rect 15084 6634 15140 6668
rect 15174 6634 15230 6668
rect 15264 6634 15320 6668
rect 15354 6634 15413 6668
rect 14719 6630 15413 6634
rect 14719 6596 14792 6630
rect 14826 6596 14892 6630
rect 14926 6596 14992 6630
rect 15026 6596 15092 6630
rect 15126 6596 15192 6630
rect 15226 6596 15292 6630
rect 15326 6596 15413 6630
rect 14719 6578 15413 6596
rect 14719 6544 14780 6578
rect 14814 6544 14870 6578
rect 14904 6544 14960 6578
rect 14994 6544 15050 6578
rect 15084 6544 15140 6578
rect 15174 6544 15230 6578
rect 15264 6544 15320 6578
rect 15354 6544 15413 6578
rect 14719 6530 15413 6544
rect 14719 6496 14792 6530
rect 14826 6496 14892 6530
rect 14926 6496 14992 6530
rect 15026 6496 15092 6530
rect 15126 6496 15192 6530
rect 15226 6496 15292 6530
rect 15326 6496 15413 6530
rect 14719 6488 15413 6496
rect 14719 6454 14780 6488
rect 14814 6454 14870 6488
rect 14904 6454 14960 6488
rect 14994 6454 15050 6488
rect 15084 6454 15140 6488
rect 15174 6454 15230 6488
rect 15264 6454 15320 6488
rect 15354 6454 15413 6488
rect 14719 6430 15413 6454
rect 14719 6398 14792 6430
rect 14826 6398 14892 6430
rect 14926 6398 14992 6430
rect 15026 6398 15092 6430
rect 14719 6364 14780 6398
rect 14826 6396 14870 6398
rect 14926 6396 14960 6398
rect 15026 6396 15050 6398
rect 14814 6364 14870 6396
rect 14904 6364 14960 6396
rect 14994 6364 15050 6396
rect 15084 6396 15092 6398
rect 15126 6398 15192 6430
rect 15126 6396 15140 6398
rect 15084 6364 15140 6396
rect 15174 6396 15192 6398
rect 15226 6398 15292 6430
rect 15326 6398 15413 6430
rect 15226 6396 15230 6398
rect 15174 6364 15230 6396
rect 15264 6396 15292 6398
rect 15264 6364 15320 6396
rect 15354 6364 15413 6398
rect 14719 6330 15413 6364
rect 14719 6308 14792 6330
rect 14826 6308 14892 6330
rect 14926 6308 14992 6330
rect 15026 6308 15092 6330
rect 14719 6274 14780 6308
rect 14826 6296 14870 6308
rect 14926 6296 14960 6308
rect 15026 6296 15050 6308
rect 14814 6274 14870 6296
rect 14904 6274 14960 6296
rect 14994 6274 15050 6296
rect 15084 6296 15092 6308
rect 15126 6308 15192 6330
rect 15126 6296 15140 6308
rect 15084 6274 15140 6296
rect 15174 6296 15192 6308
rect 15226 6308 15292 6330
rect 15326 6308 15413 6330
rect 15226 6296 15230 6308
rect 15174 6274 15230 6296
rect 15264 6296 15292 6308
rect 15264 6274 15320 6296
rect 15354 6274 15413 6308
rect 14719 6230 15413 6274
rect 14719 6218 14792 6230
rect 14826 6218 14892 6230
rect 14926 6218 14992 6230
rect 15026 6218 15092 6230
rect 14719 6184 14780 6218
rect 14826 6196 14870 6218
rect 14926 6196 14960 6218
rect 15026 6196 15050 6218
rect 14814 6184 14870 6196
rect 14904 6184 14960 6196
rect 14994 6184 15050 6196
rect 15084 6196 15092 6218
rect 15126 6218 15192 6230
rect 15126 6196 15140 6218
rect 15084 6184 15140 6196
rect 15174 6196 15192 6218
rect 15226 6218 15292 6230
rect 15326 6218 15413 6230
rect 15226 6196 15230 6218
rect 15174 6184 15230 6196
rect 15264 6196 15292 6218
rect 15264 6184 15320 6196
rect 15354 6184 15413 6218
rect 14719 6123 15413 6184
rect 15475 6766 15547 6822
rect 15475 6732 15494 6766
rect 15528 6732 15547 6766
rect 15475 6676 15547 6732
rect 15475 6642 15494 6676
rect 15528 6642 15547 6676
rect 15475 6586 15547 6642
rect 15475 6552 15494 6586
rect 15528 6552 15547 6586
rect 15475 6496 15547 6552
rect 15475 6462 15494 6496
rect 15528 6462 15547 6496
rect 15475 6406 15547 6462
rect 15475 6372 15494 6406
rect 15528 6372 15547 6406
rect 15475 6316 15547 6372
rect 15475 6282 15494 6316
rect 15528 6282 15547 6316
rect 15475 6226 15547 6282
rect 15475 6192 15494 6226
rect 15528 6192 15547 6226
rect 15475 6136 15547 6192
rect 14585 6061 14657 6121
rect 15475 6102 15494 6136
rect 15528 6102 15547 6136
rect 15475 6061 15547 6102
rect 14585 6060 15547 6061
rect 14406 5976 14521 6032
rect 14406 5942 14456 5976
rect 14490 5942 14521 5976
rect 14406 5925 14521 5942
rect 14566 6042 15547 6060
rect 14566 6008 14682 6042
rect 14716 6008 14772 6042
rect 14806 6008 14862 6042
rect 14896 6008 14952 6042
rect 14986 6008 15042 6042
rect 15076 6008 15132 6042
rect 15166 6008 15222 6042
rect 15256 6008 15312 6042
rect 15346 6008 15402 6042
rect 15436 6008 15547 6042
rect 14566 5989 15547 6008
rect 15611 6932 15643 6966
rect 15677 6932 15710 6966
rect 15611 6876 15710 6932
rect 15611 6842 15643 6876
rect 15677 6842 15710 6876
rect 15611 6786 15710 6842
rect 15611 6752 15643 6786
rect 15677 6752 15710 6786
rect 15611 6696 15710 6752
rect 15611 6662 15643 6696
rect 15677 6662 15710 6696
rect 15611 6606 15710 6662
rect 15611 6572 15643 6606
rect 15677 6572 15710 6606
rect 15611 6516 15710 6572
rect 15611 6482 15643 6516
rect 15677 6482 15710 6516
rect 15611 6426 15710 6482
rect 15611 6392 15643 6426
rect 15677 6392 15710 6426
rect 15611 6336 15710 6392
rect 15611 6302 15643 6336
rect 15677 6302 15710 6336
rect 15611 6246 15710 6302
rect 15611 6212 15643 6246
rect 15677 6212 15710 6246
rect 15611 6156 15710 6212
rect 15611 6122 15643 6156
rect 15677 6122 15710 6156
rect 15611 6066 15710 6122
rect 15611 6032 15643 6066
rect 15677 6032 15710 6066
rect 14566 5925 15526 5989
rect 15611 5976 15710 6032
rect 15611 5942 15643 5976
rect 15677 5942 15710 5976
rect 15611 5925 15710 5942
rect 14406 5892 15710 5925
rect 14406 5858 14552 5892
rect 14586 5858 14642 5892
rect 14676 5858 14732 5892
rect 14766 5858 14822 5892
rect 14856 5858 14912 5892
rect 14946 5858 15002 5892
rect 15036 5858 15092 5892
rect 15126 5858 15182 5892
rect 15216 5858 15272 5892
rect 15306 5858 15362 5892
rect 15396 5858 15452 5892
rect 15486 5858 15542 5892
rect 15576 5858 15710 5892
rect 14406 5826 15710 5858
rect 17012 7119 17046 7206
rect 16114 7085 16210 7104
rect 16080 7051 16210 7085
rect 16114 7017 16210 7051
rect 16080 6983 16210 7017
rect 16114 6949 16210 6983
rect 16080 6915 16210 6949
rect 16114 6881 16210 6915
rect 16080 6847 16210 6881
rect 16114 6813 16210 6847
rect 16080 6779 16210 6813
rect 16114 6745 16210 6779
rect 16080 6711 16210 6745
rect 16114 6678 16210 6711
rect 16842 6678 16846 7102
rect 16916 7085 17012 7102
rect 16916 7051 17046 7085
rect 16916 7017 17012 7051
rect 16916 6983 17046 7017
rect 16916 6949 17012 6983
rect 16916 6915 17046 6949
rect 16916 6881 17012 6915
rect 16916 6847 17046 6881
rect 16916 6813 17012 6847
rect 16916 6779 17046 6813
rect 16916 6745 17012 6779
rect 16916 6711 17046 6745
rect 16916 6678 17012 6711
rect 16114 6677 16280 6678
rect 16080 6666 16280 6677
rect 16842 6677 17012 6678
rect 16080 6643 16114 6666
rect 16842 6664 17046 6677
rect 16080 6575 16114 6609
rect 16080 6507 16114 6541
rect 16080 6439 16114 6473
rect 16080 6371 16114 6405
rect 16080 6303 16114 6337
rect 16080 6235 16114 6269
rect 16080 6167 16114 6201
rect 16080 6099 16114 6133
rect 16080 6031 16114 6065
rect 16080 5963 16114 5997
rect 16080 5895 16114 5929
rect 16080 5827 16114 5861
rect 12756 5734 12856 5796
rect 12916 5780 13876 5796
rect 14406 5754 14506 5826
rect 14566 5810 15526 5826
rect 16080 5759 16114 5793
rect 12756 5699 14060 5734
rect 12756 5676 12902 5699
rect 12756 5642 12806 5676
rect 12840 5665 12902 5676
rect 12936 5665 12992 5699
rect 13026 5665 13082 5699
rect 13116 5665 13172 5699
rect 13206 5665 13262 5699
rect 13296 5665 13352 5699
rect 13386 5665 13442 5699
rect 13476 5665 13532 5699
rect 13566 5665 13622 5699
rect 13656 5665 13712 5699
rect 13746 5665 13802 5699
rect 13836 5665 13892 5699
rect 13926 5676 14060 5699
rect 13926 5665 13993 5676
rect 12840 5642 13993 5665
rect 14027 5642 14060 5676
rect 12756 5635 14060 5642
rect 12756 5586 12871 5635
rect 12756 5552 12806 5586
rect 12840 5552 12871 5586
rect 13961 5586 14060 5635
rect 12756 5496 12871 5552
rect 12756 5462 12806 5496
rect 12840 5462 12871 5496
rect 12756 5406 12871 5462
rect 12756 5372 12806 5406
rect 12840 5372 12871 5406
rect 12756 5316 12871 5372
rect -7992 5279 -3406 5289
rect -7992 5245 -7773 5279
rect -7739 5245 -7705 5279
rect -7671 5245 -7637 5279
rect -7603 5245 -7569 5279
rect -7535 5245 -7501 5279
rect -7467 5245 -7433 5279
rect -7399 5245 -7365 5279
rect -7331 5245 -7297 5279
rect -7263 5245 -7229 5279
rect -7195 5245 -7161 5279
rect -7127 5245 -7093 5279
rect -7059 5245 -7025 5279
rect -6991 5245 -6957 5279
rect -6923 5245 -6889 5279
rect -6855 5245 -6821 5279
rect -6787 5245 -6753 5279
rect -6719 5245 -6685 5279
rect -6651 5245 -6617 5279
rect -6583 5245 -6549 5279
rect -6515 5245 -6481 5279
rect -6447 5245 -6413 5279
rect -6379 5245 -6345 5279
rect -6311 5245 -6277 5279
rect -6243 5245 -6209 5279
rect -6175 5245 -6141 5279
rect -6107 5245 -6073 5279
rect -6039 5245 -6005 5279
rect -5971 5245 -5937 5279
rect -5903 5245 -5869 5279
rect -5835 5245 -5801 5279
rect -5767 5245 -5733 5279
rect -5699 5245 -5665 5279
rect -5631 5245 -5597 5279
rect -5563 5245 -5529 5279
rect -5495 5245 -5461 5279
rect -5427 5245 -5393 5279
rect -5359 5245 -5325 5279
rect -5291 5245 -5257 5279
rect -5223 5245 -5189 5279
rect -5155 5245 -5121 5279
rect -5087 5245 -5053 5279
rect -5019 5245 -4985 5279
rect -4951 5245 -4917 5279
rect -4883 5245 -4849 5279
rect -4815 5245 -4781 5279
rect -4747 5245 -4713 5279
rect -4679 5245 -4645 5279
rect -4611 5245 -4577 5279
rect -4543 5245 -4509 5279
rect -4475 5245 -4441 5279
rect -4407 5245 -4373 5279
rect -4339 5245 -4305 5279
rect -4271 5245 -4237 5279
rect -4203 5245 -4169 5279
rect -4135 5245 -4101 5279
rect -4067 5245 -4033 5279
rect -3999 5245 -3965 5279
rect -3931 5245 -3897 5279
rect -3863 5245 -3829 5279
rect -3795 5245 -3761 5279
rect -3727 5245 -3693 5279
rect -3659 5245 -3625 5279
rect -3591 5245 -3406 5279
rect -7992 5011 -3406 5245
rect 12756 5282 12806 5316
rect 12840 5282 12871 5316
rect 12756 5226 12871 5282
rect 12756 5192 12806 5226
rect 12840 5192 12871 5226
rect 12756 5136 12871 5192
rect 12756 5102 12806 5136
rect 12840 5102 12871 5136
rect 12756 5046 12871 5102
rect 12756 5012 12806 5046
rect 12840 5012 12871 5046
rect -8298 4213 -3006 5011
rect 12756 4956 12871 5012
rect 12756 4922 12806 4956
rect 12840 4922 12871 4956
rect 12756 4866 12871 4922
rect 12756 4832 12806 4866
rect 12840 4832 12871 4866
rect 12756 4776 12871 4832
rect 12756 4742 12806 4776
rect 12840 4742 12871 4776
rect 12756 4686 12871 4742
rect 12935 5552 13897 5571
rect 12935 5518 13066 5552
rect 13100 5518 13156 5552
rect 13190 5518 13246 5552
rect 13280 5518 13336 5552
rect 13370 5518 13426 5552
rect 13460 5518 13516 5552
rect 13550 5518 13606 5552
rect 13640 5518 13696 5552
rect 13730 5518 13786 5552
rect 13820 5518 13897 5552
rect 12935 5499 13897 5518
rect 12935 5495 13007 5499
rect 12935 5461 12954 5495
rect 12988 5461 13007 5495
rect 12935 5405 13007 5461
rect 13825 5476 13897 5499
rect 13825 5442 13844 5476
rect 13878 5442 13897 5476
rect 12935 5371 12954 5405
rect 12988 5371 13007 5405
rect 12935 5315 13007 5371
rect 12935 5281 12954 5315
rect 12988 5281 13007 5315
rect 12935 5225 13007 5281
rect 12935 5191 12954 5225
rect 12988 5191 13007 5225
rect 12935 5135 13007 5191
rect 12935 5101 12954 5135
rect 12988 5101 13007 5135
rect 12935 5045 13007 5101
rect 12935 5011 12954 5045
rect 12988 5011 13007 5045
rect 12935 4955 13007 5011
rect 12935 4921 12954 4955
rect 12988 4921 13007 4955
rect 12935 4865 13007 4921
rect 12935 4831 12954 4865
rect 12988 4831 13007 4865
rect 12935 4775 13007 4831
rect 12935 4741 12954 4775
rect 12988 4741 13007 4775
rect 13069 5378 13763 5437
rect 13069 5344 13130 5378
rect 13164 5350 13220 5378
rect 13254 5350 13310 5378
rect 13344 5350 13400 5378
rect 13176 5344 13220 5350
rect 13276 5344 13310 5350
rect 13376 5344 13400 5350
rect 13434 5350 13490 5378
rect 13434 5344 13442 5350
rect 13069 5316 13142 5344
rect 13176 5316 13242 5344
rect 13276 5316 13342 5344
rect 13376 5316 13442 5344
rect 13476 5344 13490 5350
rect 13524 5350 13580 5378
rect 13524 5344 13542 5350
rect 13476 5316 13542 5344
rect 13576 5344 13580 5350
rect 13614 5350 13670 5378
rect 13614 5344 13642 5350
rect 13704 5344 13763 5378
rect 13576 5316 13642 5344
rect 13676 5316 13763 5344
rect 13069 5288 13763 5316
rect 13069 5254 13130 5288
rect 13164 5254 13220 5288
rect 13254 5254 13310 5288
rect 13344 5254 13400 5288
rect 13434 5254 13490 5288
rect 13524 5254 13580 5288
rect 13614 5254 13670 5288
rect 13704 5254 13763 5288
rect 13069 5250 13763 5254
rect 13069 5216 13142 5250
rect 13176 5216 13242 5250
rect 13276 5216 13342 5250
rect 13376 5216 13442 5250
rect 13476 5216 13542 5250
rect 13576 5216 13642 5250
rect 13676 5216 13763 5250
rect 13069 5198 13763 5216
rect 13069 5164 13130 5198
rect 13164 5164 13220 5198
rect 13254 5164 13310 5198
rect 13344 5164 13400 5198
rect 13434 5164 13490 5198
rect 13524 5164 13580 5198
rect 13614 5164 13670 5198
rect 13704 5164 13763 5198
rect 13069 5150 13763 5164
rect 13069 5116 13142 5150
rect 13176 5116 13242 5150
rect 13276 5116 13342 5150
rect 13376 5116 13442 5150
rect 13476 5116 13542 5150
rect 13576 5116 13642 5150
rect 13676 5116 13763 5150
rect 13069 5108 13763 5116
rect 13069 5074 13130 5108
rect 13164 5074 13220 5108
rect 13254 5074 13310 5108
rect 13344 5074 13400 5108
rect 13434 5074 13490 5108
rect 13524 5074 13580 5108
rect 13614 5074 13670 5108
rect 13704 5074 13763 5108
rect 13069 5050 13763 5074
rect 13069 5018 13142 5050
rect 13176 5018 13242 5050
rect 13276 5018 13342 5050
rect 13376 5018 13442 5050
rect 13069 4984 13130 5018
rect 13176 5016 13220 5018
rect 13276 5016 13310 5018
rect 13376 5016 13400 5018
rect 13164 4984 13220 5016
rect 13254 4984 13310 5016
rect 13344 4984 13400 5016
rect 13434 5016 13442 5018
rect 13476 5018 13542 5050
rect 13476 5016 13490 5018
rect 13434 4984 13490 5016
rect 13524 5016 13542 5018
rect 13576 5018 13642 5050
rect 13676 5018 13763 5050
rect 13576 5016 13580 5018
rect 13524 4984 13580 5016
rect 13614 5016 13642 5018
rect 13614 4984 13670 5016
rect 13704 4984 13763 5018
rect 13069 4950 13763 4984
rect 13069 4928 13142 4950
rect 13176 4928 13242 4950
rect 13276 4928 13342 4950
rect 13376 4928 13442 4950
rect 13069 4894 13130 4928
rect 13176 4916 13220 4928
rect 13276 4916 13310 4928
rect 13376 4916 13400 4928
rect 13164 4894 13220 4916
rect 13254 4894 13310 4916
rect 13344 4894 13400 4916
rect 13434 4916 13442 4928
rect 13476 4928 13542 4950
rect 13476 4916 13490 4928
rect 13434 4894 13490 4916
rect 13524 4916 13542 4928
rect 13576 4928 13642 4950
rect 13676 4928 13763 4950
rect 13576 4916 13580 4928
rect 13524 4894 13580 4916
rect 13614 4916 13642 4928
rect 13614 4894 13670 4916
rect 13704 4894 13763 4928
rect 13069 4850 13763 4894
rect 13069 4838 13142 4850
rect 13176 4838 13242 4850
rect 13276 4838 13342 4850
rect 13376 4838 13442 4850
rect 13069 4804 13130 4838
rect 13176 4816 13220 4838
rect 13276 4816 13310 4838
rect 13376 4816 13400 4838
rect 13164 4804 13220 4816
rect 13254 4804 13310 4816
rect 13344 4804 13400 4816
rect 13434 4816 13442 4838
rect 13476 4838 13542 4850
rect 13476 4816 13490 4838
rect 13434 4804 13490 4816
rect 13524 4816 13542 4838
rect 13576 4838 13642 4850
rect 13676 4838 13763 4850
rect 13576 4816 13580 4838
rect 13524 4804 13580 4816
rect 13614 4816 13642 4838
rect 13614 4804 13670 4816
rect 13704 4804 13763 4838
rect 13069 4743 13763 4804
rect 13825 5386 13897 5442
rect 13825 5352 13844 5386
rect 13878 5352 13897 5386
rect 13825 5296 13897 5352
rect 13825 5262 13844 5296
rect 13878 5262 13897 5296
rect 13825 5206 13897 5262
rect 13825 5172 13844 5206
rect 13878 5172 13897 5206
rect 13825 5116 13897 5172
rect 13825 5082 13844 5116
rect 13878 5082 13897 5116
rect 13825 5026 13897 5082
rect 13825 4992 13844 5026
rect 13878 4992 13897 5026
rect 13825 4936 13897 4992
rect 13825 4902 13844 4936
rect 13878 4902 13897 4936
rect 13825 4846 13897 4902
rect 13825 4812 13844 4846
rect 13878 4812 13897 4846
rect 13825 4756 13897 4812
rect 12935 4691 13007 4741
rect 13825 4722 13844 4756
rect 13878 4722 13897 4756
rect 13825 4691 13897 4722
rect 12756 4652 12806 4686
rect 12840 4652 12871 4686
rect 12756 4596 12871 4652
rect 12756 4562 12806 4596
rect 12840 4562 12871 4596
rect 12756 4560 12871 4562
rect 12916 4662 13897 4691
rect 12916 4628 13032 4662
rect 13066 4628 13122 4662
rect 13156 4628 13212 4662
rect 13246 4628 13302 4662
rect 13336 4628 13392 4662
rect 13426 4628 13482 4662
rect 13516 4628 13572 4662
rect 13606 4628 13662 4662
rect 13696 4628 13752 4662
rect 13786 4628 13897 4662
rect 12916 4609 13897 4628
rect 13961 5552 13993 5586
rect 14027 5552 14060 5586
rect 13961 5496 14060 5552
rect 13961 5462 13993 5496
rect 14027 5462 14060 5496
rect 13961 5406 14060 5462
rect 13961 5372 13993 5406
rect 14027 5372 14060 5406
rect 13961 5316 14060 5372
rect 13961 5282 13993 5316
rect 14027 5282 14060 5316
rect 13961 5226 14060 5282
rect 13961 5192 13993 5226
rect 14027 5192 14060 5226
rect 13961 5136 14060 5192
rect 13961 5102 13993 5136
rect 14027 5102 14060 5136
rect 13961 5046 14060 5102
rect 13961 5012 13993 5046
rect 14027 5012 14060 5046
rect 13961 4956 14060 5012
rect 13961 4922 13993 4956
rect 14027 4922 14060 4956
rect 13961 4866 14060 4922
rect 13961 4832 13993 4866
rect 14027 4832 14060 4866
rect 13961 4776 14060 4832
rect 13961 4742 13993 4776
rect 14027 4742 14060 4776
rect 13961 4686 14060 4742
rect 13961 4652 13993 4686
rect 14027 4652 14060 4686
rect 12916 4560 13876 4609
rect 13961 4596 14060 4652
rect 13961 4562 13993 4596
rect 14027 4562 14060 4596
rect 13961 4560 14060 4562
rect 14406 5719 15710 5754
rect 14406 5696 14552 5719
rect 14406 5662 14456 5696
rect 14490 5685 14552 5696
rect 14586 5685 14642 5719
rect 14676 5685 14732 5719
rect 14766 5685 14822 5719
rect 14856 5685 14912 5719
rect 14946 5685 15002 5719
rect 15036 5685 15092 5719
rect 15126 5685 15182 5719
rect 15216 5685 15272 5719
rect 15306 5685 15362 5719
rect 15396 5685 15452 5719
rect 15486 5685 15542 5719
rect 15576 5696 15710 5719
rect 15576 5685 15643 5696
rect 14490 5662 15643 5685
rect 15677 5662 15710 5696
rect 14406 5655 15710 5662
rect 14406 5606 14521 5655
rect 14406 5572 14456 5606
rect 14490 5572 14521 5606
rect 15611 5606 15710 5655
rect 14406 5516 14521 5572
rect 14406 5482 14456 5516
rect 14490 5482 14521 5516
rect 14406 5426 14521 5482
rect 14406 5392 14456 5426
rect 14490 5392 14521 5426
rect 14406 5336 14521 5392
rect 14406 5302 14456 5336
rect 14490 5302 14521 5336
rect 14406 5246 14521 5302
rect 14406 5212 14456 5246
rect 14490 5212 14521 5246
rect 14406 5156 14521 5212
rect 14406 5122 14456 5156
rect 14490 5122 14521 5156
rect 14406 5066 14521 5122
rect 14406 5032 14456 5066
rect 14490 5032 14521 5066
rect 14406 4976 14521 5032
rect 14406 4942 14456 4976
rect 14490 4942 14521 4976
rect 14406 4886 14521 4942
rect 14406 4852 14456 4886
rect 14490 4852 14521 4886
rect 14406 4796 14521 4852
rect 14406 4762 14456 4796
rect 14490 4762 14521 4796
rect 14406 4706 14521 4762
rect 14406 4672 14456 4706
rect 14490 4672 14521 4706
rect 14585 5572 15547 5591
rect 14585 5538 14716 5572
rect 14750 5538 14806 5572
rect 14840 5538 14896 5572
rect 14930 5538 14986 5572
rect 15020 5538 15076 5572
rect 15110 5538 15166 5572
rect 15200 5538 15256 5572
rect 15290 5538 15346 5572
rect 15380 5538 15436 5572
rect 15470 5538 15547 5572
rect 14585 5519 15547 5538
rect 14585 5515 14657 5519
rect 14585 5481 14604 5515
rect 14638 5481 14657 5515
rect 14585 5425 14657 5481
rect 15475 5496 15547 5519
rect 15475 5462 15494 5496
rect 15528 5462 15547 5496
rect 14585 5391 14604 5425
rect 14638 5391 14657 5425
rect 14585 5335 14657 5391
rect 14585 5301 14604 5335
rect 14638 5301 14657 5335
rect 14585 5245 14657 5301
rect 14585 5211 14604 5245
rect 14638 5211 14657 5245
rect 14585 5155 14657 5211
rect 14585 5121 14604 5155
rect 14638 5121 14657 5155
rect 14585 5065 14657 5121
rect 14585 5031 14604 5065
rect 14638 5031 14657 5065
rect 14585 4975 14657 5031
rect 14585 4941 14604 4975
rect 14638 4941 14657 4975
rect 14585 4885 14657 4941
rect 14585 4851 14604 4885
rect 14638 4851 14657 4885
rect 14585 4795 14657 4851
rect 14585 4761 14604 4795
rect 14638 4761 14657 4795
rect 14719 5398 15413 5457
rect 14719 5364 14780 5398
rect 14814 5370 14870 5398
rect 14904 5370 14960 5398
rect 14994 5370 15050 5398
rect 14826 5364 14870 5370
rect 14926 5364 14960 5370
rect 15026 5364 15050 5370
rect 15084 5370 15140 5398
rect 15084 5364 15092 5370
rect 14719 5336 14792 5364
rect 14826 5336 14892 5364
rect 14926 5336 14992 5364
rect 15026 5336 15092 5364
rect 15126 5364 15140 5370
rect 15174 5370 15230 5398
rect 15174 5364 15192 5370
rect 15126 5336 15192 5364
rect 15226 5364 15230 5370
rect 15264 5370 15320 5398
rect 15264 5364 15292 5370
rect 15354 5364 15413 5398
rect 15226 5336 15292 5364
rect 15326 5336 15413 5364
rect 14719 5308 15413 5336
rect 14719 5274 14780 5308
rect 14814 5274 14870 5308
rect 14904 5274 14960 5308
rect 14994 5274 15050 5308
rect 15084 5274 15140 5308
rect 15174 5274 15230 5308
rect 15264 5274 15320 5308
rect 15354 5274 15413 5308
rect 14719 5270 15413 5274
rect 14719 5236 14792 5270
rect 14826 5236 14892 5270
rect 14926 5236 14992 5270
rect 15026 5236 15092 5270
rect 15126 5236 15192 5270
rect 15226 5236 15292 5270
rect 15326 5236 15413 5270
rect 14719 5218 15413 5236
rect 14719 5184 14780 5218
rect 14814 5184 14870 5218
rect 14904 5184 14960 5218
rect 14994 5184 15050 5218
rect 15084 5184 15140 5218
rect 15174 5184 15230 5218
rect 15264 5184 15320 5218
rect 15354 5184 15413 5218
rect 14719 5170 15413 5184
rect 14719 5136 14792 5170
rect 14826 5136 14892 5170
rect 14926 5136 14992 5170
rect 15026 5136 15092 5170
rect 15126 5136 15192 5170
rect 15226 5136 15292 5170
rect 15326 5136 15413 5170
rect 14719 5128 15413 5136
rect 14719 5094 14780 5128
rect 14814 5094 14870 5128
rect 14904 5094 14960 5128
rect 14994 5094 15050 5128
rect 15084 5094 15140 5128
rect 15174 5094 15230 5128
rect 15264 5094 15320 5128
rect 15354 5094 15413 5128
rect 14719 5070 15413 5094
rect 14719 5038 14792 5070
rect 14826 5038 14892 5070
rect 14926 5038 14992 5070
rect 15026 5038 15092 5070
rect 14719 5004 14780 5038
rect 14826 5036 14870 5038
rect 14926 5036 14960 5038
rect 15026 5036 15050 5038
rect 14814 5004 14870 5036
rect 14904 5004 14960 5036
rect 14994 5004 15050 5036
rect 15084 5036 15092 5038
rect 15126 5038 15192 5070
rect 15126 5036 15140 5038
rect 15084 5004 15140 5036
rect 15174 5036 15192 5038
rect 15226 5038 15292 5070
rect 15326 5038 15413 5070
rect 15226 5036 15230 5038
rect 15174 5004 15230 5036
rect 15264 5036 15292 5038
rect 15264 5004 15320 5036
rect 15354 5004 15413 5038
rect 14719 4970 15413 5004
rect 14719 4948 14792 4970
rect 14826 4948 14892 4970
rect 14926 4948 14992 4970
rect 15026 4948 15092 4970
rect 14719 4914 14780 4948
rect 14826 4936 14870 4948
rect 14926 4936 14960 4948
rect 15026 4936 15050 4948
rect 14814 4914 14870 4936
rect 14904 4914 14960 4936
rect 14994 4914 15050 4936
rect 15084 4936 15092 4948
rect 15126 4948 15192 4970
rect 15126 4936 15140 4948
rect 15084 4914 15140 4936
rect 15174 4936 15192 4948
rect 15226 4948 15292 4970
rect 15326 4948 15413 4970
rect 15226 4936 15230 4948
rect 15174 4914 15230 4936
rect 15264 4936 15292 4948
rect 15264 4914 15320 4936
rect 15354 4914 15413 4948
rect 14719 4870 15413 4914
rect 14719 4858 14792 4870
rect 14826 4858 14892 4870
rect 14926 4858 14992 4870
rect 15026 4858 15092 4870
rect 14719 4824 14780 4858
rect 14826 4836 14870 4858
rect 14926 4836 14960 4858
rect 15026 4836 15050 4858
rect 14814 4824 14870 4836
rect 14904 4824 14960 4836
rect 14994 4824 15050 4836
rect 15084 4836 15092 4858
rect 15126 4858 15192 4870
rect 15126 4836 15140 4858
rect 15084 4824 15140 4836
rect 15174 4836 15192 4858
rect 15226 4858 15292 4870
rect 15326 4858 15413 4870
rect 15226 4836 15230 4858
rect 15174 4824 15230 4836
rect 15264 4836 15292 4858
rect 15264 4824 15320 4836
rect 15354 4824 15413 4858
rect 14719 4763 15413 4824
rect 15475 5406 15547 5462
rect 15475 5372 15494 5406
rect 15528 5372 15547 5406
rect 15475 5316 15547 5372
rect 15475 5282 15494 5316
rect 15528 5282 15547 5316
rect 15475 5226 15547 5282
rect 15475 5192 15494 5226
rect 15528 5192 15547 5226
rect 15475 5136 15547 5192
rect 15475 5102 15494 5136
rect 15528 5102 15547 5136
rect 15475 5046 15547 5102
rect 15475 5012 15494 5046
rect 15528 5012 15547 5046
rect 15475 4956 15547 5012
rect 15475 4922 15494 4956
rect 15528 4922 15547 4956
rect 15475 4866 15547 4922
rect 15475 4832 15494 4866
rect 15528 4832 15547 4866
rect 15475 4776 15547 4832
rect 14585 4701 14657 4761
rect 15475 4742 15494 4776
rect 15528 4742 15547 4776
rect 15475 4701 15547 4742
rect 14585 4682 15547 4701
rect 14585 4680 14682 4682
rect 14406 4616 14521 4672
rect 14406 4582 14456 4616
rect 14490 4582 14521 4616
rect 14406 4565 14521 4582
rect 14566 4648 14682 4680
rect 14716 4648 14772 4682
rect 14806 4648 14862 4682
rect 14896 4648 14952 4682
rect 14986 4648 15042 4682
rect 15076 4648 15132 4682
rect 15166 4648 15222 4682
rect 15256 4648 15312 4682
rect 15346 4648 15402 4682
rect 15436 4648 15547 4682
rect 14566 4629 15547 4648
rect 15611 5572 15643 5606
rect 15677 5572 15710 5606
rect 15611 5516 15710 5572
rect 15611 5482 15643 5516
rect 15677 5482 15710 5516
rect 15611 5426 15710 5482
rect 15611 5392 15643 5426
rect 15677 5392 15710 5426
rect 15611 5336 15710 5392
rect 15611 5302 15643 5336
rect 15677 5302 15710 5336
rect 15611 5246 15710 5302
rect 15611 5212 15643 5246
rect 15677 5212 15710 5246
rect 15611 5156 15710 5212
rect 15611 5122 15643 5156
rect 15677 5122 15710 5156
rect 15611 5066 15710 5122
rect 15611 5032 15643 5066
rect 15677 5032 15710 5066
rect 15611 4976 15710 5032
rect 15611 4942 15643 4976
rect 15677 4942 15710 4976
rect 15611 4886 15710 4942
rect 15611 4852 15643 4886
rect 15677 4852 15710 4886
rect 15611 4796 15710 4852
rect 15611 4762 15643 4796
rect 15677 4762 15710 4796
rect 15611 4706 15710 4762
rect 15611 4672 15643 4706
rect 15677 4672 15710 4706
rect 14566 4565 15526 4629
rect 15611 4616 15710 4672
rect 15611 4582 15643 4616
rect 15677 4582 15710 4616
rect 15611 4565 15710 4582
rect 14406 4560 15710 4565
rect 12756 4538 15710 4560
rect 16080 5691 16114 5725
rect 16080 5623 16114 5657
rect 16080 5555 16114 5589
rect 16080 5487 16114 5521
rect 16080 5419 16114 5453
rect 16080 5351 16114 5385
rect 16080 5283 16114 5317
rect 16080 5215 16114 5249
rect 16080 5147 16114 5181
rect 16080 5079 16114 5113
rect 17012 6643 17046 6664
rect 17012 6575 17046 6609
rect 17012 6507 17046 6541
rect 17012 6439 17046 6473
rect 17012 6371 17046 6405
rect 17012 6303 17046 6337
rect 17012 6235 17046 6269
rect 17012 6167 17046 6201
rect 17012 6099 17046 6133
rect 17012 6031 17046 6065
rect 17012 5963 17046 5997
rect 17012 5895 17046 5929
rect 17012 5827 17046 5861
rect 17012 5759 17046 5793
rect 17012 5691 17046 5725
rect 17012 5623 17046 5657
rect 17012 5555 17046 5589
rect 17012 5487 17046 5521
rect 17012 5419 17046 5453
rect 17012 5351 17046 5385
rect 17012 5283 17046 5317
rect 17012 5215 17046 5249
rect 17012 5147 17046 5181
rect 17012 5079 17046 5113
rect 16114 5045 16210 5072
rect 16080 5011 16210 5045
rect 16114 4977 16210 5011
rect 16080 4943 16210 4977
rect 16114 4909 16210 4943
rect 16080 4875 16210 4909
rect 16114 4841 16210 4875
rect 16080 4807 16210 4841
rect 16114 4773 16210 4807
rect 16080 4739 16210 4773
rect 16114 4705 16210 4739
rect 16080 4671 16210 4705
rect 16114 4646 16210 4671
rect 16844 4646 16846 5070
rect 16916 5045 17012 5070
rect 16916 5011 17046 5045
rect 16916 4977 17012 5011
rect 16916 4943 17046 4977
rect 16916 4909 17012 4943
rect 16916 4875 17046 4909
rect 16916 4841 17012 4875
rect 16916 4807 17046 4841
rect 16916 4773 17012 4807
rect 16916 4739 17046 4773
rect 16916 4705 17012 4739
rect 16916 4671 17046 4705
rect 16916 4646 17012 4671
rect 16114 4637 16280 4646
rect 16080 4634 16280 4637
rect 16844 4637 17012 4646
rect 16080 4550 16114 4634
rect 16844 4632 17046 4637
rect 17012 4550 17046 4632
rect 16080 4544 16206 4550
rect 16048 4538 16206 4544
rect 12747 4532 16206 4538
rect 12747 4512 14552 4532
rect 12747 4478 12902 4512
rect 12936 4478 12992 4512
rect 13026 4478 13082 4512
rect 13116 4478 13172 4512
rect 13206 4478 13262 4512
rect 13296 4478 13352 4512
rect 13386 4478 13442 4512
rect 13476 4478 13532 4512
rect 13566 4478 13622 4512
rect 13656 4478 13712 4512
rect 13746 4478 13802 4512
rect 13836 4478 13892 4512
rect 13926 4498 14552 4512
rect 14586 4498 14642 4532
rect 14676 4498 14732 4532
rect 14766 4498 14822 4532
rect 14856 4498 14912 4532
rect 14946 4498 15002 4532
rect 15036 4498 15092 4532
rect 15126 4498 15182 4532
rect 15216 4498 15272 4532
rect 15306 4498 15362 4532
rect 15396 4498 15452 4532
rect 15486 4498 15542 4532
rect 15576 4516 16206 4532
rect 16240 4516 16274 4550
rect 16308 4516 16342 4550
rect 16376 4516 16410 4550
rect 16444 4516 16478 4550
rect 16512 4516 16546 4550
rect 16580 4516 16614 4550
rect 16648 4516 16682 4550
rect 16716 4516 16750 4550
rect 16784 4516 16818 4550
rect 16852 4516 16886 4550
rect 16920 4544 17046 4550
rect 17300 7221 17334 7255
rect 17300 7153 17334 7187
rect 17300 7085 17334 7119
rect 17300 7017 17334 7051
rect 17300 6949 17334 6983
rect 17300 6881 17334 6915
rect 17300 6813 17334 6847
rect 17300 6745 17334 6779
rect 17300 6677 17334 6711
rect 17300 6609 17334 6643
rect 17300 6541 17334 6575
rect 17300 6473 17334 6507
rect 17300 6405 17334 6439
rect 17300 6337 17334 6371
rect 17300 6269 17334 6303
rect 17300 6201 17334 6235
rect 17300 6133 17334 6167
rect 17300 6065 17334 6099
rect 17300 5997 17334 6031
rect 17300 5929 17334 5963
rect 17300 5861 17334 5895
rect 17300 5793 17334 5827
rect 17300 5725 17334 5759
rect 17300 5657 17334 5691
rect 17300 5589 17334 5623
rect 17300 5521 17334 5555
rect 17300 5453 17334 5487
rect 17300 5385 17334 5419
rect 17300 5317 17334 5351
rect 17300 5249 17334 5283
rect 17300 5181 17334 5215
rect 17300 5113 17334 5147
rect 17300 5045 17334 5079
rect 17300 4977 17334 5011
rect 17300 4909 17334 4943
rect 17300 4841 17334 4875
rect 17300 4773 17334 4807
rect 17300 4705 17334 4739
rect 17300 4637 17334 4671
rect 17300 4569 17334 4603
rect 16920 4516 17062 4544
rect 15576 4498 17062 4516
rect 13926 4478 17062 4498
rect 12747 4408 17062 4478
rect 17434 7527 17468 7552
rect 17434 7459 17468 7471
rect 17434 7391 17468 7399
rect 17434 7323 17468 7327
rect 17434 7217 17468 7221
rect 17434 7145 17468 7153
rect 17434 7073 17468 7085
rect 17434 7001 17468 7017
rect 17434 6929 17468 6949
rect 17434 6857 17468 6881
rect 17434 6785 17468 6813
rect 17434 6713 17468 6745
rect 17434 6643 17468 6677
rect 17434 6575 17468 6607
rect 17434 6507 17468 6535
rect 17434 6439 17468 6463
rect 17434 6371 17468 6391
rect 17434 6303 17468 6319
rect 17434 6235 17468 6247
rect 17434 6167 17468 6175
rect 17434 6099 17468 6103
rect 17434 5993 17468 5997
rect 17434 5921 17468 5929
rect 17434 5849 17468 5861
rect 17434 5777 17468 5793
rect 17434 5705 17468 5725
rect 17434 5633 17468 5657
rect 17434 5561 17468 5589
rect 17434 5489 17468 5521
rect 17434 5419 17468 5453
rect 17434 5351 17468 5383
rect 17434 5283 17468 5311
rect 17434 5215 17468 5239
rect 17434 5147 17468 5167
rect 17434 5079 17468 5095
rect 17434 5011 17468 5023
rect 17434 4943 17468 4951
rect 17434 4875 17468 4879
rect 17434 4769 17468 4773
rect 17434 4697 17468 4705
rect 17434 4625 17468 4637
rect 17434 4544 17468 4569
rect 18492 7527 18526 7552
rect 18492 7459 18526 7471
rect 18492 7391 18526 7399
rect 18492 7323 18526 7327
rect 18492 7217 18526 7221
rect 18492 7145 18526 7153
rect 18492 7073 18526 7085
rect 18492 7001 18526 7017
rect 18492 6929 18526 6949
rect 18492 6857 18526 6881
rect 18492 6785 18526 6813
rect 18492 6713 18526 6745
rect 18492 6643 18526 6677
rect 18492 6575 18526 6607
rect 18492 6507 18526 6535
rect 18492 6439 18526 6463
rect 18492 6371 18526 6391
rect 18492 6303 18526 6319
rect 18492 6235 18526 6247
rect 18492 6167 18526 6175
rect 18492 6099 18526 6103
rect 18492 5993 18526 5997
rect 18492 5921 18526 5929
rect 18492 5849 18526 5861
rect 18492 5777 18526 5793
rect 18492 5705 18526 5725
rect 18492 5633 18526 5657
rect 18492 5561 18526 5589
rect 18492 5489 18526 5521
rect 18492 5419 18526 5453
rect 18492 5351 18526 5383
rect 18492 5283 18526 5311
rect 18492 5215 18526 5239
rect 18492 5147 18526 5167
rect 18492 5079 18526 5095
rect 18492 5011 18526 5023
rect 18492 4943 18526 4951
rect 18492 4875 18526 4879
rect 18492 4769 18526 4773
rect 18492 4697 18526 4705
rect 18492 4625 18526 4637
rect 18492 4544 18526 4569
rect 18626 7493 18660 7527
rect 18626 7425 18660 7459
rect 18626 7357 18660 7391
rect 18626 7289 18660 7323
rect 18626 7221 18660 7255
rect 18626 7153 18660 7187
rect 18626 7085 18660 7119
rect 18626 7017 18660 7051
rect 18626 6949 18660 6983
rect 18626 6881 18660 6915
rect 18626 6813 18660 6847
rect 18626 6745 18660 6779
rect 18626 6677 18660 6711
rect 18626 6609 18660 6643
rect 18626 6541 18660 6575
rect 18626 6473 18660 6507
rect 18626 6405 18660 6439
rect 18626 6337 18660 6371
rect 18626 6269 18660 6303
rect 18626 6201 18660 6235
rect 18626 6133 18660 6167
rect 18626 6065 18660 6099
rect 18626 5997 18660 6031
rect 18626 5929 18660 5963
rect 18626 5861 18660 5895
rect 18626 5793 18660 5827
rect 18626 5725 18660 5759
rect 18626 5657 18660 5691
rect 18626 5589 18660 5623
rect 18626 5521 18660 5555
rect 18626 5453 18660 5487
rect 18626 5385 18660 5419
rect 18626 5317 18660 5351
rect 18626 5249 18660 5283
rect 18626 5181 18660 5215
rect 18626 5113 18660 5147
rect 18626 5045 18660 5079
rect 18626 4977 18660 5011
rect 18626 4909 18660 4943
rect 18626 4841 18660 4875
rect 18626 4773 18660 4807
rect 18626 4705 18660 4739
rect 18626 4637 18660 4671
rect 18626 4569 18660 4603
rect 17300 4501 17334 4535
rect 17480 4476 17521 4510
rect 17565 4476 17589 4510
rect 17637 4476 17657 4510
rect 17709 4476 17725 4510
rect 17781 4476 17793 4510
rect 17853 4476 17861 4510
rect 17925 4476 17929 4510
rect 18031 4476 18035 4510
rect 18099 4476 18107 4510
rect 18167 4476 18179 4510
rect 18235 4476 18251 4510
rect 18303 4476 18323 4510
rect 18371 4476 18395 4510
rect 18439 4476 18480 4510
rect 18626 4501 18660 4535
rect 12747 4364 17170 4408
rect 17300 4372 17334 4467
rect 18626 4372 18660 4467
rect 12747 4352 17240 4364
rect 17300 4352 17419 4372
rect 12747 4338 17419 4352
rect 17453 4338 17487 4372
rect 17521 4338 17555 4372
rect 17589 4338 17623 4372
rect 17657 4338 17691 4372
rect 17725 4338 17759 4372
rect 17793 4338 17827 4372
rect 17861 4338 17895 4372
rect 17929 4338 17963 4372
rect 17997 4338 18031 4372
rect 18065 4338 18099 4372
rect 18133 4338 18167 4372
rect 18201 4338 18235 4372
rect 18269 4338 18303 4372
rect 18337 4338 18371 4372
rect 18405 4338 18439 4372
rect 18473 4338 18507 4372
rect 18541 4352 18660 4372
rect 18750 7724 18869 7758
rect 18903 7724 18937 7758
rect 18971 7724 19005 7758
rect 19039 7724 19073 7758
rect 19107 7724 19141 7758
rect 19175 7724 19209 7758
rect 19243 7724 19277 7758
rect 19311 7724 19345 7758
rect 19379 7724 19413 7758
rect 19447 7724 19481 7758
rect 19515 7724 19549 7758
rect 19583 7724 19617 7758
rect 19651 7724 19685 7758
rect 19719 7724 19753 7758
rect 19787 7724 19821 7758
rect 19855 7724 19889 7758
rect 19923 7724 19957 7758
rect 19991 7724 20110 7758
rect 18750 7629 18784 7724
rect 20076 7629 20110 7724
rect 18750 7561 18784 7595
rect 18930 7586 18971 7620
rect 19015 7586 19039 7620
rect 19087 7586 19107 7620
rect 19159 7586 19175 7620
rect 19231 7586 19243 7620
rect 19303 7586 19311 7620
rect 19375 7586 19379 7620
rect 19481 7586 19485 7620
rect 19549 7586 19557 7620
rect 19617 7586 19629 7620
rect 19685 7586 19701 7620
rect 19753 7586 19773 7620
rect 19821 7586 19845 7620
rect 19889 7586 19930 7620
rect 20076 7561 20110 7595
rect 18750 7493 18784 7527
rect 18750 7425 18784 7459
rect 18750 7357 18784 7391
rect 18750 7289 18784 7323
rect 18750 7221 18784 7255
rect 18750 7153 18784 7187
rect 18750 7085 18784 7119
rect 18750 7017 18784 7051
rect 18750 6949 18784 6983
rect 18750 6881 18784 6915
rect 18750 6813 18784 6847
rect 18750 6745 18784 6779
rect 18750 6677 18784 6711
rect 18750 6609 18784 6643
rect 18750 6541 18784 6575
rect 18750 6473 18784 6507
rect 18750 6405 18784 6439
rect 18750 6337 18784 6371
rect 18750 6269 18784 6303
rect 18750 6201 18784 6235
rect 18750 6133 18784 6167
rect 18750 6065 18784 6099
rect 18750 5997 18784 6031
rect 18750 5929 18784 5963
rect 18750 5861 18784 5895
rect 18750 5793 18784 5827
rect 18750 5725 18784 5759
rect 18750 5657 18784 5691
rect 18750 5589 18784 5623
rect 18750 5521 18784 5555
rect 18750 5453 18784 5487
rect 18750 5385 18784 5419
rect 18750 5317 18784 5351
rect 18750 5249 18784 5283
rect 18750 5181 18784 5215
rect 18750 5113 18784 5147
rect 18750 5045 18784 5079
rect 18750 4977 18784 5011
rect 18750 4909 18784 4943
rect 18750 4841 18784 4875
rect 18750 4773 18784 4807
rect 18750 4705 18784 4739
rect 18750 4637 18784 4671
rect 18750 4569 18784 4603
rect 18884 7527 18918 7552
rect 18884 7459 18918 7471
rect 18884 7391 18918 7399
rect 18884 7323 18918 7327
rect 18884 7217 18918 7221
rect 18884 7145 18918 7153
rect 18884 7073 18918 7085
rect 18884 7001 18918 7017
rect 18884 6929 18918 6949
rect 18884 6857 18918 6881
rect 18884 6785 18918 6813
rect 18884 6713 18918 6745
rect 18884 6643 18918 6677
rect 18884 6575 18918 6607
rect 18884 6507 18918 6535
rect 18884 6439 18918 6463
rect 18884 6371 18918 6391
rect 18884 6303 18918 6319
rect 18884 6235 18918 6247
rect 18884 6167 18918 6175
rect 18884 6099 18918 6103
rect 18884 5993 18918 5997
rect 18884 5921 18918 5929
rect 18884 5849 18918 5861
rect 18884 5777 18918 5793
rect 18884 5705 18918 5725
rect 18884 5633 18918 5657
rect 18884 5561 18918 5589
rect 18884 5489 18918 5521
rect 18884 5419 18918 5453
rect 18884 5351 18918 5383
rect 18884 5283 18918 5311
rect 18884 5215 18918 5239
rect 18884 5147 18918 5167
rect 18884 5079 18918 5095
rect 18884 5011 18918 5023
rect 18884 4943 18918 4951
rect 18884 4875 18918 4879
rect 18884 4769 18918 4773
rect 18884 4697 18918 4705
rect 18884 4625 18918 4637
rect 18884 4544 18918 4569
rect 19942 7527 19976 7552
rect 19942 7459 19976 7471
rect 19942 7391 19976 7399
rect 19942 7323 19976 7327
rect 19942 7217 19976 7221
rect 19942 7145 19976 7153
rect 19942 7073 19976 7085
rect 19942 7001 19976 7017
rect 19942 6929 19976 6949
rect 19942 6857 19976 6881
rect 19942 6785 19976 6813
rect 19942 6713 19976 6745
rect 19942 6643 19976 6677
rect 19942 6575 19976 6607
rect 19942 6507 19976 6535
rect 19942 6439 19976 6463
rect 19942 6371 19976 6391
rect 19942 6303 19976 6319
rect 19942 6235 19976 6247
rect 19942 6167 19976 6175
rect 19942 6099 19976 6103
rect 19942 5993 19976 5997
rect 19942 5921 19976 5929
rect 19942 5849 19976 5861
rect 19942 5777 19976 5793
rect 19942 5705 19976 5725
rect 19942 5633 19976 5657
rect 19942 5561 19976 5589
rect 19942 5489 19976 5521
rect 19942 5419 19976 5453
rect 19942 5351 19976 5383
rect 19942 5283 19976 5311
rect 19942 5215 19976 5239
rect 19942 5147 19976 5167
rect 19942 5079 19976 5095
rect 19942 5011 19976 5023
rect 19942 4943 19976 4951
rect 19942 4875 19976 4879
rect 19942 4769 19976 4773
rect 19942 4697 19976 4705
rect 19942 4625 19976 4637
rect 19942 4544 19976 4569
rect 20076 7493 20110 7527
rect 20076 7425 20110 7459
rect 20076 7357 20110 7391
rect 20076 7289 20110 7323
rect 20076 7221 20110 7255
rect 20076 7153 20110 7187
rect 20076 7085 20110 7119
rect 20076 7017 20110 7051
rect 20076 6949 20110 6983
rect 20076 6881 20110 6915
rect 20076 6813 20110 6847
rect 20076 6745 20110 6779
rect 20076 6677 20110 6711
rect 20076 6609 20110 6643
rect 20076 6541 20110 6575
rect 20076 6473 20110 6507
rect 20076 6405 20110 6439
rect 20076 6337 20110 6371
rect 20076 6269 20110 6303
rect 20076 6201 20110 6235
rect 20076 6133 20110 6167
rect 20076 6065 20110 6099
rect 20076 5997 20110 6031
rect 20076 5929 20110 5963
rect 20076 5861 20110 5895
rect 20076 5793 20110 5827
rect 20076 5725 20110 5759
rect 20076 5657 20110 5691
rect 20076 5589 20110 5623
rect 20076 5521 20110 5555
rect 20076 5453 20110 5487
rect 20076 5385 20110 5419
rect 20076 5317 20110 5351
rect 20076 5249 20110 5283
rect 20076 5181 20110 5215
rect 20076 5113 20110 5147
rect 20076 5045 20110 5079
rect 20076 4977 20110 5011
rect 20076 4909 20110 4943
rect 20076 4841 20110 4875
rect 20076 4773 20110 4807
rect 20076 4705 20110 4739
rect 20076 4637 20110 4671
rect 20076 4569 20110 4603
rect 20382 7742 20416 7776
rect 20382 7674 20416 7708
rect 20382 7606 20416 7640
rect 20382 7538 20416 7572
rect 20382 7470 20416 7504
rect 20382 7402 20416 7436
rect 20382 7334 20416 7368
rect 20382 7266 20416 7300
rect 20382 7198 20416 7232
rect 20382 7130 20416 7164
rect 20382 7062 20416 7096
rect 20382 6994 20416 7028
rect 20382 6926 20416 6960
rect 20382 6858 20416 6892
rect 20382 6790 20416 6824
rect 20382 6722 20416 6756
rect 20382 6654 20416 6688
rect 20382 6586 20416 6620
rect 20382 6518 20416 6552
rect 20382 6450 20416 6484
rect 20382 6382 20416 6416
rect 20382 6314 20416 6348
rect 20382 6246 20416 6280
rect 20382 6178 20416 6212
rect 20382 6110 20416 6144
rect 20382 6042 20416 6076
rect 20382 5974 20416 6008
rect 20382 5906 20416 5940
rect 20382 5838 20416 5872
rect 20382 5770 20416 5804
rect 20382 5702 20416 5736
rect 20382 5634 20416 5668
rect 20382 5566 20416 5600
rect 20382 5498 20416 5532
rect 20382 5430 20416 5464
rect 20382 5362 20416 5396
rect 20382 5294 20416 5328
rect 20382 5226 20416 5260
rect 20382 5160 20416 5192
rect 21666 14038 21670 14066
rect 21632 13998 21666 14032
rect 21632 13930 21666 13964
rect 21862 13922 22482 14952
rect 23110 15817 24398 15852
rect 23110 15794 23240 15817
rect 23110 15760 23144 15794
rect 23178 15783 23240 15794
rect 23274 15783 23330 15817
rect 23364 15783 23420 15817
rect 23454 15783 23510 15817
rect 23544 15783 23600 15817
rect 23634 15783 23690 15817
rect 23724 15783 23780 15817
rect 23814 15783 23870 15817
rect 23904 15783 23960 15817
rect 23994 15783 24050 15817
rect 24084 15783 24140 15817
rect 24174 15783 24230 15817
rect 24264 15794 24398 15817
rect 24264 15783 24331 15794
rect 23178 15760 24331 15783
rect 24365 15760 24398 15794
rect 23110 15753 24398 15760
rect 23110 15704 23209 15753
rect 23110 15670 23144 15704
rect 23178 15670 23209 15704
rect 24299 15704 24398 15753
rect 23110 15614 23209 15670
rect 23110 15580 23144 15614
rect 23178 15580 23209 15614
rect 23110 15524 23209 15580
rect 23110 15490 23144 15524
rect 23178 15490 23209 15524
rect 23110 15434 23209 15490
rect 23110 15400 23144 15434
rect 23178 15400 23209 15434
rect 23110 15344 23209 15400
rect 23110 15310 23144 15344
rect 23178 15310 23209 15344
rect 23110 15254 23209 15310
rect 23110 15220 23144 15254
rect 23178 15220 23209 15254
rect 23110 15164 23209 15220
rect 23110 15130 23144 15164
rect 23178 15130 23209 15164
rect 23110 15074 23209 15130
rect 23110 15040 23144 15074
rect 23178 15040 23209 15074
rect 23110 14984 23209 15040
rect 23110 14950 23144 14984
rect 23178 14950 23209 14984
rect 23110 14894 23209 14950
rect 23110 14860 23144 14894
rect 23178 14860 23209 14894
rect 23110 14804 23209 14860
rect 23110 14770 23144 14804
rect 23178 14770 23209 14804
rect 23110 14714 23209 14770
rect 23273 15670 24235 15689
rect 23273 15636 23404 15670
rect 23438 15636 23494 15670
rect 23528 15636 23584 15670
rect 23618 15636 23674 15670
rect 23708 15636 23764 15670
rect 23798 15636 23854 15670
rect 23888 15636 23944 15670
rect 23978 15636 24034 15670
rect 24068 15636 24124 15670
rect 24158 15636 24235 15670
rect 23273 15617 24235 15636
rect 23273 15613 23345 15617
rect 23273 15579 23292 15613
rect 23326 15579 23345 15613
rect 23273 15523 23345 15579
rect 24163 15594 24235 15617
rect 24163 15560 24182 15594
rect 24216 15560 24235 15594
rect 23273 15489 23292 15523
rect 23326 15489 23345 15523
rect 23273 15433 23345 15489
rect 23273 15399 23292 15433
rect 23326 15399 23345 15433
rect 23273 15343 23345 15399
rect 23273 15309 23292 15343
rect 23326 15309 23345 15343
rect 23273 15253 23345 15309
rect 23273 15219 23292 15253
rect 23326 15219 23345 15253
rect 23273 15163 23345 15219
rect 23273 15129 23292 15163
rect 23326 15129 23345 15163
rect 23273 15073 23345 15129
rect 23273 15039 23292 15073
rect 23326 15039 23345 15073
rect 23273 14983 23345 15039
rect 23273 14949 23292 14983
rect 23326 14949 23345 14983
rect 23273 14893 23345 14949
rect 23273 14859 23292 14893
rect 23326 14859 23345 14893
rect 23407 15496 24101 15555
rect 23407 15462 23468 15496
rect 23502 15468 23558 15496
rect 23592 15468 23648 15496
rect 23682 15468 23738 15496
rect 23514 15462 23558 15468
rect 23614 15462 23648 15468
rect 23714 15462 23738 15468
rect 23772 15468 23828 15496
rect 23772 15462 23780 15468
rect 23407 15434 23480 15462
rect 23514 15434 23580 15462
rect 23614 15434 23680 15462
rect 23714 15434 23780 15462
rect 23814 15462 23828 15468
rect 23862 15468 23918 15496
rect 23862 15462 23880 15468
rect 23814 15434 23880 15462
rect 23914 15462 23918 15468
rect 23952 15468 24008 15496
rect 23952 15462 23980 15468
rect 24042 15462 24101 15496
rect 23914 15434 23980 15462
rect 24014 15434 24101 15462
rect 23407 15406 24101 15434
rect 23407 15372 23468 15406
rect 23502 15372 23558 15406
rect 23592 15372 23648 15406
rect 23682 15372 23738 15406
rect 23772 15372 23828 15406
rect 23862 15372 23918 15406
rect 23952 15372 24008 15406
rect 24042 15372 24101 15406
rect 23407 15368 24101 15372
rect 23407 15334 23480 15368
rect 23514 15334 23580 15368
rect 23614 15334 23680 15368
rect 23714 15334 23780 15368
rect 23814 15334 23880 15368
rect 23914 15334 23980 15368
rect 24014 15334 24101 15368
rect 24163 15504 24235 15560
rect 24163 15470 24182 15504
rect 24216 15470 24235 15504
rect 24163 15414 24235 15470
rect 24163 15380 24182 15414
rect 24216 15380 24235 15414
rect 24163 15348 24235 15380
rect 24299 15670 24331 15704
rect 24365 15670 24398 15704
rect 24299 15614 24398 15670
rect 24299 15580 24331 15614
rect 24365 15580 24398 15614
rect 24299 15524 24398 15580
rect 24299 15490 24331 15524
rect 24365 15490 24398 15524
rect 24299 15434 24398 15490
rect 24299 15400 24331 15434
rect 24365 15400 24398 15434
rect 24299 15348 24398 15400
rect 24460 15830 24494 15864
rect 24460 15762 24494 15796
rect 24460 15694 24494 15728
rect 27650 15898 27684 15932
rect 27650 15830 27684 15864
rect 27650 15762 27684 15796
rect 27650 15694 27684 15728
rect 24460 15626 24494 15660
rect 27650 15626 27684 15660
rect 24460 15558 24494 15592
rect 24460 15490 24494 15524
rect 24460 15422 24494 15456
rect 27650 15558 27684 15592
rect 27650 15490 27684 15524
rect 27650 15422 27684 15456
rect 24460 15354 24494 15388
rect 23407 15316 24101 15334
rect 23407 15282 23468 15316
rect 23502 15282 23558 15316
rect 23592 15282 23648 15316
rect 23682 15282 23738 15316
rect 23772 15282 23828 15316
rect 23862 15282 23918 15316
rect 23952 15282 24008 15316
rect 24042 15282 24101 15316
rect 23407 15268 24101 15282
rect 23407 15234 23480 15268
rect 23514 15234 23580 15268
rect 23614 15234 23680 15268
rect 23714 15234 23780 15268
rect 23814 15234 23880 15268
rect 23914 15234 23980 15268
rect 24014 15234 24101 15268
rect 23407 15226 24101 15234
rect 23407 15192 23468 15226
rect 23502 15192 23558 15226
rect 23592 15192 23648 15226
rect 23682 15192 23738 15226
rect 23772 15192 23828 15226
rect 23862 15192 23918 15226
rect 23952 15192 24008 15226
rect 24042 15192 24101 15226
rect 23407 15168 24101 15192
rect 23407 15136 23480 15168
rect 23514 15136 23580 15168
rect 23614 15136 23680 15168
rect 23714 15136 23780 15168
rect 23407 15102 23468 15136
rect 23514 15134 23558 15136
rect 23614 15134 23648 15136
rect 23714 15134 23738 15136
rect 23502 15102 23558 15134
rect 23592 15102 23648 15134
rect 23682 15102 23738 15134
rect 23772 15134 23780 15136
rect 23814 15136 23880 15168
rect 23814 15134 23828 15136
rect 23772 15102 23828 15134
rect 23862 15134 23880 15136
rect 23914 15136 23980 15168
rect 24014 15136 24101 15168
rect 24162 15344 24460 15348
rect 24162 15324 24331 15344
rect 24162 15290 24182 15324
rect 24216 15310 24331 15324
rect 24365 15320 24460 15344
rect 27122 15388 27650 15390
rect 37706 16216 41165 16265
rect 37706 16182 37962 16216
rect 37996 16182 38030 16216
rect 38064 16182 38098 16216
rect 38132 16182 38166 16216
rect 38200 16182 38234 16216
rect 38268 16182 38302 16216
rect 38336 16182 38370 16216
rect 38404 16182 38438 16216
rect 38472 16182 38506 16216
rect 38540 16182 38574 16216
rect 38608 16182 38642 16216
rect 38676 16182 38710 16216
rect 38744 16182 38778 16216
rect 38812 16182 38846 16216
rect 38880 16182 38914 16216
rect 38948 16182 38982 16216
rect 39016 16182 39050 16216
rect 39084 16182 39118 16216
rect 39152 16182 39186 16216
rect 39220 16182 39254 16216
rect 39288 16182 39322 16216
rect 39356 16182 39390 16216
rect 39424 16182 39458 16216
rect 39492 16182 39526 16216
rect 39560 16182 39594 16216
rect 39628 16182 39662 16216
rect 39696 16182 39730 16216
rect 39764 16182 39798 16216
rect 39832 16182 39866 16216
rect 39900 16182 39934 16216
rect 39968 16182 40002 16216
rect 40036 16182 40070 16216
rect 40104 16182 40138 16216
rect 40172 16182 40206 16216
rect 40240 16182 40274 16216
rect 40308 16182 40342 16216
rect 40376 16182 40410 16216
rect 40444 16182 40478 16216
rect 40512 16182 40546 16216
rect 40580 16182 40614 16216
rect 40648 16182 40682 16216
rect 40716 16182 40750 16216
rect 40784 16182 40818 16216
rect 40852 16182 40886 16216
rect 40920 16182 41165 16216
rect 37706 16131 41165 16182
rect 37706 16058 37839 16131
rect 37706 16024 37749 16058
rect 37783 16024 37839 16058
rect 37706 15990 37839 16024
rect 37706 15956 37749 15990
rect 37783 15956 37839 15990
rect 41047 16018 41165 16131
rect 41047 15984 41089 16018
rect 41123 15984 41165 16018
rect 37706 15922 37839 15956
rect 37706 15888 37749 15922
rect 37783 15888 37839 15922
rect 37706 15854 37839 15888
rect 37706 15820 37749 15854
rect 37783 15820 37839 15854
rect 37706 15786 37839 15820
rect 37706 15752 37749 15786
rect 37783 15752 37839 15786
rect 37706 15718 37839 15752
rect 37706 15684 37749 15718
rect 37783 15684 37839 15718
rect 37706 15650 37839 15684
rect 38454 15913 38866 15962
rect 38454 15807 38517 15913
rect 38767 15807 38866 15913
rect 38454 15718 38866 15807
rect 38454 15684 38512 15718
rect 38546 15684 38772 15718
rect 38806 15684 38866 15718
rect 39497 15912 39895 15963
rect 39497 15806 39533 15912
rect 39855 15806 39895 15912
rect 39497 15731 39895 15806
rect 40531 15921 40679 15962
rect 40531 15887 40586 15921
rect 40620 15887 40679 15921
rect 40531 15849 40679 15887
rect 40531 15815 40586 15849
rect 40620 15815 40679 15849
rect 39497 15707 39896 15731
rect 38454 15652 38866 15684
rect 38903 15662 39463 15706
rect 37706 15616 37749 15650
rect 37783 15616 37839 15650
rect 37706 15582 37839 15616
rect 37706 15548 37749 15582
rect 37783 15548 37839 15582
rect 37706 15514 37839 15548
rect 37706 15480 37749 15514
rect 37783 15480 37839 15514
rect 37706 15446 37839 15480
rect 37706 15412 37749 15446
rect 37783 15412 37839 15446
rect 28834 15390 28960 15392
rect 27684 15388 28960 15390
rect 27122 15358 28960 15388
rect 28994 15358 29028 15392
rect 29062 15358 29096 15392
rect 29130 15358 29164 15392
rect 29198 15358 29232 15392
rect 29266 15358 29300 15392
rect 29334 15358 29368 15392
rect 29402 15358 29436 15392
rect 29470 15358 29504 15392
rect 29538 15358 29572 15392
rect 29606 15358 29640 15392
rect 29674 15358 29800 15392
rect 27122 15354 29040 15358
rect 27122 15348 27650 15354
rect 24494 15320 24590 15348
rect 24365 15310 24590 15320
rect 24216 15290 24590 15310
rect 24162 15286 24590 15290
rect 24162 15254 24460 15286
rect 24162 15234 24331 15254
rect 24162 15200 24182 15234
rect 24216 15220 24331 15234
rect 24365 15252 24460 15254
rect 24494 15278 24590 15286
rect 24494 15252 25022 15278
rect 24365 15220 25022 15252
rect 24216 15200 25022 15220
rect 24162 15182 25022 15200
rect 27554 15320 27650 15348
rect 27684 15320 29040 15354
rect 27554 15286 29040 15320
rect 27554 15278 27650 15286
rect 27122 15252 27650 15278
rect 27684 15275 29040 15286
rect 27684 15252 28834 15275
rect 27122 15241 28834 15252
rect 28868 15262 29040 15275
rect 29766 15275 29800 15358
rect 28868 15241 28964 15262
rect 27122 15207 28964 15241
rect 27122 15182 28834 15207
rect 24162 15164 24559 15182
rect 24162 15148 24331 15164
rect 23914 15134 23918 15136
rect 23862 15102 23918 15134
rect 23952 15134 23980 15136
rect 23952 15102 24008 15134
rect 24042 15102 24101 15136
rect 23407 15068 24101 15102
rect 23407 15046 23480 15068
rect 23514 15046 23580 15068
rect 23614 15046 23680 15068
rect 23714 15046 23780 15068
rect 23407 15012 23468 15046
rect 23514 15034 23558 15046
rect 23614 15034 23648 15046
rect 23714 15034 23738 15046
rect 23502 15012 23558 15034
rect 23592 15012 23648 15034
rect 23682 15012 23738 15034
rect 23772 15034 23780 15046
rect 23814 15046 23880 15068
rect 23814 15034 23828 15046
rect 23772 15012 23828 15034
rect 23862 15034 23880 15046
rect 23914 15046 23980 15068
rect 24014 15046 24101 15068
rect 23914 15034 23918 15046
rect 23862 15012 23918 15034
rect 23952 15034 23980 15046
rect 23952 15012 24008 15034
rect 24042 15012 24101 15046
rect 23407 14968 24101 15012
rect 23407 14956 23480 14968
rect 23514 14956 23580 14968
rect 23614 14956 23680 14968
rect 23714 14956 23780 14968
rect 23407 14922 23468 14956
rect 23514 14934 23558 14956
rect 23614 14934 23648 14956
rect 23714 14934 23738 14956
rect 23502 14922 23558 14934
rect 23592 14922 23648 14934
rect 23682 14922 23738 14934
rect 23772 14934 23780 14956
rect 23814 14956 23880 14968
rect 23814 14934 23828 14956
rect 23772 14922 23828 14934
rect 23862 14934 23880 14956
rect 23914 14956 23980 14968
rect 24014 14956 24101 14968
rect 23914 14934 23918 14956
rect 23862 14922 23918 14934
rect 23952 14934 23980 14956
rect 23952 14922 24008 14934
rect 24042 14922 24101 14956
rect 23407 14861 24101 14922
rect 24163 15144 24235 15148
rect 24163 15110 24182 15144
rect 24216 15110 24235 15144
rect 24163 15054 24235 15110
rect 24163 15020 24182 15054
rect 24216 15020 24235 15054
rect 24163 14964 24235 15020
rect 24163 14930 24182 14964
rect 24216 14930 24235 14964
rect 24163 14874 24235 14930
rect 23273 14799 23345 14859
rect 24163 14840 24182 14874
rect 24216 14840 24235 14874
rect 24163 14799 24235 14840
rect 23273 14780 24235 14799
rect 23273 14746 23370 14780
rect 23404 14746 23460 14780
rect 23494 14746 23550 14780
rect 23584 14746 23640 14780
rect 23674 14746 23730 14780
rect 23764 14746 23820 14780
rect 23854 14746 23910 14780
rect 23944 14746 24000 14780
rect 24034 14746 24090 14780
rect 24124 14746 24235 14780
rect 23273 14727 24235 14746
rect 24299 15130 24331 15148
rect 24365 15148 24559 15164
rect 24593 15148 24627 15182
rect 24661 15148 24695 15182
rect 24729 15148 24763 15182
rect 24797 15148 24831 15182
rect 24865 15148 24899 15182
rect 24933 15148 24967 15182
rect 25001 15148 25035 15182
rect 25069 15148 25103 15182
rect 25137 15148 25171 15182
rect 25205 15148 25239 15182
rect 25273 15148 25307 15182
rect 25341 15148 25375 15182
rect 25409 15148 25443 15182
rect 25477 15148 25511 15182
rect 25545 15148 25579 15182
rect 25613 15148 25647 15182
rect 25681 15148 25715 15182
rect 25749 15148 25783 15182
rect 25817 15148 25851 15182
rect 25885 15148 25919 15182
rect 25953 15148 25987 15182
rect 26021 15148 26055 15182
rect 26089 15148 26123 15182
rect 26157 15148 26191 15182
rect 26225 15148 26259 15182
rect 26293 15148 26327 15182
rect 26361 15148 26395 15182
rect 26429 15148 26463 15182
rect 26497 15148 26531 15182
rect 26565 15148 26599 15182
rect 26633 15148 26667 15182
rect 26701 15148 26735 15182
rect 26769 15148 26803 15182
rect 26837 15148 26871 15182
rect 26905 15148 26939 15182
rect 26973 15148 27007 15182
rect 27041 15148 27075 15182
rect 27109 15148 27143 15182
rect 27177 15148 27211 15182
rect 27245 15148 27279 15182
rect 27313 15148 27347 15182
rect 27381 15148 27415 15182
rect 27449 15148 27483 15182
rect 27517 15148 27551 15182
rect 27585 15173 28834 15182
rect 28868 15173 28964 15207
rect 27585 15149 28964 15173
rect 27585 15148 27684 15149
rect 24365 15130 24398 15148
rect 24299 15074 24398 15130
rect 24299 15040 24331 15074
rect 24365 15040 24398 15074
rect 24299 14984 24398 15040
rect 24299 14950 24331 14984
rect 24365 14950 24398 14984
rect 24299 14894 24398 14950
rect 24299 14860 24331 14894
rect 24365 14860 24398 14894
rect 24299 14804 24398 14860
rect 24299 14770 24331 14804
rect 24365 14770 24398 14804
rect 23110 14680 23144 14714
rect 23178 14680 23209 14714
rect 23110 14663 23209 14680
rect 24299 14714 24398 14770
rect 24299 14680 24331 14714
rect 24365 14680 24398 14714
rect 24299 14663 24398 14680
rect 23110 14630 24398 14663
rect 23110 14596 23240 14630
rect 23274 14596 23330 14630
rect 23364 14596 23420 14630
rect 23454 14596 23510 14630
rect 23544 14596 23600 14630
rect 23634 14596 23690 14630
rect 23724 14596 23780 14630
rect 23814 14596 23870 14630
rect 23904 14596 23960 14630
rect 23994 14596 24050 14630
rect 24084 14596 24140 14630
rect 24174 14596 24230 14630
rect 24264 14596 24398 14630
rect 23110 14564 24398 14596
rect 28834 15139 28964 15149
rect 28868 15105 28964 15139
rect 28834 15071 28964 15105
rect 28868 15037 28964 15071
rect 28834 15003 28964 15037
rect 28868 14969 28964 15003
rect 28834 14935 28964 14969
rect 28868 14901 28964 14935
rect 28834 14867 28964 14901
rect 28868 14833 28964 14867
rect 28834 14830 28964 14833
rect 29034 14830 29040 15262
rect 29670 15241 29766 15262
rect 37706 15378 37839 15412
rect 37706 15344 37749 15378
rect 37783 15344 37839 15378
rect 37706 15310 37839 15344
rect 37706 15276 37749 15310
rect 37783 15276 37839 15310
rect 29800 15241 29806 15262
rect 29670 15207 29806 15241
rect 29670 15173 29766 15207
rect 29800 15173 29806 15207
rect 29670 15139 29806 15173
rect 29670 15105 29766 15139
rect 29800 15105 29806 15139
rect 29670 15071 29806 15105
rect 29670 15037 29766 15071
rect 29800 15037 29806 15071
rect 29670 15003 29806 15037
rect 29670 14969 29766 15003
rect 29800 14969 29806 15003
rect 29670 14935 29806 14969
rect 29670 14901 29766 14935
rect 29800 14901 29806 14935
rect 29670 14867 29806 14901
rect 29670 14833 29766 14867
rect 29800 14833 29806 14867
rect 29670 14830 29806 14833
rect 37706 15242 37839 15276
rect 37706 15208 37749 15242
rect 37783 15208 37839 15242
rect 37706 15174 37839 15208
rect 37706 15140 37749 15174
rect 37783 15140 37839 15174
rect 37706 15106 37839 15140
rect 37706 15072 37749 15106
rect 37783 15072 37839 15106
rect 37706 15038 37839 15072
rect 37706 15004 37749 15038
rect 37783 15004 37839 15038
rect 37706 14970 37839 15004
rect 37706 14936 37749 14970
rect 37783 14936 37839 14970
rect 37706 14902 37839 14936
rect 37706 14868 37749 14902
rect 37783 14868 37839 14902
rect 37706 14834 37839 14868
rect 28834 14799 28868 14830
rect 28834 14731 28868 14765
rect 28834 14663 28868 14697
rect 28834 14595 28868 14629
rect 28834 14527 28868 14561
rect 28834 14459 28868 14493
rect 28834 14391 28868 14425
rect 28834 14323 28868 14357
rect 28834 14255 28868 14289
rect 28834 14190 28868 14221
rect 29766 14799 29800 14830
rect 29766 14731 29800 14765
rect 29766 14663 29800 14697
rect 29766 14595 29800 14629
rect 29766 14527 29800 14561
rect 29766 14459 29800 14493
rect 29766 14391 29800 14425
rect 29766 14323 29800 14357
rect 29766 14255 29800 14289
rect 29766 14192 29800 14221
rect 37706 14800 37749 14834
rect 37783 14800 37839 14834
rect 37706 14766 37839 14800
rect 37706 14732 37749 14766
rect 37783 14732 37839 14766
rect 37706 14698 37839 14732
rect 37706 14664 37749 14698
rect 37783 14664 37839 14698
rect 37706 14630 37839 14664
rect 37706 14596 37749 14630
rect 37783 14596 37839 14630
rect 37706 14562 37839 14596
rect 37706 14528 37749 14562
rect 37783 14528 37839 14562
rect 37706 14494 37839 14528
rect 37706 14460 37749 14494
rect 37783 14460 37839 14494
rect 37706 14426 37839 14460
rect 37706 14392 37749 14426
rect 37783 14392 37839 14426
rect 37706 14358 37839 14392
rect 37706 14324 37749 14358
rect 37783 14324 37839 14358
rect 37706 14290 37839 14324
rect 37706 14256 37749 14290
rect 37783 14256 37839 14290
rect 37706 14222 37839 14256
rect 29604 14190 29804 14192
rect 28834 14187 28964 14190
rect 28868 14153 28964 14187
rect 28834 14119 28964 14153
rect 28868 14085 28964 14119
rect 28834 14051 28964 14085
rect 28868 14017 28964 14051
rect 28834 13983 28964 14017
rect 28868 13949 28964 13983
rect 21632 13862 21666 13896
rect 21632 13794 21666 13828
rect 21632 13726 21666 13760
rect 21632 13658 21666 13692
rect 21632 13590 21666 13624
rect 21632 13522 21666 13556
rect 21632 13454 21666 13488
rect 21852 13490 26012 13922
rect 28834 13915 28964 13949
rect 28868 13881 28964 13915
rect 28834 13847 28964 13881
rect 28868 13813 28964 13847
rect 28834 13779 28964 13813
rect 28868 13758 28964 13779
rect 29034 13758 29040 14190
rect 29670 14187 29804 14190
rect 29670 14153 29766 14187
rect 29800 14153 29804 14187
rect 29670 14119 29804 14153
rect 29670 14085 29766 14119
rect 29800 14085 29804 14119
rect 29670 14051 29804 14085
rect 29670 14017 29766 14051
rect 29800 14017 29804 14051
rect 29670 13983 29804 14017
rect 29670 13949 29766 13983
rect 29800 13949 29804 13983
rect 29670 13915 29804 13949
rect 29670 13881 29766 13915
rect 29800 13881 29804 13915
rect 29670 13847 29804 13881
rect 29670 13813 29766 13847
rect 29800 13813 29804 13847
rect 29670 13779 29804 13813
rect 29670 13760 29766 13779
rect 28834 13662 28868 13745
rect 29800 13760 29804 13779
rect 37706 14188 37749 14222
rect 37783 14188 37839 14222
rect 37706 14154 37839 14188
rect 37706 14120 37749 14154
rect 37783 14120 37839 14154
rect 37706 14086 37839 14120
rect 37706 14052 37749 14086
rect 37783 14052 37839 14086
rect 37706 14018 37839 14052
rect 37706 13984 37749 14018
rect 37783 13984 37839 14018
rect 37706 13950 37839 13984
rect 37706 13916 37749 13950
rect 37783 13916 37839 13950
rect 37706 13882 37839 13916
rect 37706 13848 37749 13882
rect 37783 13848 37839 13882
rect 37706 13814 37839 13848
rect 37706 13780 37749 13814
rect 37783 13780 37839 13814
rect 29766 13662 29800 13745
rect 37706 13746 37839 13780
rect 37706 13712 37749 13746
rect 37783 13712 37839 13746
rect 37706 13678 37839 13712
rect 28834 13628 28960 13662
rect 28994 13628 29028 13662
rect 29062 13628 29096 13662
rect 29130 13628 29164 13662
rect 29198 13628 29232 13662
rect 29266 13628 29300 13662
rect 29334 13628 29368 13662
rect 29402 13628 29436 13662
rect 29470 13628 29504 13662
rect 29538 13628 29572 13662
rect 29606 13628 29640 13662
rect 29674 13628 29806 13662
rect 21852 13456 23114 13490
rect 23148 13456 23182 13490
rect 23216 13456 23250 13490
rect 23284 13456 23318 13490
rect 23352 13456 23386 13490
rect 23420 13456 23454 13490
rect 23488 13456 23522 13490
rect 23556 13456 23590 13490
rect 23624 13456 23658 13490
rect 23692 13456 23726 13490
rect 23760 13456 23794 13490
rect 23828 13456 23862 13490
rect 23896 13456 23930 13490
rect 23964 13456 23998 13490
rect 24032 13456 24066 13490
rect 24100 13456 24134 13490
rect 24168 13456 24202 13490
rect 24236 13456 24270 13490
rect 24304 13484 26012 13490
rect 24304 13456 24674 13484
rect 21852 13450 24674 13456
rect 24708 13450 24742 13484
rect 24776 13450 24810 13484
rect 24844 13450 24878 13484
rect 24912 13450 24946 13484
rect 24980 13450 25014 13484
rect 25048 13450 25082 13484
rect 25116 13450 25150 13484
rect 25184 13450 25218 13484
rect 25252 13450 25286 13484
rect 25320 13450 25354 13484
rect 25388 13450 25422 13484
rect 25456 13450 25490 13484
rect 25524 13450 25558 13484
rect 25592 13450 25626 13484
rect 25660 13450 25694 13484
rect 25728 13450 25762 13484
rect 25796 13450 25830 13484
rect 25864 13450 26012 13484
rect 21852 13422 26012 13450
rect 26398 13440 26524 13474
rect 26558 13440 26592 13474
rect 26626 13440 26660 13474
rect 26694 13440 26728 13474
rect 26762 13440 26796 13474
rect 26830 13440 26864 13474
rect 26898 13440 26932 13474
rect 26966 13440 27000 13474
rect 27034 13440 27068 13474
rect 27102 13440 27136 13474
rect 27170 13440 27204 13474
rect 27238 13440 27364 13474
rect 28840 13458 29806 13628
rect 37706 13644 37749 13678
rect 37783 13644 37839 13678
rect 37706 13610 37839 13644
rect 37706 13576 37749 13610
rect 37783 13576 37839 13610
rect 38133 15554 38167 15589
rect 38133 15486 38167 15504
rect 38133 15418 38167 15432
rect 38133 15350 38167 15360
rect 38133 15282 38167 15288
rect 38133 15214 38167 15216
rect 38133 15178 38167 15180
rect 38133 15106 38167 15112
rect 38133 15034 38167 15044
rect 38133 14962 38167 14976
rect 38133 14890 38167 14908
rect 38133 14818 38167 14840
rect 38133 14746 38167 14772
rect 38133 14674 38167 14704
rect 38133 14602 38167 14636
rect 38133 14534 38167 14568
rect 38133 14466 38167 14496
rect 38133 14398 38167 14424
rect 38133 14330 38167 14352
rect 38133 14262 38167 14280
rect 38133 14194 38167 14208
rect 38133 14126 38167 14136
rect 38133 14058 38167 14064
rect 38133 13990 38167 13992
rect 38133 13954 38167 13956
rect 38133 13882 38167 13888
rect 38133 13810 38167 13820
rect 38133 13738 38167 13752
rect 38133 13666 38167 13684
rect 38391 15554 38425 15589
rect 38391 15486 38425 15504
rect 38391 15418 38425 15432
rect 38391 15350 38425 15360
rect 38391 15282 38425 15288
rect 38391 15214 38425 15216
rect 38391 15178 38425 15180
rect 38391 15106 38425 15112
rect 38391 15034 38425 15044
rect 38391 14962 38425 14976
rect 38391 14890 38425 14908
rect 38391 14818 38425 14840
rect 38391 14746 38425 14772
rect 38391 14674 38425 14704
rect 38391 14602 38425 14636
rect 38391 14534 38425 14568
rect 38391 14466 38425 14496
rect 38391 14398 38425 14424
rect 38391 14330 38425 14352
rect 38391 14262 38425 14280
rect 38391 14194 38425 14208
rect 38391 14126 38425 14136
rect 38391 14058 38425 14064
rect 38391 13990 38425 13992
rect 38391 13954 38425 13956
rect 38391 13882 38425 13888
rect 38391 13810 38425 13820
rect 38391 13738 38425 13752
rect 38391 13666 38425 13684
rect 38133 13581 38167 13616
rect 38385 13616 38391 13621
rect 38649 15554 38683 15589
rect 38649 15486 38683 15504
rect 38649 15418 38683 15432
rect 38649 15350 38683 15360
rect 38649 15282 38683 15288
rect 38649 15214 38683 15216
rect 38649 15178 38683 15180
rect 38649 15106 38683 15112
rect 38649 15034 38683 15044
rect 38649 14962 38683 14976
rect 38649 14890 38683 14908
rect 38649 14818 38683 14840
rect 38649 14746 38683 14772
rect 38649 14674 38683 14704
rect 38649 14602 38683 14636
rect 38649 14534 38683 14568
rect 38649 14466 38683 14496
rect 38649 14398 38683 14424
rect 38649 14330 38683 14352
rect 38649 14262 38683 14280
rect 38649 14194 38683 14208
rect 38649 14126 38683 14136
rect 38649 14058 38683 14064
rect 38649 13990 38683 13992
rect 38649 13954 38683 13956
rect 38649 13882 38683 13888
rect 38649 13810 38683 13820
rect 38649 13738 38683 13752
rect 38649 13666 38683 13684
rect 38425 13616 38429 13621
rect 37706 13542 37839 13576
rect 37706 13508 37749 13542
rect 37783 13508 37839 13542
rect 37706 13474 37839 13508
rect 38385 13513 38429 13616
rect 38649 13581 38683 13616
rect 38903 15554 38947 15662
rect 38903 15504 38907 15554
rect 38941 15504 38947 15554
rect 38903 15486 38947 15504
rect 38903 15432 38907 15486
rect 38941 15432 38947 15486
rect 38903 15418 38947 15432
rect 38903 15360 38907 15418
rect 38941 15360 38947 15418
rect 38903 15350 38947 15360
rect 38903 15288 38907 15350
rect 38941 15288 38947 15350
rect 38903 15282 38947 15288
rect 38903 15216 38907 15282
rect 38941 15216 38947 15282
rect 38903 15214 38947 15216
rect 38903 15180 38907 15214
rect 38941 15180 38947 15214
rect 38903 15178 38947 15180
rect 38903 15112 38907 15178
rect 38941 15112 38947 15178
rect 38903 15106 38947 15112
rect 38903 15044 38907 15106
rect 38941 15044 38947 15106
rect 38903 15034 38947 15044
rect 38903 14976 38907 15034
rect 38941 14976 38947 15034
rect 38903 14962 38947 14976
rect 38903 14908 38907 14962
rect 38941 14908 38947 14962
rect 38903 14890 38947 14908
rect 38903 14840 38907 14890
rect 38941 14840 38947 14890
rect 38903 14818 38947 14840
rect 38903 14772 38907 14818
rect 38941 14772 38947 14818
rect 38903 14746 38947 14772
rect 38903 14704 38907 14746
rect 38941 14704 38947 14746
rect 38903 14674 38947 14704
rect 38903 14636 38907 14674
rect 38941 14636 38947 14674
rect 38903 14602 38947 14636
rect 38903 14568 38907 14602
rect 38941 14568 38947 14602
rect 38903 14534 38947 14568
rect 38903 14496 38907 14534
rect 38941 14496 38947 14534
rect 38903 14466 38947 14496
rect 38903 14424 38907 14466
rect 38941 14424 38947 14466
rect 38903 14398 38947 14424
rect 38903 14352 38907 14398
rect 38941 14352 38947 14398
rect 38903 14330 38947 14352
rect 38903 14280 38907 14330
rect 38941 14280 38947 14330
rect 38903 14262 38947 14280
rect 38903 14208 38907 14262
rect 38941 14208 38947 14262
rect 38903 14194 38947 14208
rect 38903 14136 38907 14194
rect 38941 14136 38947 14194
rect 38903 14126 38947 14136
rect 38903 14064 38907 14126
rect 38941 14064 38947 14126
rect 38903 14058 38947 14064
rect 38903 13992 38907 14058
rect 38941 13992 38947 14058
rect 38903 13990 38947 13992
rect 38903 13956 38907 13990
rect 38941 13956 38947 13990
rect 38903 13954 38947 13956
rect 38903 13888 38907 13954
rect 38941 13888 38947 13954
rect 38903 13882 38947 13888
rect 38903 13820 38907 13882
rect 38941 13820 38947 13882
rect 38903 13810 38947 13820
rect 38903 13752 38907 13810
rect 38941 13752 38947 13810
rect 38903 13738 38947 13752
rect 38903 13684 38907 13738
rect 38941 13684 38947 13738
rect 38903 13666 38947 13684
rect 38903 13616 38907 13666
rect 38941 13616 38947 13666
rect 38903 13533 38947 13616
rect 39165 15554 39199 15589
rect 39165 15486 39199 15504
rect 39165 15418 39199 15432
rect 39165 15350 39199 15360
rect 39165 15282 39199 15288
rect 39165 15214 39199 15216
rect 39165 15178 39199 15180
rect 39165 15106 39199 15112
rect 39165 15034 39199 15044
rect 39165 14962 39199 14976
rect 39165 14890 39199 14908
rect 39165 14818 39199 14840
rect 39165 14746 39199 14772
rect 39165 14674 39199 14704
rect 39165 14602 39199 14636
rect 39165 14534 39199 14568
rect 39165 14466 39199 14496
rect 39165 14398 39199 14424
rect 39165 14330 39199 14352
rect 39165 14262 39199 14280
rect 39165 14194 39199 14208
rect 39165 14126 39199 14136
rect 39165 14058 39199 14064
rect 39165 13990 39199 13992
rect 39165 13954 39199 13956
rect 39165 13882 39199 13888
rect 39165 13810 39199 13820
rect 39165 13738 39199 13752
rect 39165 13666 39199 13684
rect 39165 13581 39199 13616
rect 39419 15554 39463 15662
rect 39497 15673 39564 15707
rect 39598 15694 39896 15707
rect 40126 15704 40366 15714
rect 39598 15673 39814 15694
rect 39497 15660 39814 15673
rect 39848 15660 39896 15694
rect 39497 15624 39896 15660
rect 39932 15685 40491 15704
rect 39932 15660 40156 15685
rect 39419 15504 39423 15554
rect 39457 15504 39463 15554
rect 39419 15486 39463 15504
rect 39419 15432 39423 15486
rect 39457 15432 39463 15486
rect 39419 15418 39463 15432
rect 39419 15360 39423 15418
rect 39457 15360 39463 15418
rect 39419 15350 39463 15360
rect 39419 15288 39423 15350
rect 39457 15288 39463 15350
rect 39419 15282 39463 15288
rect 39419 15216 39423 15282
rect 39457 15216 39463 15282
rect 39419 15214 39463 15216
rect 39419 15180 39423 15214
rect 39457 15180 39463 15214
rect 39419 15178 39463 15180
rect 39419 15112 39423 15178
rect 39457 15112 39463 15178
rect 39419 15106 39463 15112
rect 39419 15044 39423 15106
rect 39457 15044 39463 15106
rect 39419 15034 39463 15044
rect 39419 14976 39423 15034
rect 39457 14976 39463 15034
rect 39419 14962 39463 14976
rect 39419 14908 39423 14962
rect 39457 14908 39463 14962
rect 39419 14890 39463 14908
rect 39419 14840 39423 14890
rect 39457 14840 39463 14890
rect 39419 14818 39463 14840
rect 39419 14772 39423 14818
rect 39457 14772 39463 14818
rect 39419 14746 39463 14772
rect 39419 14704 39423 14746
rect 39457 14704 39463 14746
rect 39419 14674 39463 14704
rect 39419 14636 39423 14674
rect 39457 14636 39463 14674
rect 39419 14602 39463 14636
rect 39419 14568 39423 14602
rect 39457 14568 39463 14602
rect 39419 14534 39463 14568
rect 39419 14496 39423 14534
rect 39457 14496 39463 14534
rect 39419 14466 39463 14496
rect 39419 14424 39423 14466
rect 39457 14424 39463 14466
rect 39419 14398 39463 14424
rect 39419 14352 39423 14398
rect 39457 14352 39463 14398
rect 39419 14330 39463 14352
rect 39419 14280 39423 14330
rect 39457 14280 39463 14330
rect 39419 14262 39463 14280
rect 39419 14208 39423 14262
rect 39457 14208 39463 14262
rect 39419 14194 39463 14208
rect 39419 14136 39423 14194
rect 39457 14136 39463 14194
rect 39419 14126 39463 14136
rect 39419 14064 39423 14126
rect 39457 14064 39463 14126
rect 39419 14058 39463 14064
rect 39419 13992 39423 14058
rect 39457 13992 39463 14058
rect 39419 13990 39463 13992
rect 39419 13956 39423 13990
rect 39457 13956 39463 13990
rect 39419 13954 39463 13956
rect 39419 13888 39423 13954
rect 39457 13888 39463 13954
rect 39419 13882 39463 13888
rect 39419 13820 39423 13882
rect 39457 13820 39463 13882
rect 39419 13810 39463 13820
rect 39419 13752 39423 13810
rect 39457 13752 39463 13810
rect 39419 13738 39463 13752
rect 39419 13684 39423 13738
rect 39457 13684 39463 13738
rect 39419 13666 39463 13684
rect 39419 13616 39423 13666
rect 39457 13616 39463 13666
rect 38718 13513 38947 13533
rect 38385 13508 38947 13513
rect 21632 13386 21666 13420
rect 21632 13318 21666 13352
rect 21632 13250 21666 13284
rect 21632 13182 21666 13216
rect 21632 13114 21666 13148
rect 21632 13046 21666 13080
rect 21632 12978 21666 13012
rect 21632 12910 21666 12944
rect 21632 12842 21666 12876
rect 21632 12774 21666 12808
rect 21632 12706 21666 12740
rect 21632 12638 21666 12672
rect 21632 12570 21666 12604
rect 21632 12502 21666 12536
rect 21632 12434 21666 12468
rect 21632 12366 21666 12400
rect 21632 12298 21666 12332
rect 21632 12230 21666 12264
rect 21632 12162 21666 12196
rect 21632 12094 21666 12128
rect 21632 12026 21666 12060
rect 21632 11958 21666 11992
rect 21632 11890 21666 11924
rect 21632 11822 21666 11856
rect 21632 11754 21666 11788
rect 21632 11686 21666 11720
rect 21632 11618 21666 11652
rect 21632 11550 21666 11584
rect 21632 11482 21666 11516
rect 21632 11414 21666 11448
rect 21632 11346 21666 11380
rect 21632 11278 21666 11312
rect 21632 11210 21666 11244
rect 21632 11142 21666 11176
rect 21632 11074 21666 11108
rect 21632 11006 21666 11040
rect 21632 10938 21666 10972
rect 21632 10870 21666 10904
rect 21632 10802 21666 10836
rect 21632 10734 21666 10768
rect 21632 10666 21666 10700
rect 21632 10598 21666 10632
rect 21632 10530 21666 10564
rect 21632 10462 21666 10496
rect 21632 10394 21666 10428
rect 21632 10326 21666 10360
rect 21632 10258 21666 10292
rect 21632 10190 21666 10224
rect 21632 10122 21666 10156
rect 21632 10054 21666 10088
rect 21632 9986 21666 10020
rect 21632 9918 21666 9952
rect 21632 9850 21666 9884
rect 21632 9782 21666 9816
rect 21632 9714 21666 9748
rect 21632 9646 21666 9680
rect 21632 9578 21666 9612
rect 21632 9510 21666 9544
rect 21632 9442 21666 9476
rect 21632 9374 21666 9408
rect 21632 9306 21666 9340
rect 21632 9238 21666 9272
rect 21632 9170 21666 9204
rect 21632 9102 21666 9136
rect 21632 9034 21666 9068
rect 21632 8966 21666 9000
rect 21632 8898 21666 8932
rect 21632 8830 21666 8864
rect 21632 8762 21666 8796
rect 21632 8694 21666 8728
rect 21632 8626 21666 8660
rect 21632 8558 21666 8592
rect 21632 8490 21666 8524
rect 21632 8422 21666 8456
rect 21632 8354 21666 8388
rect 21632 8286 21666 8320
rect 21632 8218 21666 8252
rect 21632 8150 21666 8184
rect 21632 8082 21666 8116
rect 21632 8014 21666 8048
rect 21632 7946 21666 7980
rect 21632 7878 21666 7912
rect 21632 7810 21666 7844
rect 21632 7742 21666 7776
rect 21632 7674 21666 7708
rect 21632 7606 21666 7640
rect 21632 7538 21666 7572
rect 21632 7470 21666 7504
rect 21632 7402 21666 7436
rect 21632 7334 21666 7368
rect 21632 7266 21666 7300
rect 21632 7198 21666 7232
rect 21632 7130 21666 7164
rect 21632 7062 21666 7096
rect 21862 7631 22482 13422
rect 22990 13371 23024 13422
rect 23292 13356 23572 13422
rect 24394 13371 24428 13422
rect 22990 13303 23024 13337
rect 23205 13322 23224 13356
rect 23284 13322 23296 13356
rect 23352 13322 23368 13356
rect 23420 13322 23440 13356
rect 23488 13322 23512 13356
rect 23556 13322 23584 13356
rect 23624 13322 23656 13356
rect 23692 13322 23726 13356
rect 23762 13322 23794 13356
rect 23834 13322 23862 13356
rect 23906 13322 23930 13356
rect 23978 13322 23998 13356
rect 24050 13322 24066 13356
rect 24122 13322 24134 13356
rect 24194 13322 24213 13356
rect 22990 13235 23024 13269
rect 22990 13167 23024 13201
rect 22990 13099 23024 13133
rect 22990 13031 23024 13065
rect 22990 12963 23024 12997
rect 22990 12895 23024 12929
rect 22990 12827 23024 12861
rect 22990 12759 23024 12793
rect 22990 12691 23024 12725
rect 22990 12623 23024 12657
rect 22990 12555 23024 12589
rect 22990 12487 23024 12521
rect 22990 12419 23024 12453
rect 22990 12351 23024 12385
rect 22990 12283 23024 12317
rect 23128 13269 23162 13310
rect 23128 13201 23162 13225
rect 23128 13133 23162 13153
rect 23128 13065 23162 13081
rect 23128 12997 23162 13009
rect 23128 12929 23162 12937
rect 23128 12861 23162 12865
rect 23128 12755 23162 12759
rect 23128 12683 23162 12691
rect 23128 12611 23162 12623
rect 23128 12539 23162 12555
rect 23128 12467 23162 12487
rect 23128 12395 23162 12419
rect 23128 12310 23162 12351
rect 24256 13269 24290 13310
rect 24256 13201 24290 13225
rect 24256 13133 24290 13153
rect 24256 13065 24290 13081
rect 24256 12997 24290 13009
rect 24256 12929 24290 12937
rect 24256 12861 24290 12865
rect 24256 12755 24290 12759
rect 24256 12683 24290 12691
rect 24256 12611 24290 12623
rect 24256 12539 24290 12555
rect 24256 12467 24290 12487
rect 24256 12395 24290 12419
rect 24256 12310 24290 12351
rect 24394 13303 24428 13337
rect 24394 13235 24428 13269
rect 24394 13167 24428 13201
rect 24394 13099 24428 13133
rect 24394 13031 24428 13065
rect 24394 12963 24428 12997
rect 24394 12895 24428 12929
rect 24394 12827 24428 12861
rect 24394 12759 24428 12793
rect 24394 12691 24428 12725
rect 24394 12623 24428 12657
rect 24394 12555 24428 12589
rect 24394 12487 24428 12521
rect 24394 12419 24428 12453
rect 24394 12351 24428 12385
rect 23205 12264 23224 12298
rect 23284 12264 23296 12298
rect 23352 12264 23368 12298
rect 23420 12264 23440 12298
rect 23488 12264 23512 12298
rect 23556 12264 23584 12298
rect 23624 12264 23656 12298
rect 23692 12264 23726 12298
rect 23762 12264 23794 12298
rect 23834 12264 23862 12298
rect 23906 12264 23930 12298
rect 23978 12264 23998 12298
rect 24050 12264 24066 12298
rect 24122 12264 24134 12298
rect 24194 12264 24213 12298
rect 24394 12283 24428 12317
rect 22990 12164 23024 12249
rect 24394 12164 24428 12249
rect 22990 12130 23114 12164
rect 23148 12130 23182 12164
rect 23216 12130 23250 12164
rect 23284 12130 23318 12164
rect 23352 12130 23386 12164
rect 23420 12130 23454 12164
rect 23488 12130 23522 12164
rect 23556 12130 23590 12164
rect 23624 12130 23658 12164
rect 23692 12130 23726 12164
rect 23760 12130 23794 12164
rect 23828 12130 23862 12164
rect 23896 12130 23930 12164
rect 23964 12130 23998 12164
rect 24032 12130 24066 12164
rect 24100 12130 24134 12164
rect 24168 12130 24202 12164
rect 24236 12130 24270 12164
rect 24304 12130 24428 12164
rect 24550 13376 24584 13422
rect 24972 13350 25232 13422
rect 25954 13376 25988 13422
rect 24550 13308 24584 13342
rect 24765 13316 24784 13350
rect 24844 13316 24856 13350
rect 24912 13316 24928 13350
rect 24980 13316 25000 13350
rect 25048 13316 25072 13350
rect 25116 13316 25144 13350
rect 25184 13316 25216 13350
rect 25252 13316 25286 13350
rect 25322 13316 25354 13350
rect 25394 13316 25422 13350
rect 25466 13316 25490 13350
rect 25538 13316 25558 13350
rect 25610 13316 25626 13350
rect 25682 13316 25694 13350
rect 25754 13316 25773 13350
rect 24972 13312 25232 13316
rect 25954 13308 25988 13342
rect 26398 13363 26432 13440
rect 27330 13363 27364 13440
rect 26398 13322 26432 13329
rect 24550 13240 24584 13274
rect 24550 13172 24584 13206
rect 24550 13104 24584 13138
rect 24550 13036 24584 13070
rect 24550 12968 24584 13002
rect 24550 12900 24584 12934
rect 24550 12832 24584 12866
rect 24550 12764 24584 12798
rect 24550 12696 24584 12730
rect 24550 12628 24584 12662
rect 24550 12560 24584 12594
rect 24550 12492 24584 12526
rect 24550 12424 24584 12458
rect 24550 12356 24584 12390
rect 24550 12288 24584 12322
rect 24688 13263 24722 13304
rect 24688 13195 24722 13219
rect 24688 13127 24722 13147
rect 24688 13059 24722 13075
rect 24688 12991 24722 13003
rect 24688 12923 24722 12931
rect 24688 12855 24722 12859
rect 24688 12749 24722 12753
rect 24688 12677 24722 12685
rect 24688 12605 24722 12617
rect 24688 12533 24722 12549
rect 24688 12461 24722 12481
rect 24688 12389 24722 12413
rect 24688 12304 24722 12345
rect 25816 13263 25850 13304
rect 25816 13195 25850 13219
rect 25816 13127 25850 13147
rect 25816 13059 25850 13075
rect 25816 12991 25850 13003
rect 25816 12923 25850 12931
rect 25816 12855 25850 12859
rect 25816 12749 25850 12753
rect 25816 12677 25850 12685
rect 25816 12605 25850 12617
rect 25816 12533 25850 12549
rect 25816 12461 25850 12481
rect 25816 12389 25850 12413
rect 25816 12304 25850 12345
rect 25954 13240 25988 13274
rect 25954 13172 25988 13206
rect 25954 13104 25988 13138
rect 25954 13036 25988 13070
rect 25954 12968 25988 13002
rect 25954 12900 25988 12934
rect 26392 13295 26528 13322
rect 26392 13261 26398 13295
rect 26432 13261 26528 13295
rect 26392 13227 26528 13261
rect 26392 13193 26398 13227
rect 26432 13193 26528 13227
rect 26392 13159 26528 13193
rect 26392 13125 26398 13159
rect 26432 13125 26528 13159
rect 26392 13091 26528 13125
rect 26392 13057 26398 13091
rect 26432 13057 26528 13091
rect 26392 13023 26528 13057
rect 26392 12989 26398 13023
rect 26432 12989 26528 13023
rect 26392 12955 26528 12989
rect 26392 12921 26398 12955
rect 26432 12921 26528 12955
rect 26392 12912 26528 12921
rect 27152 12912 27164 13332
rect 27234 13329 27330 13332
rect 27570 13424 27686 13458
rect 27720 13424 27754 13458
rect 27788 13424 27822 13458
rect 27856 13424 27890 13458
rect 27924 13424 27958 13458
rect 27992 13424 28026 13458
rect 28060 13424 28094 13458
rect 28128 13424 28162 13458
rect 28196 13424 28230 13458
rect 28264 13424 28298 13458
rect 28332 13424 28366 13458
rect 28400 13424 28434 13458
rect 28468 13424 28502 13458
rect 28536 13424 28570 13458
rect 28604 13424 28638 13458
rect 28672 13424 28706 13458
rect 28740 13424 28774 13458
rect 28808 13424 28842 13458
rect 28876 13424 28910 13458
rect 28944 13424 28978 13458
rect 29012 13424 29046 13458
rect 29080 13424 29114 13458
rect 29148 13424 29182 13458
rect 29216 13424 29250 13458
rect 29284 13424 29318 13458
rect 29352 13424 29386 13458
rect 29420 13424 29454 13458
rect 29488 13424 29522 13458
rect 29556 13424 29590 13458
rect 29624 13424 29658 13458
rect 29692 13424 29808 13458
rect 27570 13347 27604 13424
rect 27364 13329 27570 13332
rect 27234 13313 27570 13329
rect 29774 13347 29808 13424
rect 27604 13328 27776 13332
rect 29616 13328 29774 13330
rect 27604 13313 27700 13328
rect 27234 13295 27700 13313
rect 27234 13261 27330 13295
rect 27364 13279 27700 13295
rect 27364 13261 27570 13279
rect 27234 13245 27570 13261
rect 27604 13245 27700 13279
rect 27234 13227 27700 13245
rect 27234 13193 27330 13227
rect 27364 13211 27700 13227
rect 27364 13193 27570 13211
rect 27234 13177 27570 13193
rect 27604 13177 27700 13211
rect 27234 13159 27700 13177
rect 27234 13125 27330 13159
rect 27364 13143 27700 13159
rect 27364 13125 27570 13143
rect 27234 13109 27570 13125
rect 27604 13109 27700 13143
rect 27234 13091 27700 13109
rect 27234 13057 27330 13091
rect 27364 13075 27700 13091
rect 27364 13057 27570 13075
rect 27234 13041 27570 13057
rect 27604 13041 27700 13075
rect 27234 13023 27700 13041
rect 27234 12989 27330 13023
rect 27364 13007 27700 13023
rect 27364 12989 27570 13007
rect 27234 12973 27570 12989
rect 27604 12973 27700 13007
rect 27234 12955 27700 12973
rect 27234 12921 27330 12955
rect 27364 12939 27700 12955
rect 27364 12921 27570 12939
rect 27234 12912 27570 12921
rect 26392 12902 26592 12912
rect 27152 12905 27570 12912
rect 27604 12905 27700 12939
rect 25954 12832 25988 12866
rect 25954 12764 25988 12798
rect 25954 12696 25988 12730
rect 25954 12628 25988 12662
rect 25954 12560 25988 12594
rect 25954 12492 25988 12526
rect 25954 12424 25988 12458
rect 25954 12356 25988 12390
rect 24765 12258 24784 12292
rect 24844 12258 24856 12292
rect 24912 12258 24928 12292
rect 24980 12258 25000 12292
rect 25048 12258 25072 12292
rect 25116 12258 25144 12292
rect 25184 12258 25216 12292
rect 25252 12258 25286 12292
rect 25322 12258 25354 12292
rect 25394 12258 25422 12292
rect 25466 12258 25490 12292
rect 25538 12258 25558 12292
rect 25610 12258 25626 12292
rect 25682 12258 25694 12292
rect 25754 12258 25773 12292
rect 25954 12288 25988 12322
rect 24550 12220 24584 12254
rect 24550 12152 24584 12186
rect 24550 12084 24584 12118
rect 24550 12016 24584 12050
rect 22920 11916 23035 11950
rect 23069 11916 23103 11950
rect 23137 11916 23171 11950
rect 23205 11916 23239 11950
rect 23273 11916 23307 11950
rect 23341 11916 23375 11950
rect 23409 11916 23443 11950
rect 23477 11916 23511 11950
rect 23545 11916 23579 11950
rect 23613 11916 23647 11950
rect 23681 11916 23715 11950
rect 23749 11916 23783 11950
rect 23817 11916 23851 11950
rect 23885 11916 23919 11950
rect 23953 11916 23987 11950
rect 24021 11916 24055 11950
rect 24089 11916 24123 11950
rect 24157 11916 24191 11950
rect 24225 11916 24340 11950
rect 22920 11831 22954 11916
rect 24306 11831 24340 11916
rect 22920 11763 22954 11797
rect 23126 11782 23145 11816
rect 23205 11782 23217 11816
rect 23273 11782 23289 11816
rect 23341 11782 23361 11816
rect 23409 11782 23433 11816
rect 23477 11782 23505 11816
rect 23545 11782 23577 11816
rect 23613 11782 23647 11816
rect 23683 11782 23715 11816
rect 23755 11782 23783 11816
rect 23827 11782 23851 11816
rect 23899 11782 23919 11816
rect 23971 11782 23987 11816
rect 24043 11782 24055 11816
rect 24115 11782 24134 11816
rect 22920 11695 22954 11729
rect 22920 11627 22954 11661
rect 22920 11559 22954 11593
rect 22920 11491 22954 11525
rect 22920 11423 22954 11457
rect 22920 11355 22954 11389
rect 22920 11287 22954 11321
rect 22920 11219 22954 11253
rect 22920 11151 22954 11185
rect 22920 11083 22954 11117
rect 22920 11015 22954 11049
rect 22920 10947 22954 10981
rect 22920 10879 22954 10913
rect 22920 10811 22954 10845
rect 22920 10743 22954 10777
rect 23058 11729 23092 11770
rect 23058 11661 23092 11685
rect 23058 11593 23092 11613
rect 23058 11525 23092 11541
rect 23058 11457 23092 11469
rect 23058 11389 23092 11397
rect 23058 11321 23092 11325
rect 23058 11215 23092 11219
rect 23058 11143 23092 11151
rect 23058 11071 23092 11083
rect 23058 10999 23092 11015
rect 23058 10927 23092 10947
rect 23058 10855 23092 10879
rect 23058 10770 23092 10811
rect 24168 11729 24202 11770
rect 24168 11661 24202 11685
rect 24168 11593 24202 11613
rect 24168 11525 24202 11541
rect 24168 11457 24202 11469
rect 24168 11389 24202 11397
rect 24168 11321 24202 11325
rect 24168 11215 24202 11219
rect 24168 11143 24202 11151
rect 24168 11071 24202 11083
rect 24168 10999 24202 11015
rect 24168 10927 24202 10947
rect 24168 10855 24202 10879
rect 24168 10770 24202 10811
rect 24306 11763 24340 11797
rect 24306 11695 24340 11729
rect 24306 11627 24340 11661
rect 24306 11559 24340 11593
rect 24306 11491 24340 11525
rect 24306 11423 24340 11457
rect 24306 11355 24340 11389
rect 24306 11287 24340 11321
rect 24306 11219 24340 11253
rect 24306 11151 24340 11185
rect 24306 11083 24340 11117
rect 24306 11015 24340 11049
rect 24306 10947 24340 10981
rect 24306 10879 24340 10913
rect 24306 10811 24340 10845
rect 23126 10724 23145 10758
rect 23205 10724 23217 10758
rect 23273 10724 23289 10758
rect 23341 10724 23361 10758
rect 23409 10724 23433 10758
rect 23477 10724 23505 10758
rect 23545 10724 23577 10758
rect 23613 10724 23647 10758
rect 23683 10724 23715 10758
rect 23755 10724 23783 10758
rect 23827 10724 23851 10758
rect 23899 10724 23919 10758
rect 23971 10724 23987 10758
rect 24043 10724 24055 10758
rect 24115 10724 24134 10758
rect 24306 10743 24340 10777
rect 22920 10624 22954 10709
rect 24306 10624 24340 10709
rect 22920 10590 23035 10624
rect 23069 10590 23103 10624
rect 23137 10590 23171 10624
rect 23205 10590 23239 10624
rect 23273 10590 23307 10624
rect 23341 10590 23375 10624
rect 23409 10590 23443 10624
rect 23477 10590 23511 10624
rect 23545 10590 23579 10624
rect 23613 10590 23647 10624
rect 23681 10590 23715 10624
rect 23749 10590 23783 10624
rect 23817 10590 23851 10624
rect 23885 10590 23919 10624
rect 23953 10590 23987 10624
rect 24021 10590 24055 10624
rect 24089 10590 24123 10624
rect 24157 10590 24191 10624
rect 24225 10590 24340 10624
rect 24550 11948 24584 11982
rect 24550 11880 24584 11914
rect 24550 11812 24584 11846
rect 24550 11744 24584 11778
rect 24550 11676 24584 11710
rect 24550 11608 24584 11642
rect 24550 11540 24584 11574
rect 24550 11472 24584 11506
rect 24550 11404 24584 11438
rect 24550 11336 24584 11370
rect 24550 11268 24584 11302
rect 24688 12205 24722 12246
rect 24688 12137 24722 12161
rect 24688 12069 24722 12089
rect 24688 12001 24722 12017
rect 24688 11933 24722 11945
rect 24688 11865 24722 11873
rect 24688 11797 24722 11801
rect 24688 11691 24722 11695
rect 24688 11619 24722 11627
rect 24688 11547 24722 11559
rect 24688 11475 24722 11491
rect 24688 11403 24722 11423
rect 24688 11331 24722 11355
rect 24688 11246 24722 11287
rect 25816 12205 25850 12246
rect 25816 12137 25850 12161
rect 25816 12069 25850 12089
rect 25816 12001 25850 12017
rect 25816 11933 25850 11945
rect 25816 11865 25850 11873
rect 25816 11797 25850 11801
rect 25816 11691 25850 11695
rect 25816 11619 25850 11627
rect 25816 11547 25850 11559
rect 25816 11475 25850 11491
rect 25816 11403 25850 11423
rect 25816 11331 25850 11355
rect 25816 11246 25850 11287
rect 25954 12220 25988 12254
rect 25954 12152 25988 12186
rect 25954 12084 25988 12118
rect 25954 12016 25988 12050
rect 25954 11948 25988 11982
rect 25954 11880 25988 11914
rect 25954 11812 25988 11846
rect 25954 11744 25988 11778
rect 25954 11676 25988 11710
rect 25954 11608 25988 11642
rect 25954 11540 25988 11574
rect 25954 11472 25988 11506
rect 25954 11404 25988 11438
rect 25954 11336 25988 11370
rect 25954 11268 25988 11302
rect 24550 11200 24584 11234
rect 24765 11200 24784 11234
rect 24844 11200 24856 11234
rect 24912 11200 24928 11234
rect 24980 11200 25000 11234
rect 25048 11200 25072 11234
rect 25116 11200 25144 11234
rect 25184 11200 25216 11234
rect 25252 11200 25286 11234
rect 25322 11200 25354 11234
rect 25394 11200 25422 11234
rect 25466 11200 25490 11234
rect 25538 11200 25558 11234
rect 25610 11200 25626 11234
rect 25682 11200 25694 11234
rect 25754 11200 25773 11234
rect 25954 11200 25988 11234
rect 24550 11132 24584 11166
rect 24550 11064 24584 11098
rect 24550 10996 24584 11030
rect 24550 10928 24584 10962
rect 24550 10860 24584 10894
rect 24550 10792 24584 10826
rect 24550 10724 24584 10758
rect 24550 10656 24584 10690
rect 23672 8014 23812 10590
rect 24550 10588 24584 10622
rect 24550 10520 24584 10554
rect 24550 10452 24584 10486
rect 24550 10384 24584 10418
rect 24550 10316 24584 10350
rect 24550 10248 24584 10282
rect 24550 10180 24584 10214
rect 24688 11147 24722 11188
rect 24688 11079 24722 11103
rect 24688 11011 24722 11031
rect 24688 10943 24722 10959
rect 24688 10875 24722 10887
rect 24688 10807 24722 10815
rect 24688 10739 24722 10743
rect 24688 10633 24722 10637
rect 24688 10561 24722 10569
rect 24688 10489 24722 10501
rect 24688 10417 24722 10433
rect 24688 10345 24722 10365
rect 24688 10273 24722 10297
rect 24688 10188 24722 10229
rect 25816 11147 25850 11188
rect 25816 11079 25850 11103
rect 25816 11011 25850 11031
rect 25816 10943 25850 10959
rect 25816 10875 25850 10887
rect 25816 10807 25850 10815
rect 25816 10739 25850 10743
rect 25816 10633 25850 10637
rect 25816 10561 25850 10569
rect 25816 10489 25850 10501
rect 25816 10417 25850 10433
rect 25816 10345 25850 10365
rect 25816 10273 25850 10297
rect 25816 10188 25850 10229
rect 25954 11132 25988 11166
rect 25954 11064 25988 11098
rect 25954 10996 25988 11030
rect 25954 10928 25988 10962
rect 25954 10860 25988 10894
rect 25954 10792 25988 10826
rect 25954 10724 25988 10758
rect 25954 10656 25988 10690
rect 25954 10588 25988 10622
rect 25954 10520 25988 10554
rect 25954 10452 25988 10486
rect 25954 10384 25988 10418
rect 25954 10316 25988 10350
rect 25954 10248 25988 10282
rect 25954 10180 25988 10214
rect 24550 10112 24584 10146
rect 24765 10142 24784 10176
rect 24844 10142 24856 10176
rect 24912 10142 24928 10176
rect 24980 10142 25000 10176
rect 25048 10142 25072 10176
rect 25116 10142 25144 10176
rect 25184 10142 25216 10176
rect 25252 10142 25286 10176
rect 25322 10142 25354 10176
rect 25394 10142 25422 10176
rect 25466 10142 25490 10176
rect 25538 10142 25558 10176
rect 25610 10142 25626 10176
rect 25682 10142 25694 10176
rect 25754 10142 25773 10176
rect 24550 10044 24584 10078
rect 24550 9976 24584 10010
rect 24550 9908 24584 9942
rect 24550 9840 24584 9874
rect 24550 9772 24584 9806
rect 24550 9704 24584 9738
rect 24550 9636 24584 9670
rect 24550 9568 24584 9602
rect 24550 9500 24584 9534
rect 24550 9432 24584 9466
rect 24550 9364 24584 9398
rect 24550 9296 24584 9330
rect 24550 9228 24584 9262
rect 24550 9160 24584 9194
rect 24688 10089 24722 10130
rect 24688 10021 24722 10045
rect 24688 9953 24722 9973
rect 24688 9885 24722 9901
rect 24688 9817 24722 9829
rect 24688 9749 24722 9757
rect 24688 9681 24722 9685
rect 24688 9575 24722 9579
rect 24688 9503 24722 9511
rect 24688 9431 24722 9443
rect 24688 9359 24722 9375
rect 24688 9287 24722 9307
rect 24688 9215 24722 9239
rect 24688 9130 24722 9171
rect 25816 10089 25850 10130
rect 25816 10021 25850 10045
rect 25816 9953 25850 9973
rect 25816 9885 25850 9901
rect 25816 9817 25850 9829
rect 25816 9749 25850 9757
rect 25816 9681 25850 9685
rect 25816 9575 25850 9579
rect 25816 9503 25850 9511
rect 25816 9431 25850 9443
rect 25816 9359 25850 9375
rect 25816 9287 25850 9307
rect 25816 9215 25850 9239
rect 25816 9130 25850 9171
rect 25954 10112 25988 10146
rect 25954 10044 25988 10078
rect 25954 9976 25988 10010
rect 25954 9908 25988 9942
rect 25954 9840 25988 9874
rect 25954 9772 25988 9806
rect 25954 9704 25988 9738
rect 25954 9636 25988 9670
rect 25954 9568 25988 9602
rect 25954 9500 25988 9534
rect 25954 9432 25988 9466
rect 25954 9364 25988 9398
rect 25954 9296 25988 9330
rect 25954 9228 25988 9262
rect 25954 9160 25988 9194
rect 24550 9092 24584 9126
rect 24765 9084 24784 9118
rect 24844 9084 24856 9118
rect 24912 9084 24928 9118
rect 24980 9084 25000 9118
rect 25048 9084 25072 9118
rect 25116 9084 25144 9118
rect 25184 9084 25216 9118
rect 25252 9084 25286 9118
rect 25322 9084 25354 9118
rect 25394 9084 25422 9118
rect 25466 9084 25490 9118
rect 25538 9084 25558 9118
rect 25610 9084 25626 9118
rect 25682 9084 25694 9118
rect 25754 9084 25773 9118
rect 25954 9092 25988 9126
rect 24550 8984 24584 9058
rect 25954 8984 25988 9058
rect 24550 8950 24674 8984
rect 24708 8950 24742 8984
rect 24776 8950 24810 8984
rect 24844 8950 24878 8984
rect 24912 8950 24946 8984
rect 24980 8950 25014 8984
rect 25048 8950 25082 8984
rect 25116 8950 25150 8984
rect 25184 8950 25218 8984
rect 25252 8950 25286 8984
rect 25320 8950 25354 8984
rect 25388 8950 25422 8984
rect 25456 8950 25490 8984
rect 25524 8950 25558 8984
rect 25592 8950 25626 8984
rect 25660 8950 25694 8984
rect 25728 8950 25762 8984
rect 25796 8950 25830 8984
rect 25864 8950 25988 8984
rect 26398 12887 26432 12902
rect 27152 12900 27700 12905
rect 26398 12819 26432 12853
rect 26398 12751 26432 12785
rect 26398 12683 26432 12717
rect 26398 12615 26432 12649
rect 26398 12547 26432 12581
rect 26398 12479 26432 12513
rect 26398 12411 26432 12445
rect 26398 12343 26432 12377
rect 26398 12275 26432 12309
rect 26398 12207 26432 12241
rect 26398 12139 26432 12173
rect 26398 12071 26432 12105
rect 26398 12003 26432 12037
rect 26398 11935 26432 11969
rect 26398 11867 26432 11901
rect 26398 11799 26432 11833
rect 26398 11731 26432 11765
rect 26398 11663 26432 11697
rect 26398 11595 26432 11629
rect 26398 11527 26432 11561
rect 26398 11459 26432 11493
rect 26398 11391 26432 11425
rect 26398 11323 26432 11357
rect 26398 11255 26432 11289
rect 26398 11187 26432 11221
rect 26398 11119 26432 11153
rect 26398 11051 26432 11085
rect 26398 10983 26432 11017
rect 26398 10915 26432 10949
rect 26398 10847 26432 10881
rect 26398 10779 26432 10813
rect 26398 10711 26432 10745
rect 26398 10643 26432 10677
rect 26398 10575 26432 10609
rect 26398 10507 26432 10541
rect 26398 10439 26432 10473
rect 26398 10371 26432 10405
rect 26398 10303 26432 10337
rect 26398 10235 26432 10269
rect 26398 10167 26432 10201
rect 26398 10099 26432 10133
rect 26398 10031 26432 10065
rect 26398 9963 26432 9997
rect 26398 9895 26432 9929
rect 26398 9827 26432 9861
rect 26398 9759 26432 9793
rect 26398 9691 26432 9725
rect 26398 9623 26432 9657
rect 26398 9555 26432 9589
rect 26398 9487 26432 9521
rect 26398 9419 26432 9453
rect 26398 9351 26432 9385
rect 26398 9283 26432 9317
rect 26398 9215 26432 9249
rect 26398 9147 26432 9181
rect 26398 9079 26432 9113
rect 26398 9011 26432 9045
rect 26398 8943 26432 8977
rect 26398 8875 26432 8909
rect 26398 8807 26432 8841
rect 26398 8739 26432 8773
rect 26398 8671 26432 8705
rect 26398 8603 26432 8637
rect 26398 8535 26432 8569
rect 26398 8467 26432 8501
rect 26398 8399 26432 8433
rect 26398 8331 26432 8365
rect 26398 8263 26432 8297
rect 26398 8195 26432 8229
rect 26398 8127 26432 8161
rect 26398 8059 26432 8093
rect 21862 7093 21898 7631
rect 22436 7093 22482 7631
rect 21862 7062 22482 7093
rect 23400 7980 23515 8014
rect 23549 7980 23583 8014
rect 23617 7980 23651 8014
rect 23685 7980 23719 8014
rect 23753 7980 23787 8014
rect 23821 7980 23855 8014
rect 23889 7980 23923 8014
rect 23957 7980 23991 8014
rect 24025 7980 24059 8014
rect 24093 7980 24127 8014
rect 24161 7980 24195 8014
rect 24229 7980 24263 8014
rect 24297 7980 24331 8014
rect 24365 7980 24399 8014
rect 24433 7980 24467 8014
rect 24501 7980 24535 8014
rect 24569 7980 24603 8014
rect 24637 7980 24671 8014
rect 24705 7980 24820 8014
rect 23400 7906 23434 7980
rect 23672 7962 23812 7980
rect 24786 7906 24820 7980
rect 23400 7838 23434 7872
rect 23606 7846 23625 7880
rect 23685 7846 23697 7880
rect 23753 7846 23769 7880
rect 23821 7846 23841 7880
rect 23889 7846 23913 7880
rect 23957 7846 23985 7880
rect 24025 7846 24057 7880
rect 24093 7846 24127 7880
rect 24163 7846 24195 7880
rect 24235 7846 24263 7880
rect 24307 7846 24331 7880
rect 24379 7846 24399 7880
rect 24451 7846 24467 7880
rect 24523 7846 24535 7880
rect 24595 7846 24614 7880
rect 24786 7838 24820 7872
rect 23400 7770 23434 7804
rect 23400 7702 23434 7736
rect 23400 7634 23434 7668
rect 23400 7566 23434 7600
rect 23400 7498 23434 7532
rect 23400 7430 23434 7464
rect 23400 7362 23434 7396
rect 23400 7294 23434 7328
rect 23400 7226 23434 7260
rect 23400 7158 23434 7192
rect 23400 7090 23434 7124
rect 21632 6994 21666 7028
rect 21632 6926 21666 6960
rect 21632 6858 21666 6892
rect 21632 6790 21666 6824
rect 21632 6722 21666 6756
rect 21632 6654 21666 6688
rect 21632 6586 21666 6620
rect 21632 6518 21666 6552
rect 21632 6450 21666 6484
rect 21632 6382 21666 6416
rect 21632 6314 21666 6348
rect 21632 6246 21666 6280
rect 21632 6178 21666 6212
rect 21632 6110 21666 6144
rect 21632 6042 21666 6076
rect 21632 5974 21666 6008
rect 21632 5906 21666 5940
rect 21632 5838 21666 5872
rect 21632 5770 21666 5804
rect 21632 5702 21666 5736
rect 21632 5634 21666 5668
rect 21632 5566 21666 5600
rect 21632 5498 21666 5532
rect 21632 5430 21666 5464
rect 21632 5362 21666 5396
rect 21632 5294 21666 5328
rect 21632 5226 21666 5260
rect 20382 5158 20590 5160
rect 20416 5152 20590 5158
rect 21632 5158 21666 5192
rect 21464 5152 21632 5154
rect 20416 5124 20512 5152
rect 20382 5090 20512 5124
rect 20416 5056 20512 5090
rect 20382 5022 20512 5056
rect 20416 4988 20512 5022
rect 20382 4954 20512 4988
rect 20416 4920 20512 4954
rect 20382 4886 20512 4920
rect 20416 4852 20512 4886
rect 20382 4818 20512 4852
rect 20416 4784 20512 4818
rect 20382 4750 20512 4784
rect 20416 4724 20512 4750
rect 20582 4724 20590 5152
rect 20828 4720 20830 5152
rect 20900 4720 21148 5152
rect 21464 4720 21466 5152
rect 21536 5124 21632 5152
rect 23400 7022 23434 7056
rect 23400 6954 23434 6988
rect 23400 6886 23434 6920
rect 23400 6818 23434 6852
rect 23538 7793 23572 7834
rect 23538 7725 23572 7749
rect 23538 7657 23572 7677
rect 23538 7589 23572 7605
rect 23538 7521 23572 7533
rect 23538 7453 23572 7461
rect 23538 7385 23572 7389
rect 23538 7279 23572 7283
rect 23538 7207 23572 7215
rect 23538 7135 23572 7147
rect 23538 7063 23572 7079
rect 23538 6991 23572 7011
rect 23538 6919 23572 6943
rect 23538 6834 23572 6875
rect 24648 7793 24682 7834
rect 24648 7725 24682 7749
rect 24648 7657 24682 7677
rect 24648 7589 24682 7605
rect 24648 7521 24682 7533
rect 24648 7453 24682 7461
rect 24648 7385 24682 7389
rect 24648 7279 24682 7283
rect 24648 7207 24682 7215
rect 24648 7135 24682 7147
rect 24648 7063 24682 7079
rect 24648 6991 24682 7011
rect 24648 6919 24682 6943
rect 24648 6834 24682 6875
rect 24786 7770 24820 7804
rect 24786 7702 24820 7736
rect 24786 7634 24820 7668
rect 24786 7566 24820 7600
rect 24786 7498 24820 7532
rect 24786 7430 24820 7464
rect 24786 7362 24820 7396
rect 24786 7294 24820 7328
rect 24786 7226 24820 7260
rect 24786 7158 24820 7192
rect 24786 7090 24820 7124
rect 24786 7022 24820 7056
rect 24786 6954 24820 6988
rect 24786 6886 24820 6920
rect 23606 6788 23625 6822
rect 23685 6788 23697 6822
rect 23753 6788 23769 6822
rect 23821 6788 23841 6822
rect 23889 6788 23913 6822
rect 23957 6788 23985 6822
rect 24025 6788 24057 6822
rect 24093 6788 24127 6822
rect 24163 6788 24195 6822
rect 24235 6788 24263 6822
rect 24307 6788 24331 6822
rect 24379 6788 24399 6822
rect 24451 6788 24467 6822
rect 24523 6788 24535 6822
rect 24595 6788 24614 6822
rect 24786 6818 24820 6852
rect 23400 6750 23434 6784
rect 23400 6682 23434 6716
rect 23400 6614 23434 6648
rect 23400 6546 23434 6580
rect 23400 6478 23434 6512
rect 23400 6410 23434 6444
rect 23400 6342 23434 6376
rect 23400 6274 23434 6308
rect 23400 6206 23434 6240
rect 23400 6138 23434 6172
rect 23400 6070 23434 6104
rect 23400 6002 23434 6036
rect 23400 5934 23434 5968
rect 23400 5866 23434 5900
rect 23400 5798 23434 5832
rect 23538 6735 23572 6776
rect 23538 6667 23572 6691
rect 23538 6599 23572 6619
rect 23538 6531 23572 6547
rect 23538 6463 23572 6475
rect 23538 6395 23572 6403
rect 23538 6327 23572 6331
rect 23538 6221 23572 6225
rect 23538 6149 23572 6157
rect 23538 6077 23572 6089
rect 23538 6005 23572 6021
rect 23538 5933 23572 5953
rect 23538 5861 23572 5885
rect 23538 5776 23572 5817
rect 24648 6735 24682 6776
rect 24648 6667 24682 6691
rect 24648 6599 24682 6619
rect 24648 6531 24682 6547
rect 24648 6463 24682 6475
rect 24648 6395 24682 6403
rect 24648 6327 24682 6331
rect 24648 6221 24682 6225
rect 24648 6149 24682 6157
rect 24648 6077 24682 6089
rect 24648 6005 24682 6021
rect 24648 5933 24682 5953
rect 24648 5861 24682 5885
rect 24648 5776 24682 5817
rect 24786 6750 24820 6784
rect 24786 6682 24820 6716
rect 24786 6614 24820 6648
rect 24786 6546 24820 6580
rect 24786 6478 24820 6512
rect 24786 6410 24820 6444
rect 24786 6342 24820 6376
rect 24786 6274 24820 6308
rect 24786 6206 24820 6240
rect 24786 6138 24820 6172
rect 24786 6070 24820 6104
rect 24786 6002 24820 6036
rect 24786 5934 24820 5968
rect 24786 5866 24820 5900
rect 24786 5798 24820 5832
rect 23400 5730 23434 5764
rect 23606 5730 23625 5764
rect 23685 5730 23697 5764
rect 23753 5730 23769 5764
rect 23821 5730 23841 5764
rect 23889 5730 23913 5764
rect 23957 5730 23985 5764
rect 24025 5730 24057 5764
rect 24093 5730 24127 5764
rect 24163 5730 24195 5764
rect 24235 5730 24263 5764
rect 24307 5730 24331 5764
rect 24379 5730 24399 5764
rect 24451 5730 24467 5764
rect 24523 5730 24535 5764
rect 24595 5730 24614 5764
rect 24786 5730 24820 5764
rect 23400 5662 23434 5696
rect 23400 5594 23434 5628
rect 23400 5526 23434 5560
rect 23400 5458 23434 5492
rect 23400 5390 23434 5424
rect 23400 5322 23434 5356
rect 23400 5254 23434 5288
rect 23400 5186 23434 5220
rect 21666 5124 21670 5154
rect 21536 5090 21670 5124
rect 21536 5056 21632 5090
rect 21666 5056 21670 5090
rect 21536 5022 21670 5056
rect 21536 4988 21632 5022
rect 21666 4988 21670 5022
rect 21536 4954 21670 4988
rect 21536 4920 21632 4954
rect 21666 4920 21670 4954
rect 21536 4886 21670 4920
rect 21536 4852 21632 4886
rect 21666 4852 21670 4886
rect 21536 4818 21670 4852
rect 21536 4784 21632 4818
rect 21666 4784 21670 4818
rect 21536 4750 21670 4784
rect 21536 4720 21632 4750
rect 21464 4718 21632 4720
rect 20382 4624 20416 4716
rect 21666 4718 21670 4750
rect 23400 5118 23434 5152
rect 23400 5050 23434 5084
rect 23400 4982 23434 5016
rect 23400 4914 23434 4948
rect 23400 4846 23434 4880
rect 23400 4778 23434 4812
rect 21632 4624 21666 4716
rect 20382 4590 20497 4624
rect 20531 4590 20565 4624
rect 20599 4590 20633 4624
rect 20667 4590 20701 4624
rect 20735 4590 20769 4624
rect 20803 4590 20837 4624
rect 20871 4590 20905 4624
rect 20939 4590 20973 4624
rect 21007 4590 21041 4624
rect 21075 4590 21109 4624
rect 21143 4590 21177 4624
rect 21211 4590 21245 4624
rect 21279 4590 21313 4624
rect 21347 4590 21381 4624
rect 21415 4590 21449 4624
rect 21483 4590 21517 4624
rect 21551 4618 21666 4624
rect 23400 4710 23434 4744
rect 23538 5677 23572 5718
rect 23538 5609 23572 5633
rect 23538 5541 23572 5561
rect 23538 5473 23572 5489
rect 23538 5405 23572 5417
rect 23538 5337 23572 5345
rect 23538 5269 23572 5273
rect 23538 5163 23572 5167
rect 23538 5091 23572 5099
rect 23538 5019 23572 5031
rect 23538 4947 23572 4963
rect 23538 4875 23572 4895
rect 23538 4803 23572 4827
rect 23538 4718 23572 4759
rect 24648 5677 24682 5718
rect 24648 5609 24682 5633
rect 24648 5541 24682 5561
rect 24648 5473 24682 5489
rect 24648 5405 24682 5417
rect 24648 5337 24682 5345
rect 24648 5269 24682 5273
rect 24648 5163 24682 5167
rect 24648 5091 24682 5099
rect 24648 5019 24682 5031
rect 24648 4947 24682 4963
rect 24648 4875 24682 4895
rect 24648 4803 24682 4827
rect 24648 4718 24682 4759
rect 24786 5662 24820 5696
rect 24786 5594 24820 5628
rect 24786 5526 24820 5560
rect 24786 5458 24820 5492
rect 24786 5390 24820 5424
rect 24786 5322 24820 5356
rect 24786 5254 24820 5288
rect 24786 5186 24820 5220
rect 24786 5118 24820 5152
rect 24786 5050 24820 5084
rect 24786 4982 24820 5016
rect 24786 4914 24820 4948
rect 24786 4846 24820 4880
rect 24786 4778 24820 4812
rect 24786 4710 24820 4744
rect 23400 4642 23434 4676
rect 23606 4672 23625 4706
rect 23685 4672 23697 4706
rect 23753 4672 23769 4706
rect 23821 4672 23841 4706
rect 23889 4672 23913 4706
rect 23957 4672 23985 4706
rect 24025 4672 24057 4706
rect 24093 4672 24127 4706
rect 24163 4672 24195 4706
rect 24235 4672 24263 4706
rect 24307 4672 24331 4706
rect 24379 4672 24399 4706
rect 24451 4672 24467 4706
rect 24523 4672 24535 4706
rect 24595 4672 24614 4706
rect 21551 4590 21676 4618
rect 18750 4501 18784 4535
rect 18930 4476 18971 4510
rect 19015 4476 19039 4510
rect 19087 4476 19107 4510
rect 19159 4476 19175 4510
rect 19231 4476 19243 4510
rect 19303 4476 19311 4510
rect 19375 4476 19379 4510
rect 19481 4476 19485 4510
rect 19549 4476 19557 4510
rect 19617 4476 19629 4510
rect 19685 4476 19701 4510
rect 19753 4476 19773 4510
rect 19821 4476 19845 4510
rect 19889 4476 19930 4510
rect 20076 4501 20110 4535
rect 18750 4372 18784 4467
rect 20076 4372 20110 4467
rect 18750 4352 18869 4372
rect 18541 4338 18869 4352
rect 18903 4338 18937 4372
rect 18971 4338 19005 4372
rect 19039 4338 19073 4372
rect 19107 4338 19141 4372
rect 19175 4338 19209 4372
rect 19243 4338 19277 4372
rect 19311 4338 19345 4372
rect 19379 4338 19413 4372
rect 19447 4338 19481 4372
rect 19515 4338 19549 4372
rect 19583 4338 19617 4372
rect 19651 4338 19685 4372
rect 19719 4338 19753 4372
rect 19787 4338 19821 4372
rect 19855 4338 19889 4372
rect 19923 4338 19957 4372
rect 19991 4352 20110 4372
rect 20384 4352 21676 4590
rect 23400 4574 23434 4608
rect 23400 4506 23434 4540
rect 23400 4438 23434 4472
rect 23400 4370 23434 4404
rect 19991 4338 21682 4352
rect 12747 4300 21682 4338
rect 23400 4302 23434 4336
rect -7120 787 -5286 4213
rect 12747 4209 22876 4300
rect 12747 3815 12824 4209
rect 22650 3815 22876 4209
rect 12747 3794 22876 3815
rect 12747 3760 21682 3794
rect 16016 3756 21682 3760
rect 16016 3736 17170 3756
rect 22376 3552 22876 3794
rect 23400 4234 23434 4268
rect 23400 4166 23434 4200
rect 23400 4098 23434 4132
rect 23400 4030 23434 4064
rect 23400 3962 23434 3996
rect 23400 3894 23434 3928
rect 23400 3826 23434 3860
rect 23400 3758 23434 3792
rect 23400 3690 23434 3724
rect 23538 4619 23572 4660
rect 23538 4551 23572 4575
rect 23538 4483 23572 4503
rect 23538 4415 23572 4431
rect 23538 4347 23572 4359
rect 23538 4279 23572 4287
rect 23538 4211 23572 4215
rect 23538 4105 23572 4109
rect 23538 4033 23572 4041
rect 23538 3961 23572 3973
rect 23538 3889 23572 3905
rect 23538 3817 23572 3837
rect 23538 3745 23572 3769
rect 23538 3660 23572 3701
rect 24648 4619 24682 4660
rect 24648 4551 24682 4575
rect 24648 4483 24682 4503
rect 24648 4415 24682 4431
rect 24648 4347 24682 4359
rect 24648 4279 24682 4287
rect 24648 4211 24682 4215
rect 24648 4105 24682 4109
rect 24648 4033 24682 4041
rect 24648 3961 24682 3973
rect 24648 3889 24682 3905
rect 24648 3817 24682 3837
rect 24648 3745 24682 3769
rect 24648 3660 24682 3701
rect 24786 4642 24820 4676
rect 24786 4574 24820 4608
rect 24786 4506 24820 4540
rect 24786 4438 24820 4472
rect 24786 4370 24820 4404
rect 24786 4302 24820 4336
rect 24786 4234 24820 4268
rect 24786 4166 24820 4200
rect 24786 4098 24820 4132
rect 24786 4030 24820 4064
rect 24786 3962 24820 3996
rect 24786 3894 24820 3928
rect 24786 3826 24820 3860
rect 24786 3758 24820 3792
rect 24786 3690 24820 3724
rect 23400 3622 23434 3656
rect 23606 3614 23625 3648
rect 23685 3614 23697 3648
rect 23753 3614 23769 3648
rect 23821 3614 23841 3648
rect 23889 3614 23913 3648
rect 23957 3614 23985 3648
rect 24025 3614 24057 3648
rect 24093 3614 24127 3648
rect 24163 3614 24195 3648
rect 24235 3614 24263 3648
rect 24307 3614 24331 3648
rect 24379 3614 24399 3648
rect 24451 3614 24467 3648
rect 24523 3614 24535 3648
rect 24595 3614 24614 3648
rect 24786 3622 24820 3656
rect 23400 3552 23434 3588
rect 24786 3552 24820 3588
rect 24900 7980 25015 8014
rect 25049 7980 25083 8014
rect 25117 7980 25151 8014
rect 25185 7980 25219 8014
rect 25253 7980 25287 8014
rect 25321 7980 25355 8014
rect 25389 7980 25423 8014
rect 25457 7980 25491 8014
rect 25525 7980 25559 8014
rect 25593 7980 25627 8014
rect 25661 7980 25695 8014
rect 25729 7980 25763 8014
rect 25797 7980 25831 8014
rect 25865 7980 25899 8014
rect 25933 7980 25967 8014
rect 26001 7980 26035 8014
rect 26069 7980 26103 8014
rect 26137 7980 26171 8014
rect 26205 7980 26320 8014
rect 24900 7906 24934 7980
rect 26286 7906 26320 7980
rect 24900 7838 24934 7872
rect 25106 7846 25125 7880
rect 25185 7846 25197 7880
rect 25253 7846 25269 7880
rect 25321 7846 25341 7880
rect 25389 7846 25413 7880
rect 25457 7846 25485 7880
rect 25525 7846 25557 7880
rect 25593 7846 25627 7880
rect 25663 7846 25695 7880
rect 25735 7846 25763 7880
rect 25807 7846 25831 7880
rect 25879 7846 25899 7880
rect 25951 7846 25967 7880
rect 26023 7846 26035 7880
rect 26095 7846 26114 7880
rect 26286 7838 26320 7872
rect 24900 7770 24934 7804
rect 24900 7702 24934 7736
rect 24900 7634 24934 7668
rect 24900 7566 24934 7600
rect 24900 7498 24934 7532
rect 24900 7430 24934 7464
rect 24900 7362 24934 7396
rect 24900 7294 24934 7328
rect 24900 7226 24934 7260
rect 24900 7158 24934 7192
rect 24900 7090 24934 7124
rect 24900 7022 24934 7056
rect 24900 6954 24934 6988
rect 24900 6886 24934 6920
rect 24900 6818 24934 6852
rect 25038 7793 25072 7834
rect 25038 7725 25072 7749
rect 25038 7657 25072 7677
rect 25038 7589 25072 7605
rect 25038 7521 25072 7533
rect 25038 7453 25072 7461
rect 25038 7385 25072 7389
rect 25038 7279 25072 7283
rect 25038 7207 25072 7215
rect 25038 7135 25072 7147
rect 25038 7063 25072 7079
rect 25038 6991 25072 7011
rect 25038 6919 25072 6943
rect 25038 6834 25072 6875
rect 26148 7793 26182 7834
rect 26148 7725 26182 7749
rect 26148 7657 26182 7677
rect 26148 7589 26182 7605
rect 26148 7521 26182 7533
rect 26148 7453 26182 7461
rect 26148 7385 26182 7389
rect 26148 7279 26182 7283
rect 26148 7207 26182 7215
rect 26148 7135 26182 7147
rect 26148 7063 26182 7079
rect 26148 6991 26182 7011
rect 26148 6919 26182 6943
rect 26148 6834 26182 6875
rect 26286 7770 26320 7804
rect 26286 7702 26320 7736
rect 26286 7634 26320 7668
rect 26286 7566 26320 7600
rect 26286 7498 26320 7532
rect 26286 7430 26320 7464
rect 26286 7362 26320 7396
rect 26286 7294 26320 7328
rect 26286 7226 26320 7260
rect 26286 7158 26320 7192
rect 26286 7090 26320 7124
rect 26286 7022 26320 7056
rect 26286 6954 26320 6988
rect 26286 6886 26320 6920
rect 25106 6788 25125 6822
rect 25185 6788 25197 6822
rect 25253 6788 25269 6822
rect 25321 6788 25341 6822
rect 25389 6788 25413 6822
rect 25457 6788 25485 6822
rect 25525 6788 25557 6822
rect 25593 6788 25627 6822
rect 25663 6788 25695 6822
rect 25735 6788 25763 6822
rect 25807 6788 25831 6822
rect 25879 6788 25899 6822
rect 25951 6788 25967 6822
rect 26023 6788 26035 6822
rect 26095 6788 26114 6822
rect 26286 6818 26320 6852
rect 24900 6750 24934 6784
rect 24900 6682 24934 6716
rect 24900 6614 24934 6648
rect 24900 6546 24934 6580
rect 24900 6478 24934 6512
rect 24900 6410 24934 6444
rect 24900 6342 24934 6376
rect 24900 6274 24934 6308
rect 24900 6206 24934 6240
rect 24900 6138 24934 6172
rect 24900 6070 24934 6104
rect 24900 6002 24934 6036
rect 24900 5934 24934 5968
rect 24900 5866 24934 5900
rect 24900 5798 24934 5832
rect 25038 6735 25072 6776
rect 25038 6667 25072 6691
rect 25038 6599 25072 6619
rect 25038 6531 25072 6547
rect 25038 6463 25072 6475
rect 25038 6395 25072 6403
rect 25038 6327 25072 6331
rect 25038 6221 25072 6225
rect 25038 6149 25072 6157
rect 25038 6077 25072 6089
rect 25038 6005 25072 6021
rect 25038 5933 25072 5953
rect 25038 5861 25072 5885
rect 25038 5776 25072 5817
rect 26148 6735 26182 6776
rect 26148 6667 26182 6691
rect 26148 6599 26182 6619
rect 26148 6531 26182 6547
rect 26148 6463 26182 6475
rect 26148 6395 26182 6403
rect 26148 6327 26182 6331
rect 26148 6221 26182 6225
rect 26148 6149 26182 6157
rect 26148 6077 26182 6089
rect 26148 6005 26182 6021
rect 26148 5933 26182 5953
rect 26148 5861 26182 5885
rect 26148 5776 26182 5817
rect 26286 6750 26320 6784
rect 26286 6682 26320 6716
rect 26286 6614 26320 6648
rect 26286 6546 26320 6580
rect 26286 6478 26320 6512
rect 26286 6410 26320 6444
rect 26286 6342 26320 6376
rect 26286 6274 26320 6308
rect 26286 6206 26320 6240
rect 26286 6138 26320 6172
rect 26286 6070 26320 6104
rect 26286 6002 26320 6036
rect 26286 5934 26320 5968
rect 26286 5866 26320 5900
rect 26286 5798 26320 5832
rect 24900 5730 24934 5764
rect 25106 5730 25125 5764
rect 25185 5730 25197 5764
rect 25253 5730 25269 5764
rect 25321 5730 25341 5764
rect 25389 5730 25413 5764
rect 25457 5730 25485 5764
rect 25525 5730 25557 5764
rect 25593 5730 25627 5764
rect 25663 5730 25695 5764
rect 25735 5730 25763 5764
rect 25807 5730 25831 5764
rect 25879 5730 25899 5764
rect 25951 5730 25967 5764
rect 26023 5730 26035 5764
rect 26095 5730 26114 5764
rect 26286 5730 26320 5764
rect 24900 5662 24934 5696
rect 24900 5594 24934 5628
rect 24900 5526 24934 5560
rect 24900 5458 24934 5492
rect 24900 5390 24934 5424
rect 24900 5322 24934 5356
rect 24900 5254 24934 5288
rect 24900 5186 24934 5220
rect 24900 5118 24934 5152
rect 24900 5050 24934 5084
rect 24900 4982 24934 5016
rect 24900 4914 24934 4948
rect 24900 4846 24934 4880
rect 24900 4778 24934 4812
rect 24900 4710 24934 4744
rect 25038 5677 25072 5718
rect 25038 5609 25072 5633
rect 25038 5541 25072 5561
rect 25038 5473 25072 5489
rect 25038 5405 25072 5417
rect 25038 5337 25072 5345
rect 25038 5269 25072 5273
rect 25038 5163 25072 5167
rect 25038 5091 25072 5099
rect 25038 5019 25072 5031
rect 25038 4947 25072 4963
rect 25038 4875 25072 4895
rect 25038 4803 25072 4827
rect 25038 4718 25072 4759
rect 26148 5677 26182 5718
rect 26148 5609 26182 5633
rect 26148 5541 26182 5561
rect 26148 5473 26182 5489
rect 26148 5405 26182 5417
rect 26148 5337 26182 5345
rect 26148 5269 26182 5273
rect 26148 5163 26182 5167
rect 26148 5091 26182 5099
rect 26148 5019 26182 5031
rect 26148 4947 26182 4963
rect 26148 4875 26182 4895
rect 26148 4803 26182 4827
rect 26148 4718 26182 4759
rect 26286 5662 26320 5696
rect 26286 5594 26320 5628
rect 26286 5526 26320 5560
rect 26286 5458 26320 5492
rect 26286 5390 26320 5424
rect 26286 5322 26320 5356
rect 26286 5254 26320 5288
rect 26286 5186 26320 5220
rect 26286 5118 26320 5152
rect 26286 5050 26320 5084
rect 26286 4982 26320 5016
rect 26286 4914 26320 4948
rect 26286 4846 26320 4880
rect 26286 4778 26320 4812
rect 26286 4710 26320 4744
rect 24900 4642 24934 4676
rect 25106 4672 25125 4706
rect 25185 4672 25197 4706
rect 25253 4672 25269 4706
rect 25321 4672 25341 4706
rect 25389 4672 25413 4706
rect 25457 4672 25485 4706
rect 25525 4672 25557 4706
rect 25593 4672 25627 4706
rect 25663 4672 25695 4706
rect 25735 4672 25763 4706
rect 25807 4672 25831 4706
rect 25879 4672 25899 4706
rect 25951 4672 25967 4706
rect 26023 4672 26035 4706
rect 26095 4672 26114 4706
rect 24900 4574 24934 4608
rect 24900 4506 24934 4540
rect 24900 4438 24934 4472
rect 24900 4370 24934 4404
rect 24900 4302 24934 4336
rect 24900 4234 24934 4268
rect 24900 4166 24934 4200
rect 24900 4098 24934 4132
rect 24900 4030 24934 4064
rect 24900 3962 24934 3996
rect 24900 3894 24934 3928
rect 24900 3826 24934 3860
rect 24900 3758 24934 3792
rect 24900 3690 24934 3724
rect 25038 4619 25072 4660
rect 25038 4551 25072 4575
rect 25038 4483 25072 4503
rect 25038 4415 25072 4431
rect 25038 4347 25072 4359
rect 25038 4279 25072 4287
rect 25038 4211 25072 4215
rect 25038 4105 25072 4109
rect 25038 4033 25072 4041
rect 25038 3961 25072 3973
rect 25038 3889 25072 3905
rect 25038 3817 25072 3837
rect 25038 3745 25072 3769
rect 25038 3660 25072 3701
rect 26148 4619 26182 4660
rect 26148 4551 26182 4575
rect 26148 4483 26182 4503
rect 26148 4415 26182 4431
rect 26148 4347 26182 4359
rect 26148 4279 26182 4287
rect 26148 4211 26182 4215
rect 26148 4105 26182 4109
rect 26148 4033 26182 4041
rect 26148 3961 26182 3973
rect 26148 3889 26182 3905
rect 26148 3817 26182 3837
rect 26148 3745 26182 3769
rect 26148 3660 26182 3701
rect 26286 4642 26320 4676
rect 26286 4574 26320 4608
rect 26286 4506 26320 4540
rect 26286 4438 26320 4472
rect 26286 4370 26320 4404
rect 26286 4302 26320 4336
rect 26286 4234 26320 4268
rect 26286 4166 26320 4200
rect 26286 4098 26320 4132
rect 26286 4030 26320 4064
rect 26286 3962 26320 3996
rect 26286 3894 26320 3928
rect 26286 3826 26320 3860
rect 26286 3758 26320 3792
rect 26286 3690 26320 3724
rect 24900 3622 24934 3656
rect 25106 3614 25125 3648
rect 25185 3614 25197 3648
rect 25253 3614 25269 3648
rect 25321 3614 25341 3648
rect 25389 3614 25413 3648
rect 25457 3614 25485 3648
rect 25525 3614 25557 3648
rect 25593 3614 25627 3648
rect 25663 3614 25695 3648
rect 25735 3614 25763 3648
rect 25807 3614 25831 3648
rect 25879 3614 25899 3648
rect 25951 3614 25967 3648
rect 26023 3614 26035 3648
rect 26095 3614 26114 3648
rect 26286 3622 26320 3656
rect 24900 3552 24934 3588
rect 26286 3552 26320 3588
rect 26398 7991 26432 8025
rect 26398 7923 26432 7957
rect 26398 7855 26432 7889
rect 26398 7787 26432 7821
rect 26398 7719 26432 7753
rect 26398 7651 26432 7685
rect 26398 7583 26432 7617
rect 26398 7515 26432 7549
rect 26398 7447 26432 7481
rect 26398 7379 26432 7413
rect 26398 7311 26432 7345
rect 26398 7243 26432 7277
rect 26398 7175 26432 7209
rect 26398 7107 26432 7141
rect 26398 7039 26432 7073
rect 26398 6971 26432 7005
rect 26398 6903 26432 6937
rect 26398 6835 26432 6869
rect 26398 6767 26432 6801
rect 26398 6699 26432 6733
rect 26398 6631 26432 6665
rect 26398 6563 26432 6597
rect 26398 6495 26432 6529
rect 27318 12887 27612 12900
rect 27770 12900 27776 13328
rect 29678 13313 29774 13328
rect 37706 13440 37749 13474
rect 37783 13440 37839 13474
rect 37706 13406 37839 13440
rect 37706 13372 37749 13406
rect 37783 13372 37839 13406
rect 38200 13471 38346 13504
rect 38200 13437 38249 13471
rect 38283 13437 38346 13471
rect 38385 13474 38752 13508
rect 38786 13474 38824 13508
rect 38858 13474 38947 13508
rect 39419 13512 39463 13616
rect 39681 15554 39715 15589
rect 39681 15486 39715 15504
rect 39681 15418 39715 15432
rect 39681 15350 39715 15360
rect 39681 15282 39715 15288
rect 39681 15214 39715 15216
rect 39681 15178 39715 15180
rect 39681 15106 39715 15112
rect 39681 15034 39715 15044
rect 39681 14962 39715 14976
rect 39681 14890 39715 14908
rect 39681 14818 39715 14840
rect 39681 14746 39715 14772
rect 39681 14674 39715 14704
rect 39681 14602 39715 14636
rect 39681 14534 39715 14568
rect 39681 14466 39715 14496
rect 39681 14398 39715 14424
rect 39681 14330 39715 14352
rect 39681 14262 39715 14280
rect 39681 14194 39715 14208
rect 39681 14126 39715 14136
rect 39681 14058 39715 14064
rect 39681 13990 39715 13992
rect 39681 13954 39715 13956
rect 39681 13882 39715 13888
rect 39681 13810 39715 13820
rect 39681 13738 39715 13752
rect 39681 13666 39715 13684
rect 39681 13581 39715 13616
rect 39932 15554 39976 15660
rect 40126 15651 40156 15660
rect 40190 15651 40228 15685
rect 40262 15651 40300 15685
rect 40334 15660 40491 15685
rect 40334 15651 40366 15660
rect 40126 15624 40366 15651
rect 39932 15504 39939 15554
rect 39973 15504 39976 15554
rect 39932 15486 39976 15504
rect 39932 15432 39939 15486
rect 39973 15432 39976 15486
rect 39932 15418 39976 15432
rect 39932 15360 39939 15418
rect 39973 15360 39976 15418
rect 39932 15350 39976 15360
rect 39932 15288 39939 15350
rect 39973 15288 39976 15350
rect 39932 15282 39976 15288
rect 39932 15216 39939 15282
rect 39973 15216 39976 15282
rect 39932 15214 39976 15216
rect 39932 15180 39939 15214
rect 39973 15180 39976 15214
rect 39932 15178 39976 15180
rect 39932 15112 39939 15178
rect 39973 15112 39976 15178
rect 39932 15106 39976 15112
rect 39932 15044 39939 15106
rect 39973 15044 39976 15106
rect 39932 15034 39976 15044
rect 39932 14976 39939 15034
rect 39973 14976 39976 15034
rect 39932 14962 39976 14976
rect 39932 14908 39939 14962
rect 39973 14908 39976 14962
rect 39932 14890 39976 14908
rect 39932 14840 39939 14890
rect 39973 14840 39976 14890
rect 39932 14818 39976 14840
rect 39932 14772 39939 14818
rect 39973 14772 39976 14818
rect 39932 14746 39976 14772
rect 39932 14704 39939 14746
rect 39973 14704 39976 14746
rect 39932 14674 39976 14704
rect 39932 14636 39939 14674
rect 39973 14636 39976 14674
rect 39932 14602 39976 14636
rect 39932 14568 39939 14602
rect 39973 14568 39976 14602
rect 39932 14534 39976 14568
rect 39932 14496 39939 14534
rect 39973 14496 39976 14534
rect 39932 14466 39976 14496
rect 39932 14424 39939 14466
rect 39973 14424 39976 14466
rect 39932 14398 39976 14424
rect 39932 14352 39939 14398
rect 39973 14352 39976 14398
rect 39932 14330 39976 14352
rect 39932 14280 39939 14330
rect 39973 14280 39976 14330
rect 39932 14262 39976 14280
rect 39932 14208 39939 14262
rect 39973 14208 39976 14262
rect 39932 14194 39976 14208
rect 39932 14136 39939 14194
rect 39973 14136 39976 14194
rect 39932 14126 39976 14136
rect 39932 14064 39939 14126
rect 39973 14064 39976 14126
rect 39932 14058 39976 14064
rect 39932 13992 39939 14058
rect 39973 13992 39976 14058
rect 39932 13990 39976 13992
rect 39932 13956 39939 13990
rect 39973 13956 39976 13990
rect 39932 13954 39976 13956
rect 39932 13888 39939 13954
rect 39973 13888 39976 13954
rect 39932 13882 39976 13888
rect 39932 13820 39939 13882
rect 39973 13820 39976 13882
rect 39932 13810 39976 13820
rect 39932 13752 39939 13810
rect 39973 13752 39976 13810
rect 39932 13738 39976 13752
rect 39932 13684 39939 13738
rect 39973 13684 39976 13738
rect 39932 13666 39976 13684
rect 39932 13616 39939 13666
rect 39973 13616 39976 13666
rect 39932 13512 39976 13616
rect 40197 15554 40231 15589
rect 40447 15554 40491 15660
rect 40531 15698 40679 15815
rect 40531 15664 40585 15698
rect 40619 15664 40679 15698
rect 40531 15659 40679 15664
rect 41047 15950 41165 15984
rect 41047 15916 41089 15950
rect 41123 15916 41165 15950
rect 41047 15882 41165 15916
rect 41047 15848 41089 15882
rect 41123 15848 41165 15882
rect 41047 15814 41165 15848
rect 41047 15780 41089 15814
rect 41123 15780 41165 15814
rect 41047 15746 41165 15780
rect 41047 15712 41089 15746
rect 41123 15712 41165 15746
rect 41047 15678 41165 15712
rect 40531 15624 40671 15659
rect 41047 15644 41089 15678
rect 41123 15644 41165 15678
rect 41047 15610 41165 15644
rect 40447 15527 40455 15554
rect 40197 15486 40231 15504
rect 40197 15418 40231 15432
rect 40197 15350 40231 15360
rect 40197 15282 40231 15288
rect 40197 15214 40231 15216
rect 40197 15178 40231 15180
rect 40197 15106 40231 15112
rect 40197 15034 40231 15044
rect 40197 14962 40231 14976
rect 40197 14890 40231 14908
rect 40197 14818 40231 14840
rect 40197 14746 40231 14772
rect 40197 14674 40231 14704
rect 40197 14602 40231 14636
rect 40197 14534 40231 14568
rect 40197 14466 40231 14496
rect 40197 14398 40231 14424
rect 40197 14330 40231 14352
rect 40197 14262 40231 14280
rect 40197 14194 40231 14208
rect 40197 14126 40231 14136
rect 40197 14058 40231 14064
rect 40197 13990 40231 13992
rect 40197 13954 40231 13956
rect 40197 13882 40231 13888
rect 40197 13810 40231 13820
rect 40197 13738 40231 13752
rect 40197 13666 40231 13684
rect 40197 13581 40231 13616
rect 40489 15527 40491 15554
rect 40713 15554 40747 15589
rect 40455 15486 40489 15504
rect 40455 15418 40489 15432
rect 40455 15350 40489 15360
rect 40455 15282 40489 15288
rect 40455 15214 40489 15216
rect 40455 15178 40489 15180
rect 40455 15106 40489 15112
rect 40455 15034 40489 15044
rect 40455 14962 40489 14976
rect 40455 14890 40489 14908
rect 40455 14818 40489 14840
rect 40455 14746 40489 14772
rect 40455 14674 40489 14704
rect 40455 14602 40489 14636
rect 40455 14534 40489 14568
rect 40455 14466 40489 14496
rect 40455 14398 40489 14424
rect 40455 14330 40489 14352
rect 40455 14262 40489 14280
rect 40455 14194 40489 14208
rect 40455 14126 40489 14136
rect 40455 14058 40489 14064
rect 40455 13990 40489 13992
rect 40455 13954 40489 13956
rect 40455 13882 40489 13888
rect 40455 13810 40489 13820
rect 40455 13738 40489 13752
rect 40455 13666 40489 13684
rect 40455 13581 40489 13616
rect 40713 15486 40747 15504
rect 40713 15418 40747 15432
rect 40713 15350 40747 15360
rect 40713 15282 40747 15288
rect 40713 15214 40747 15216
rect 40713 15178 40747 15180
rect 40713 15106 40747 15112
rect 40713 15034 40747 15044
rect 40713 14962 40747 14976
rect 40713 14890 40747 14908
rect 40713 14818 40747 14840
rect 40713 14746 40747 14772
rect 40713 14674 40747 14704
rect 40713 14602 40747 14636
rect 40713 14534 40747 14568
rect 40713 14466 40747 14496
rect 40713 14398 40747 14424
rect 40713 14330 40747 14352
rect 40713 14262 40747 14280
rect 40713 14194 40747 14208
rect 40713 14126 40747 14136
rect 40713 14058 40747 14064
rect 40713 13990 40747 13992
rect 40713 13954 40747 13956
rect 40713 13882 40747 13888
rect 40713 13810 40747 13820
rect 40713 13738 40747 13752
rect 40713 13666 40747 13684
rect 40713 13581 40747 13616
rect 41047 15576 41089 15610
rect 41123 15576 41165 15610
rect 41047 15542 41165 15576
rect 41047 15508 41089 15542
rect 41123 15508 41165 15542
rect 41047 15474 41165 15508
rect 41047 15440 41089 15474
rect 41123 15440 41165 15474
rect 41047 15406 41165 15440
rect 41047 15372 41089 15406
rect 41123 15372 41165 15406
rect 41047 15338 41165 15372
rect 41047 15304 41089 15338
rect 41123 15304 41165 15338
rect 41047 15270 41165 15304
rect 41047 15236 41089 15270
rect 41123 15236 41165 15270
rect 41047 15202 41165 15236
rect 41047 15168 41089 15202
rect 41123 15168 41165 15202
rect 41047 15134 41165 15168
rect 41047 15100 41089 15134
rect 41123 15100 41165 15134
rect 41047 15066 41165 15100
rect 41047 15032 41089 15066
rect 41123 15032 41165 15066
rect 41047 14998 41165 15032
rect 41047 14964 41089 14998
rect 41123 14964 41165 14998
rect 41047 14930 41165 14964
rect 41047 14896 41089 14930
rect 41123 14896 41165 14930
rect 41047 14862 41165 14896
rect 41047 14828 41089 14862
rect 41123 14828 41165 14862
rect 41047 14794 41165 14828
rect 41047 14760 41089 14794
rect 41123 14760 41165 14794
rect 41047 14726 41165 14760
rect 41047 14692 41089 14726
rect 41123 14692 41165 14726
rect 41047 14658 41165 14692
rect 41047 14624 41089 14658
rect 41123 14624 41165 14658
rect 41047 14590 41165 14624
rect 41047 14556 41089 14590
rect 41123 14556 41165 14590
rect 41047 14522 41165 14556
rect 41047 14488 41089 14522
rect 41123 14488 41165 14522
rect 41047 14454 41165 14488
rect 41047 14420 41089 14454
rect 41123 14420 41165 14454
rect 41047 14386 41165 14420
rect 41047 14352 41089 14386
rect 41123 14352 41165 14386
rect 41047 14318 41165 14352
rect 41047 14284 41089 14318
rect 41123 14284 41165 14318
rect 41047 14250 41165 14284
rect 41047 14216 41089 14250
rect 41123 14216 41165 14250
rect 41047 14182 41165 14216
rect 41047 14148 41089 14182
rect 41123 14148 41165 14182
rect 41047 14114 41165 14148
rect 41047 14080 41089 14114
rect 41123 14080 41165 14114
rect 41047 14046 41165 14080
rect 41047 14012 41089 14046
rect 41123 14012 41165 14046
rect 41047 13978 41165 14012
rect 41047 13944 41089 13978
rect 41123 13944 41165 13978
rect 41047 13910 41165 13944
rect 41047 13876 41089 13910
rect 41123 13876 41165 13910
rect 41047 13842 41165 13876
rect 41047 13808 41089 13842
rect 41123 13808 41165 13842
rect 41047 13774 41165 13808
rect 41047 13740 41089 13774
rect 41123 13740 41165 13774
rect 41047 13706 41165 13740
rect 41047 13672 41089 13706
rect 41123 13672 41165 13706
rect 41047 13638 41165 13672
rect 41047 13604 41089 13638
rect 41123 13604 41165 13638
rect 38385 13469 38947 13474
rect 38984 13479 39135 13505
rect 38718 13457 38946 13469
rect 38200 13387 38346 13437
rect 38984 13445 39045 13479
rect 39079 13445 39135 13479
rect 37706 13338 37839 13372
rect 29808 13313 29812 13330
rect 29678 13279 29812 13313
rect 29678 13245 29774 13279
rect 29808 13245 29812 13279
rect 29678 13211 29812 13245
rect 29678 13177 29774 13211
rect 29808 13177 29812 13211
rect 29678 13143 29812 13177
rect 29678 13109 29774 13143
rect 29808 13109 29812 13143
rect 29678 13075 29812 13109
rect 29678 13041 29774 13075
rect 29808 13041 29812 13075
rect 29678 13007 29812 13041
rect 37706 13304 37749 13338
rect 37783 13304 37839 13338
rect 37706 13270 37839 13304
rect 37706 13236 37749 13270
rect 37783 13236 37839 13270
rect 37706 13202 37839 13236
rect 37706 13168 37749 13202
rect 37783 13168 37839 13202
rect 37706 13134 37839 13168
rect 38199 13302 38347 13387
rect 38199 13268 38253 13302
rect 38287 13268 38347 13302
rect 38199 13230 38347 13268
rect 38199 13196 38253 13230
rect 38287 13196 38347 13230
rect 38199 13150 38347 13196
rect 38984 13310 39135 13445
rect 38984 13276 39042 13310
rect 39076 13276 39135 13310
rect 38984 13238 39135 13276
rect 38984 13204 39042 13238
rect 39076 13204 39135 13238
rect 38984 13151 39135 13204
rect 39233 13474 39381 13504
rect 39233 13440 39282 13474
rect 39316 13440 39381 13474
rect 39419 13468 39976 13512
rect 41047 13570 41165 13604
rect 41047 13536 41089 13570
rect 41123 13536 41165 13570
rect 40019 13476 40164 13505
rect 41047 13502 41165 13536
rect 39233 13312 39381 13440
rect 39233 13278 39282 13312
rect 39316 13278 39381 13312
rect 39233 13240 39381 13278
rect 39233 13206 39282 13240
rect 39316 13206 39381 13240
rect 39233 13153 39381 13206
rect 40019 13442 40076 13476
rect 40110 13442 40164 13476
rect 40019 13307 40164 13442
rect 40019 13273 40061 13307
rect 40095 13273 40164 13307
rect 40019 13235 40164 13273
rect 40019 13201 40061 13235
rect 40095 13201 40164 13235
rect 40019 13153 40164 13201
rect 40271 13476 40427 13501
rect 40271 13442 40331 13476
rect 40365 13442 40427 13476
rect 40271 13320 40427 13442
rect 40271 13286 40330 13320
rect 40364 13286 40427 13320
rect 40271 13248 40427 13286
rect 40271 13214 40330 13248
rect 40364 13214 40427 13248
rect 40271 13153 40427 13214
rect 41047 13468 41089 13502
rect 41123 13468 41165 13502
rect 41047 13434 41165 13468
rect 41047 13400 41089 13434
rect 41123 13400 41165 13434
rect 41047 13366 41165 13400
rect 41047 13332 41089 13366
rect 41123 13332 41165 13366
rect 41047 13298 41165 13332
rect 41047 13264 41089 13298
rect 41123 13264 41165 13298
rect 41047 13230 41165 13264
rect 41047 13196 41089 13230
rect 41123 13196 41165 13230
rect 41047 13162 41165 13196
rect 37706 13100 37749 13134
rect 37783 13100 37839 13134
rect 37706 13028 37839 13100
rect 41047 13128 41089 13162
rect 41123 13128 41165 13162
rect 41047 13094 41165 13128
rect 41582 15751 41696 15785
rect 41730 15751 41764 15785
rect 41798 15751 41912 15785
rect 41582 15664 41616 15751
rect 41878 15664 41912 15751
rect 41582 15596 41616 15630
rect 41582 15528 41616 15562
rect 41582 15460 41616 15494
rect 41582 15392 41616 15426
rect 41582 15324 41616 15358
rect 41582 15256 41616 15290
rect 41878 15596 41912 15630
rect 41878 15528 41912 15562
rect 41878 15460 41912 15494
rect 41878 15392 41912 15426
rect 41878 15324 41912 15358
rect 41878 15256 41912 15290
rect 41582 15188 41616 15222
rect 41582 15120 41616 15154
rect 41582 15052 41616 15086
rect 41582 14984 41616 15018
rect 41582 14916 41616 14950
rect 41582 14848 41616 14882
rect 41582 14780 41616 14814
rect 41582 14712 41616 14746
rect 41582 14644 41616 14678
rect 41582 14576 41616 14610
rect 41582 14508 41616 14542
rect 41582 14440 41616 14474
rect 41582 14372 41616 14406
rect 41582 14304 41616 14338
rect 41582 14236 41616 14270
rect 41582 14168 41616 14202
rect 41582 14100 41616 14134
rect 41582 14032 41616 14066
rect 41582 13964 41616 13998
rect 41582 13896 41616 13930
rect 41582 13828 41616 13862
rect 41582 13760 41616 13794
rect 41582 13692 41616 13726
rect 41582 13624 41616 13658
rect 41878 15188 41912 15222
rect 41878 15120 41912 15154
rect 41878 15052 41912 15086
rect 41878 14984 41912 15018
rect 41878 14916 41912 14950
rect 41878 14848 41912 14882
rect 41878 14780 41912 14814
rect 41878 14712 41912 14746
rect 41878 14644 41912 14678
rect 41878 14576 41912 14610
rect 41878 14508 41912 14542
rect 41878 14440 41912 14474
rect 41878 14372 41912 14406
rect 41878 14304 41912 14338
rect 41878 14236 41912 14270
rect 41878 14168 41912 14202
rect 41878 14100 41912 14134
rect 41878 14032 41912 14066
rect 41878 13964 41912 13998
rect 41878 13896 41912 13930
rect 41878 13828 41912 13862
rect 41878 13760 41912 13794
rect 41878 13692 41912 13726
rect 41878 13624 41912 13658
rect 41582 13556 41616 13590
rect 41582 13488 41616 13522
rect 41582 13420 41616 13454
rect 41582 13352 41616 13386
rect 41582 13284 41616 13318
rect 41582 13216 41616 13250
rect 41878 13556 41912 13590
rect 41878 13488 41912 13522
rect 41878 13420 41912 13454
rect 41878 13352 41912 13386
rect 41878 13284 41912 13318
rect 41878 13216 41912 13250
rect 41582 13105 41616 13182
rect 41878 13105 41912 13182
rect 41047 13060 41089 13094
rect 41123 13060 41165 13094
rect 41510 13095 41966 13105
rect 41510 13076 41696 13095
rect 41047 13028 41165 13060
rect 41506 13061 41696 13076
rect 41730 13061 41764 13095
rect 41798 13061 41966 13095
rect 29678 12973 29774 13007
rect 29808 12973 29812 13007
rect 29678 12939 29812 12973
rect 29678 12905 29774 12939
rect 29808 12905 29812 12939
rect 37704 12986 41171 13028
rect 37704 12952 38022 12986
rect 38056 12952 38090 12986
rect 38124 12952 38158 12986
rect 38192 12952 38226 12986
rect 38260 12952 38294 12986
rect 38328 12952 38362 12986
rect 38396 12952 38430 12986
rect 38464 12952 38498 12986
rect 38532 12952 38566 12986
rect 38600 12952 38634 12986
rect 38668 12952 38702 12986
rect 38736 12952 38770 12986
rect 38804 12952 38838 12986
rect 38872 12952 38906 12986
rect 38940 12952 38974 12986
rect 39008 12952 39042 12986
rect 39076 12952 39110 12986
rect 39144 12952 39178 12986
rect 39212 12952 39246 12986
rect 39280 12952 39314 12986
rect 39348 12952 39382 12986
rect 39416 12952 39450 12986
rect 39484 12952 39518 12986
rect 39552 12952 39586 12986
rect 39620 12952 39654 12986
rect 39688 12952 39722 12986
rect 39756 12952 39790 12986
rect 39824 12952 39858 12986
rect 39892 12952 39926 12986
rect 39960 12952 39994 12986
rect 40028 12952 40062 12986
rect 40096 12952 40130 12986
rect 40164 12952 40198 12986
rect 40232 12952 40266 12986
rect 40300 12952 40334 12986
rect 40368 12952 40402 12986
rect 40436 12952 40470 12986
rect 40504 12952 40538 12986
rect 40572 12952 40606 12986
rect 40640 12952 40674 12986
rect 40708 12952 40742 12986
rect 40776 12952 40810 12986
rect 40844 12952 40878 12986
rect 40912 12952 40946 12986
rect 40980 12952 41171 12986
rect 37704 12934 41171 12952
rect 41506 12934 41966 13061
rect 37704 12913 41966 12934
rect 29678 12900 29812 12905
rect 27318 12853 27330 12887
rect 27364 12871 27612 12887
rect 27364 12853 27570 12871
rect 27318 12837 27570 12853
rect 27604 12837 27612 12871
rect 27318 12819 27612 12837
rect 27318 12785 27330 12819
rect 27364 12803 27612 12819
rect 27364 12785 27570 12803
rect 27318 12769 27570 12785
rect 27604 12769 27612 12803
rect 27318 12751 27612 12769
rect 27318 12717 27330 12751
rect 27364 12735 27612 12751
rect 27364 12717 27570 12735
rect 27318 12701 27570 12717
rect 27604 12701 27612 12735
rect 27318 12683 27612 12701
rect 27318 12649 27330 12683
rect 27364 12667 27612 12683
rect 27364 12649 27570 12667
rect 27318 12633 27570 12649
rect 27604 12633 27612 12667
rect 27318 12615 27612 12633
rect 27318 12581 27330 12615
rect 27364 12599 27612 12615
rect 27364 12581 27570 12599
rect 27318 12565 27570 12581
rect 27604 12565 27612 12599
rect 27318 12547 27612 12565
rect 27318 12513 27330 12547
rect 27364 12531 27612 12547
rect 27364 12513 27570 12531
rect 27318 12497 27570 12513
rect 27604 12497 27612 12531
rect 27318 12479 27612 12497
rect 27318 12445 27330 12479
rect 27364 12463 27612 12479
rect 27364 12445 27570 12463
rect 27318 12429 27570 12445
rect 27604 12429 27612 12463
rect 27318 12411 27612 12429
rect 27318 12377 27330 12411
rect 27364 12395 27612 12411
rect 27364 12377 27570 12395
rect 27318 12361 27570 12377
rect 27604 12361 27612 12395
rect 27318 12343 27612 12361
rect 27318 12309 27330 12343
rect 27364 12327 27612 12343
rect 27364 12309 27570 12327
rect 27318 12293 27570 12309
rect 27604 12293 27612 12327
rect 27318 12275 27612 12293
rect 27318 12241 27330 12275
rect 27364 12259 27612 12275
rect 27364 12241 27570 12259
rect 27318 12225 27570 12241
rect 27604 12225 27612 12259
rect 27318 12207 27612 12225
rect 27318 12173 27330 12207
rect 27364 12191 27612 12207
rect 27364 12173 27570 12191
rect 27318 12157 27570 12173
rect 27604 12157 27612 12191
rect 27318 12139 27612 12157
rect 27318 12105 27330 12139
rect 27364 12123 27612 12139
rect 27364 12105 27570 12123
rect 27318 12089 27570 12105
rect 27604 12089 27612 12123
rect 27318 12071 27612 12089
rect 27318 12037 27330 12071
rect 27364 12055 27612 12071
rect 27364 12037 27570 12055
rect 27318 12021 27570 12037
rect 27604 12021 27612 12055
rect 27318 12003 27612 12021
rect 27318 11969 27330 12003
rect 27364 11987 27612 12003
rect 27364 11969 27570 11987
rect 27318 11953 27570 11969
rect 27604 11953 27612 11987
rect 27318 11935 27612 11953
rect 27318 11901 27330 11935
rect 27364 11919 27612 11935
rect 27364 11901 27570 11919
rect 27318 11885 27570 11901
rect 27604 11885 27612 11919
rect 27318 11867 27612 11885
rect 27318 11833 27330 11867
rect 27364 11851 27612 11867
rect 27364 11833 27570 11851
rect 27318 11817 27570 11833
rect 27604 11817 27612 11851
rect 27318 11799 27612 11817
rect 27318 11765 27330 11799
rect 27364 11783 27612 11799
rect 27364 11765 27570 11783
rect 27318 11749 27570 11765
rect 27604 11749 27612 11783
rect 27318 11731 27612 11749
rect 27318 11697 27330 11731
rect 27364 11715 27612 11731
rect 27364 11697 27570 11715
rect 27318 11681 27570 11697
rect 27604 11681 27612 11715
rect 27318 11663 27612 11681
rect 27318 11629 27330 11663
rect 27364 11647 27612 11663
rect 27364 11629 27570 11647
rect 27318 11613 27570 11629
rect 27604 11613 27612 11647
rect 27318 11595 27612 11613
rect 27318 11561 27330 11595
rect 27364 11579 27612 11595
rect 27364 11561 27570 11579
rect 27318 11545 27570 11561
rect 27604 11545 27612 11579
rect 27318 11527 27612 11545
rect 27318 11493 27330 11527
rect 27364 11511 27612 11527
rect 27364 11493 27570 11511
rect 27318 11477 27570 11493
rect 27604 11477 27612 11511
rect 27318 11459 27612 11477
rect 27318 11425 27330 11459
rect 27364 11443 27612 11459
rect 27364 11425 27570 11443
rect 27318 11409 27570 11425
rect 27604 11409 27612 11443
rect 27318 11391 27612 11409
rect 27318 11357 27330 11391
rect 27364 11375 27612 11391
rect 27364 11357 27570 11375
rect 27318 11341 27570 11357
rect 27604 11341 27612 11375
rect 27318 11323 27612 11341
rect 27318 11289 27330 11323
rect 27364 11307 27612 11323
rect 27364 11289 27570 11307
rect 27318 11273 27570 11289
rect 27604 11273 27612 11307
rect 27318 11255 27612 11273
rect 27318 11221 27330 11255
rect 27364 11239 27612 11255
rect 27364 11221 27570 11239
rect 27318 11205 27570 11221
rect 27604 11205 27612 11239
rect 27318 11187 27612 11205
rect 27318 11153 27330 11187
rect 27364 11171 27612 11187
rect 27364 11153 27570 11171
rect 27318 11137 27570 11153
rect 27604 11137 27612 11171
rect 27318 11119 27612 11137
rect 27318 11085 27330 11119
rect 27364 11103 27612 11119
rect 27364 11085 27570 11103
rect 27318 11069 27570 11085
rect 27604 11069 27612 11103
rect 27318 11051 27612 11069
rect 27318 11017 27330 11051
rect 27364 11035 27612 11051
rect 27364 11017 27570 11035
rect 27318 11001 27570 11017
rect 27604 11001 27612 11035
rect 27318 10983 27612 11001
rect 27318 10949 27330 10983
rect 27364 10967 27612 10983
rect 27364 10949 27570 10967
rect 27318 10933 27570 10949
rect 27604 10933 27612 10967
rect 27318 10915 27612 10933
rect 27318 10881 27330 10915
rect 27364 10899 27612 10915
rect 27364 10881 27570 10899
rect 27318 10865 27570 10881
rect 27604 10865 27612 10899
rect 27318 10847 27612 10865
rect 27318 10813 27330 10847
rect 27364 10831 27612 10847
rect 27364 10813 27570 10831
rect 27318 10797 27570 10813
rect 27604 10797 27612 10831
rect 27318 10779 27612 10797
rect 27318 10745 27330 10779
rect 27364 10763 27612 10779
rect 27364 10745 27570 10763
rect 27318 10729 27570 10745
rect 27604 10729 27612 10763
rect 27318 10711 27612 10729
rect 27318 10677 27330 10711
rect 27364 10695 27612 10711
rect 27364 10677 27570 10695
rect 27318 10661 27570 10677
rect 27604 10661 27612 10695
rect 27318 10643 27612 10661
rect 27318 10609 27330 10643
rect 27364 10627 27612 10643
rect 27364 10609 27570 10627
rect 27318 10593 27570 10609
rect 27604 10593 27612 10627
rect 27318 10575 27612 10593
rect 27318 10541 27330 10575
rect 27364 10559 27612 10575
rect 27364 10541 27570 10559
rect 27318 10525 27570 10541
rect 27604 10525 27612 10559
rect 27318 10507 27612 10525
rect 27318 10473 27330 10507
rect 27364 10491 27612 10507
rect 27364 10473 27570 10491
rect 27318 10457 27570 10473
rect 27604 10457 27612 10491
rect 27318 10439 27612 10457
rect 27318 10405 27330 10439
rect 27364 10423 27612 10439
rect 27364 10405 27570 10423
rect 27318 10389 27570 10405
rect 27604 10389 27612 10423
rect 27318 10371 27612 10389
rect 27318 10337 27330 10371
rect 27364 10355 27612 10371
rect 27364 10337 27570 10355
rect 27318 10321 27570 10337
rect 27604 10321 27612 10355
rect 27318 10303 27612 10321
rect 27318 10269 27330 10303
rect 27364 10287 27612 10303
rect 27364 10269 27570 10287
rect 27318 10253 27570 10269
rect 27604 10253 27612 10287
rect 27318 10235 27612 10253
rect 27318 10201 27330 10235
rect 27364 10219 27612 10235
rect 27364 10201 27570 10219
rect 27318 10185 27570 10201
rect 27604 10185 27612 10219
rect 27318 10167 27612 10185
rect 27318 10133 27330 10167
rect 27364 10151 27612 10167
rect 27364 10133 27570 10151
rect 27318 10117 27570 10133
rect 27604 10117 27612 10151
rect 27318 10099 27612 10117
rect 27318 10065 27330 10099
rect 27364 10083 27612 10099
rect 27364 10065 27570 10083
rect 27318 10049 27570 10065
rect 27604 10049 27612 10083
rect 27318 10031 27612 10049
rect 27318 9997 27330 10031
rect 27364 10015 27612 10031
rect 27364 9997 27570 10015
rect 27318 9981 27570 9997
rect 27604 9981 27612 10015
rect 27318 9963 27612 9981
rect 27318 9929 27330 9963
rect 27364 9947 27612 9963
rect 27364 9929 27570 9947
rect 27318 9913 27570 9929
rect 27604 9913 27612 9947
rect 27318 9895 27612 9913
rect 27318 9861 27330 9895
rect 27364 9879 27612 9895
rect 27364 9861 27570 9879
rect 27318 9845 27570 9861
rect 27604 9845 27612 9879
rect 27318 9827 27612 9845
rect 27318 9793 27330 9827
rect 27364 9811 27612 9827
rect 27364 9793 27570 9811
rect 27318 9777 27570 9793
rect 27604 9777 27612 9811
rect 27318 9759 27612 9777
rect 27318 9725 27330 9759
rect 27364 9743 27612 9759
rect 27364 9725 27570 9743
rect 27318 9709 27570 9725
rect 27604 9709 27612 9743
rect 27318 9691 27612 9709
rect 27318 9657 27330 9691
rect 27364 9675 27612 9691
rect 27364 9657 27570 9675
rect 27318 9641 27570 9657
rect 27604 9641 27612 9675
rect 27318 9623 27612 9641
rect 27318 9589 27330 9623
rect 27364 9607 27612 9623
rect 27364 9589 27570 9607
rect 27318 9573 27570 9589
rect 27604 9573 27612 9607
rect 27318 9555 27612 9573
rect 27318 9521 27330 9555
rect 27364 9539 27612 9555
rect 27364 9521 27570 9539
rect 27318 9505 27570 9521
rect 27604 9505 27612 9539
rect 27318 9487 27612 9505
rect 27318 9453 27330 9487
rect 27364 9471 27612 9487
rect 27364 9453 27570 9471
rect 27318 9437 27570 9453
rect 27604 9437 27612 9471
rect 27318 9419 27612 9437
rect 27318 9385 27330 9419
rect 27364 9403 27612 9419
rect 27364 9385 27570 9403
rect 27318 9369 27570 9385
rect 27604 9369 27612 9403
rect 27318 9351 27612 9369
rect 27318 9317 27330 9351
rect 27364 9335 27612 9351
rect 27364 9317 27570 9335
rect 27318 9301 27570 9317
rect 27604 9301 27612 9335
rect 27318 9283 27612 9301
rect 27318 9249 27330 9283
rect 27364 9267 27612 9283
rect 27364 9249 27570 9267
rect 27318 9233 27570 9249
rect 27604 9233 27612 9267
rect 27318 9215 27612 9233
rect 27318 9181 27330 9215
rect 27364 9199 27612 9215
rect 27364 9181 27570 9199
rect 27318 9165 27570 9181
rect 27604 9165 27612 9199
rect 27318 9147 27612 9165
rect 27318 9113 27330 9147
rect 27364 9131 27612 9147
rect 27364 9113 27570 9131
rect 27318 9097 27570 9113
rect 27604 9097 27612 9131
rect 27318 9079 27612 9097
rect 27318 9045 27330 9079
rect 27364 9063 27612 9079
rect 27364 9045 27570 9063
rect 27318 9029 27570 9045
rect 27604 9029 27612 9063
rect 27318 9011 27612 9029
rect 27318 8977 27330 9011
rect 27364 8995 27612 9011
rect 27364 8977 27570 8995
rect 27318 8961 27570 8977
rect 27604 8961 27612 8995
rect 27318 8943 27612 8961
rect 27318 8909 27330 8943
rect 27364 8927 27612 8943
rect 27364 8909 27570 8927
rect 27318 8893 27570 8909
rect 27604 8893 27612 8927
rect 27318 8875 27612 8893
rect 27318 8841 27330 8875
rect 27364 8859 27612 8875
rect 27364 8841 27570 8859
rect 27318 8825 27570 8841
rect 27604 8825 27612 8859
rect 27318 8807 27612 8825
rect 27318 8773 27330 8807
rect 27364 8791 27612 8807
rect 27364 8773 27570 8791
rect 27318 8757 27570 8773
rect 27604 8757 27612 8791
rect 27318 8739 27612 8757
rect 27318 8705 27330 8739
rect 27364 8723 27612 8739
rect 27364 8705 27570 8723
rect 27318 8689 27570 8705
rect 27604 8689 27612 8723
rect 27318 8671 27612 8689
rect 27318 8637 27330 8671
rect 27364 8655 27612 8671
rect 27364 8637 27570 8655
rect 27318 8621 27570 8637
rect 27604 8621 27612 8655
rect 27318 8603 27612 8621
rect 27318 8569 27330 8603
rect 27364 8587 27612 8603
rect 27364 8569 27570 8587
rect 27318 8553 27570 8569
rect 27604 8553 27612 8587
rect 27318 8535 27612 8553
rect 27318 8501 27330 8535
rect 27364 8519 27612 8535
rect 27364 8501 27570 8519
rect 27318 8485 27570 8501
rect 27604 8485 27612 8519
rect 27318 8467 27612 8485
rect 27318 8433 27330 8467
rect 27364 8451 27612 8467
rect 27364 8433 27570 8451
rect 27318 8417 27570 8433
rect 27604 8417 27612 8451
rect 27318 8399 27612 8417
rect 27318 8365 27330 8399
rect 27364 8383 27612 8399
rect 27364 8365 27570 8383
rect 27318 8349 27570 8365
rect 27604 8349 27612 8383
rect 27318 8331 27612 8349
rect 27318 8297 27330 8331
rect 27364 8315 27612 8331
rect 27364 8297 27570 8315
rect 27318 8281 27570 8297
rect 27604 8281 27612 8315
rect 27318 8263 27612 8281
rect 27318 8229 27330 8263
rect 27364 8247 27612 8263
rect 27364 8229 27570 8247
rect 27318 8213 27570 8229
rect 27604 8213 27612 8247
rect 27318 8195 27612 8213
rect 27318 8161 27330 8195
rect 27364 8179 27612 8195
rect 27364 8161 27570 8179
rect 27318 8145 27570 8161
rect 27604 8145 27612 8179
rect 27318 8127 27612 8145
rect 27318 8093 27330 8127
rect 27364 8111 27612 8127
rect 27364 8093 27570 8111
rect 27318 8077 27570 8093
rect 27604 8077 27612 8111
rect 27318 8059 27612 8077
rect 27318 8025 27330 8059
rect 27364 8043 27612 8059
rect 27364 8025 27570 8043
rect 27318 8009 27570 8025
rect 27604 8009 27612 8043
rect 27318 7991 27612 8009
rect 27318 7957 27330 7991
rect 27364 7975 27612 7991
rect 27364 7957 27570 7975
rect 27318 7941 27570 7957
rect 27604 7941 27612 7975
rect 27318 7923 27612 7941
rect 27318 7889 27330 7923
rect 27364 7907 27612 7923
rect 27364 7889 27570 7907
rect 27318 7873 27570 7889
rect 27604 7873 27612 7907
rect 27318 7855 27612 7873
rect 27318 7821 27330 7855
rect 27364 7839 27612 7855
rect 27364 7821 27570 7839
rect 27318 7805 27570 7821
rect 27604 7805 27612 7839
rect 27318 7787 27612 7805
rect 27318 7753 27330 7787
rect 27364 7771 27612 7787
rect 27364 7753 27570 7771
rect 27318 7737 27570 7753
rect 27604 7737 27612 7771
rect 27318 7719 27612 7737
rect 27318 7685 27330 7719
rect 27364 7703 27612 7719
rect 27364 7685 27570 7703
rect 27318 7669 27570 7685
rect 27604 7669 27612 7703
rect 27318 7651 27612 7669
rect 27318 7617 27330 7651
rect 27364 7635 27612 7651
rect 27364 7617 27570 7635
rect 27318 7601 27570 7617
rect 27604 7601 27612 7635
rect 27318 7583 27612 7601
rect 27318 7549 27330 7583
rect 27364 7567 27612 7583
rect 27364 7549 27570 7567
rect 27318 7533 27570 7549
rect 27604 7533 27612 7567
rect 27318 7515 27612 7533
rect 27318 7481 27330 7515
rect 27364 7499 27612 7515
rect 27364 7481 27570 7499
rect 27318 7465 27570 7481
rect 27604 7465 27612 7499
rect 27318 7447 27612 7465
rect 27318 7413 27330 7447
rect 27364 7431 27612 7447
rect 27364 7413 27570 7431
rect 27318 7397 27570 7413
rect 27604 7397 27612 7431
rect 27318 7379 27612 7397
rect 27318 7345 27330 7379
rect 27364 7363 27612 7379
rect 27364 7345 27570 7363
rect 27318 7329 27570 7345
rect 27604 7329 27612 7363
rect 27318 7311 27612 7329
rect 27318 7277 27330 7311
rect 27364 7295 27612 7311
rect 27364 7277 27570 7295
rect 27318 7261 27570 7277
rect 27604 7261 27612 7295
rect 27318 7243 27612 7261
rect 27318 7209 27330 7243
rect 27364 7227 27612 7243
rect 27364 7209 27570 7227
rect 27318 7193 27570 7209
rect 27604 7193 27612 7227
rect 27318 7175 27612 7193
rect 27318 7141 27330 7175
rect 27364 7159 27612 7175
rect 27364 7141 27570 7159
rect 27318 7125 27570 7141
rect 27604 7125 27612 7159
rect 27318 7107 27612 7125
rect 27318 7073 27330 7107
rect 27364 7091 27612 7107
rect 27364 7073 27570 7091
rect 27318 7057 27570 7073
rect 27604 7057 27612 7091
rect 27318 7039 27612 7057
rect 27318 7005 27330 7039
rect 27364 7023 27612 7039
rect 27364 7005 27570 7023
rect 27318 6989 27570 7005
rect 27604 6989 27612 7023
rect 27318 6971 27612 6989
rect 27318 6937 27330 6971
rect 27364 6955 27612 6971
rect 27364 6937 27570 6955
rect 27318 6921 27570 6937
rect 27604 6921 27612 6955
rect 27318 6903 27612 6921
rect 27318 6869 27330 6903
rect 27364 6898 27612 6903
rect 29774 12871 29808 12900
rect 29774 12803 29808 12837
rect 29774 12735 29808 12769
rect 29774 12667 29808 12701
rect 29774 12599 29808 12633
rect 29774 12531 29808 12565
rect 29774 12463 29808 12497
rect 29774 12395 29808 12429
rect 29774 12327 29808 12361
rect 37686 12663 41966 12913
rect 37686 12345 41186 12663
rect 41510 12661 41966 12663
rect 29774 12259 29808 12293
rect 29774 12191 29808 12225
rect 29774 12123 29808 12157
rect 29774 12055 29808 12089
rect 29774 11987 29808 12021
rect 29774 11919 29808 11953
rect 29774 11851 29808 11885
rect 29774 11783 29808 11817
rect 29774 11715 29808 11749
rect 29774 11647 29808 11681
rect 29774 11579 29808 11613
rect 29774 11511 29808 11545
rect 29774 11443 29808 11477
rect 29774 11375 29808 11409
rect 29774 11307 29808 11341
rect 29774 11239 29808 11273
rect 29774 11171 29808 11205
rect 29774 11103 29808 11137
rect 29774 11035 29808 11069
rect 29774 10967 29808 11001
rect 29774 10899 29808 10933
rect 29774 10831 29808 10865
rect 29774 10763 29808 10797
rect 29774 10695 29808 10729
rect 29774 10627 29808 10661
rect 29774 10559 29808 10593
rect 29774 10491 29808 10525
rect 29774 10423 29808 10457
rect 29774 10355 29808 10389
rect 29774 10287 29808 10321
rect 29774 10219 29808 10253
rect 29774 10151 29808 10185
rect 29774 10083 29808 10117
rect 29774 10015 29808 10049
rect 29774 9947 29808 9981
rect 29774 9879 29808 9913
rect 29774 9811 29808 9845
rect 29774 9743 29808 9777
rect 29774 9675 29808 9709
rect 29774 9607 29808 9641
rect 29774 9539 29808 9573
rect 29774 9471 29808 9505
rect 29774 9403 29808 9437
rect 29774 9335 29808 9369
rect 29774 9267 29808 9301
rect 29774 9199 29808 9233
rect 29774 9131 29808 9165
rect 29774 9063 29808 9097
rect 36484 12315 42303 12345
rect 36484 12281 36760 12315
rect 36794 12281 36828 12315
rect 36862 12281 36896 12315
rect 36930 12281 36964 12315
rect 36998 12281 37032 12315
rect 37066 12281 37100 12315
rect 37134 12281 37168 12315
rect 37202 12281 37236 12315
rect 37270 12281 37304 12315
rect 37338 12281 37372 12315
rect 37406 12281 37440 12315
rect 37474 12281 37508 12315
rect 37542 12281 37576 12315
rect 37610 12281 37644 12315
rect 37678 12281 37712 12315
rect 37746 12281 37780 12315
rect 37814 12281 37848 12315
rect 37882 12281 37916 12315
rect 37950 12281 37984 12315
rect 38018 12281 38052 12315
rect 38086 12281 38120 12315
rect 38154 12281 38188 12315
rect 38222 12281 38256 12315
rect 38290 12281 38324 12315
rect 38358 12281 38392 12315
rect 38426 12281 38460 12315
rect 38494 12281 38528 12315
rect 38562 12281 38596 12315
rect 38630 12281 38664 12315
rect 38698 12281 38732 12315
rect 38766 12281 38800 12315
rect 38834 12281 38868 12315
rect 38902 12281 38936 12315
rect 38970 12281 39004 12315
rect 39038 12281 39072 12315
rect 39106 12281 39140 12315
rect 39174 12281 39208 12315
rect 39242 12281 39276 12315
rect 39310 12281 39344 12315
rect 39378 12281 39412 12315
rect 39446 12281 39480 12315
rect 39514 12281 39548 12315
rect 39582 12281 39616 12315
rect 39650 12281 39684 12315
rect 39718 12281 39752 12315
rect 39786 12281 39820 12315
rect 39854 12281 39888 12315
rect 39922 12281 39956 12315
rect 39990 12281 40024 12315
rect 40058 12281 40092 12315
rect 40126 12281 40160 12315
rect 40194 12281 40228 12315
rect 40262 12281 40296 12315
rect 40330 12281 40364 12315
rect 40398 12281 40432 12315
rect 40466 12281 40500 12315
rect 40534 12281 40568 12315
rect 40602 12281 40636 12315
rect 40670 12281 40704 12315
rect 40738 12281 40772 12315
rect 40806 12281 40840 12315
rect 40874 12281 40908 12315
rect 40942 12281 40976 12315
rect 41010 12281 41044 12315
rect 41078 12281 41112 12315
rect 41146 12281 41180 12315
rect 41214 12281 41248 12315
rect 41282 12281 41316 12315
rect 41350 12281 41384 12315
rect 41418 12281 41452 12315
rect 41486 12281 41520 12315
rect 41554 12281 41588 12315
rect 41622 12281 41656 12315
rect 41690 12281 41724 12315
rect 41758 12281 41792 12315
rect 41826 12281 41860 12315
rect 41894 12281 41928 12315
rect 41962 12281 41996 12315
rect 42030 12281 42303 12315
rect 36484 12251 42303 12281
rect 36484 12125 36576 12251
rect 36484 12091 36511 12125
rect 36545 12091 36576 12125
rect 36484 12057 36576 12091
rect 36484 12023 36511 12057
rect 36545 12023 36576 12057
rect 36484 11989 36576 12023
rect 36484 11955 36511 11989
rect 36545 11955 36576 11989
rect 42203 12085 42303 12251
rect 42203 12051 42237 12085
rect 42271 12051 42303 12085
rect 42203 12017 42303 12051
rect 36484 11921 36576 11955
rect 36823 11952 36870 11986
rect 36906 11952 36940 11986
rect 36976 11952 37023 11986
rect 37081 11952 37128 11986
rect 37164 11952 37198 11986
rect 37234 11952 37281 11986
rect 37339 11952 37386 11986
rect 37422 11952 37456 11986
rect 37492 11952 37539 11986
rect 37597 11952 37644 11986
rect 37680 11952 37714 11986
rect 37750 11952 37797 11986
rect 37855 11952 37902 11986
rect 37938 11952 37972 11986
rect 38008 11952 38055 11986
rect 38113 11952 38160 11986
rect 38196 11952 38230 11986
rect 38266 11952 38313 11986
rect 38371 11952 38418 11986
rect 38454 11952 38488 11986
rect 38524 11952 38571 11986
rect 38629 11952 38676 11986
rect 38712 11952 38746 11986
rect 38782 11952 38829 11986
rect 38887 11952 38934 11986
rect 38970 11952 39004 11986
rect 39040 11952 39087 11986
rect 39145 11952 39192 11986
rect 39228 11952 39262 11986
rect 39298 11952 39345 11986
rect 39403 11952 39450 11986
rect 39486 11952 39520 11986
rect 39556 11952 39603 11986
rect 39661 11952 39708 11986
rect 39744 11952 39778 11986
rect 39814 11952 39861 11986
rect 39919 11952 39966 11986
rect 40002 11952 40036 11986
rect 40072 11952 40119 11986
rect 40177 11952 40224 11986
rect 40260 11952 40294 11986
rect 40330 11952 40377 11986
rect 40435 11952 40482 11986
rect 40518 11952 40552 11986
rect 40588 11952 40635 11986
rect 40693 11952 40740 11986
rect 40776 11952 40810 11986
rect 40846 11952 40893 11986
rect 40951 11952 40998 11986
rect 41034 11952 41068 11986
rect 41104 11952 41151 11986
rect 41209 11952 41256 11986
rect 41292 11952 41326 11986
rect 41362 11952 41409 11986
rect 41467 11952 41514 11986
rect 41550 11952 41584 11986
rect 41620 11952 41667 11986
rect 41725 11952 41772 11986
rect 41808 11952 41842 11986
rect 41878 11952 41925 11986
rect 42203 11983 42237 12017
rect 42271 11983 42303 12017
rect 36484 11887 36511 11921
rect 36545 11887 36576 11921
rect 42203 11949 42303 11983
rect 36484 11853 36576 11887
rect 36484 11819 36511 11853
rect 36545 11819 36576 11853
rect 36484 11785 36576 11819
rect 36484 11751 36511 11785
rect 36545 11751 36576 11785
rect 36484 11717 36576 11751
rect 36484 11683 36511 11717
rect 36545 11683 36576 11717
rect 36484 11649 36576 11683
rect 36484 11615 36511 11649
rect 36545 11615 36576 11649
rect 36484 11581 36576 11615
rect 36484 11547 36511 11581
rect 36545 11547 36576 11581
rect 36484 11513 36576 11547
rect 36484 11479 36511 11513
rect 36545 11479 36576 11513
rect 36484 11445 36576 11479
rect 36484 11411 36511 11445
rect 36545 11411 36576 11445
rect 36484 11377 36576 11411
rect 36484 11343 36511 11377
rect 36545 11343 36576 11377
rect 36484 11309 36576 11343
rect 36484 11275 36511 11309
rect 36545 11275 36576 11309
rect 36484 11241 36576 11275
rect 36484 11207 36511 11241
rect 36545 11207 36576 11241
rect 36484 11173 36576 11207
rect 36484 11139 36511 11173
rect 36545 11139 36576 11173
rect 36484 11105 36576 11139
rect 36484 11071 36511 11105
rect 36545 11071 36576 11105
rect 36484 11037 36576 11071
rect 36484 11003 36511 11037
rect 36545 11003 36576 11037
rect 36484 10969 36576 11003
rect 36484 10935 36511 10969
rect 36545 10935 36576 10969
rect 36484 10901 36576 10935
rect 36777 11899 36811 11918
rect 36777 11827 36811 11839
rect 36777 11755 36811 11771
rect 36777 11683 36811 11703
rect 36777 11611 36811 11635
rect 36777 11539 36811 11567
rect 36777 11467 36811 11499
rect 36777 11397 36811 11431
rect 36777 11329 36811 11361
rect 36777 11261 36811 11289
rect 36777 11193 36811 11217
rect 36777 11125 36811 11145
rect 36777 11057 36811 11073
rect 36777 10989 36811 11001
rect 36777 10910 36811 10929
rect 37035 11899 37069 11918
rect 37035 11827 37069 11839
rect 37035 11755 37069 11771
rect 37035 11683 37069 11703
rect 37035 11611 37069 11635
rect 37035 11539 37069 11567
rect 37035 11467 37069 11499
rect 37035 11397 37069 11431
rect 37035 11329 37069 11361
rect 37035 11261 37069 11289
rect 37035 11193 37069 11217
rect 37035 11125 37069 11145
rect 37035 11057 37069 11073
rect 37035 10989 37069 11001
rect 37035 10910 37069 10929
rect 37293 11899 37327 11918
rect 37293 11827 37327 11839
rect 37293 11755 37327 11771
rect 37293 11683 37327 11703
rect 37293 11611 37327 11635
rect 37293 11539 37327 11567
rect 37293 11467 37327 11499
rect 37293 11397 37327 11431
rect 37293 11329 37327 11361
rect 37293 11261 37327 11289
rect 37293 11193 37327 11217
rect 37293 11125 37327 11145
rect 37293 11057 37327 11073
rect 37293 10989 37327 11001
rect 37293 10910 37327 10929
rect 37551 11899 37585 11918
rect 37551 11827 37585 11839
rect 37551 11755 37585 11771
rect 37551 11683 37585 11703
rect 37551 11611 37585 11635
rect 37551 11539 37585 11567
rect 37551 11467 37585 11499
rect 37551 11397 37585 11431
rect 37551 11329 37585 11361
rect 37551 11261 37585 11289
rect 37551 11193 37585 11217
rect 37551 11125 37585 11145
rect 37551 11057 37585 11073
rect 37551 10989 37585 11001
rect 37551 10910 37585 10929
rect 37809 11899 37843 11918
rect 37809 11827 37843 11839
rect 37809 11755 37843 11771
rect 37809 11683 37843 11703
rect 37809 11611 37843 11635
rect 37809 11539 37843 11567
rect 37809 11467 37843 11499
rect 37809 11397 37843 11431
rect 37809 11329 37843 11361
rect 37809 11261 37843 11289
rect 37809 11193 37843 11217
rect 37809 11125 37843 11145
rect 37809 11057 37843 11073
rect 37809 10989 37843 11001
rect 37809 10910 37843 10929
rect 38067 11899 38101 11918
rect 38067 11827 38101 11839
rect 38067 11755 38101 11771
rect 38067 11683 38101 11703
rect 38067 11611 38101 11635
rect 38067 11539 38101 11567
rect 38067 11467 38101 11499
rect 38067 11397 38101 11431
rect 38067 11329 38101 11361
rect 38067 11261 38101 11289
rect 38067 11193 38101 11217
rect 38067 11125 38101 11145
rect 38067 11057 38101 11073
rect 38067 10989 38101 11001
rect 38067 10910 38101 10929
rect 38325 11899 38359 11918
rect 38325 11827 38359 11839
rect 38325 11755 38359 11771
rect 38325 11683 38359 11703
rect 38325 11611 38359 11635
rect 38325 11539 38359 11567
rect 38325 11467 38359 11499
rect 38325 11397 38359 11431
rect 38325 11329 38359 11361
rect 38325 11261 38359 11289
rect 38325 11193 38359 11217
rect 38325 11125 38359 11145
rect 38325 11057 38359 11073
rect 38325 10989 38359 11001
rect 38325 10910 38359 10929
rect 38583 11899 38617 11918
rect 38583 11827 38617 11839
rect 38583 11755 38617 11771
rect 38583 11683 38617 11703
rect 38583 11611 38617 11635
rect 38583 11539 38617 11567
rect 38583 11467 38617 11499
rect 38583 11397 38617 11431
rect 38583 11329 38617 11361
rect 38583 11261 38617 11289
rect 38583 11193 38617 11217
rect 38583 11125 38617 11145
rect 38583 11057 38617 11073
rect 38583 10989 38617 11001
rect 38583 10910 38617 10929
rect 38841 11899 38875 11918
rect 38841 11827 38875 11839
rect 38841 11755 38875 11771
rect 38841 11683 38875 11703
rect 38841 11611 38875 11635
rect 38841 11539 38875 11567
rect 38841 11467 38875 11499
rect 38841 11397 38875 11431
rect 38841 11329 38875 11361
rect 38841 11261 38875 11289
rect 38841 11193 38875 11217
rect 38841 11125 38875 11145
rect 38841 11057 38875 11073
rect 38841 10989 38875 11001
rect 38841 10910 38875 10929
rect 39099 11899 39133 11918
rect 39099 11827 39133 11839
rect 39099 11755 39133 11771
rect 39099 11683 39133 11703
rect 39099 11611 39133 11635
rect 39099 11539 39133 11567
rect 39099 11467 39133 11499
rect 39099 11397 39133 11431
rect 39099 11329 39133 11361
rect 39099 11261 39133 11289
rect 39099 11193 39133 11217
rect 39099 11125 39133 11145
rect 39099 11057 39133 11073
rect 39099 10989 39133 11001
rect 39099 10910 39133 10929
rect 39357 11899 39391 11918
rect 39357 11827 39391 11839
rect 39357 11755 39391 11771
rect 39357 11683 39391 11703
rect 39357 11611 39391 11635
rect 39357 11539 39391 11567
rect 39357 11467 39391 11499
rect 39357 11397 39391 11431
rect 39357 11329 39391 11361
rect 39357 11261 39391 11289
rect 39357 11193 39391 11217
rect 39357 11125 39391 11145
rect 39357 11057 39391 11073
rect 39357 10989 39391 11001
rect 39357 10910 39391 10929
rect 39615 11899 39649 11918
rect 39615 11827 39649 11839
rect 39615 11755 39649 11771
rect 39615 11683 39649 11703
rect 39615 11611 39649 11635
rect 39615 11539 39649 11567
rect 39615 11467 39649 11499
rect 39615 11397 39649 11431
rect 39615 11329 39649 11361
rect 39615 11261 39649 11289
rect 39615 11193 39649 11217
rect 39615 11125 39649 11145
rect 39615 11057 39649 11073
rect 39615 10989 39649 11001
rect 39615 10910 39649 10929
rect 39873 11899 39907 11918
rect 39873 11827 39907 11839
rect 39873 11755 39907 11771
rect 39873 11683 39907 11703
rect 39873 11611 39907 11635
rect 39873 11539 39907 11567
rect 39873 11467 39907 11499
rect 39873 11397 39907 11431
rect 39873 11329 39907 11361
rect 39873 11261 39907 11289
rect 39873 11193 39907 11217
rect 39873 11125 39907 11145
rect 39873 11057 39907 11073
rect 39873 10989 39907 11001
rect 39873 10910 39907 10929
rect 40131 11899 40165 11918
rect 40131 11827 40165 11839
rect 40131 11755 40165 11771
rect 40131 11683 40165 11703
rect 40131 11611 40165 11635
rect 40131 11539 40165 11567
rect 40131 11467 40165 11499
rect 40131 11397 40165 11431
rect 40131 11329 40165 11361
rect 40131 11261 40165 11289
rect 40131 11193 40165 11217
rect 40131 11125 40165 11145
rect 40131 11057 40165 11073
rect 40131 10989 40165 11001
rect 40131 10910 40165 10929
rect 40389 11899 40423 11918
rect 40389 11827 40423 11839
rect 40389 11755 40423 11771
rect 40389 11683 40423 11703
rect 40389 11611 40423 11635
rect 40389 11539 40423 11567
rect 40389 11467 40423 11499
rect 40389 11397 40423 11431
rect 40389 11329 40423 11361
rect 40389 11261 40423 11289
rect 40389 11193 40423 11217
rect 40389 11125 40423 11145
rect 40389 11057 40423 11073
rect 40389 10989 40423 11001
rect 40389 10910 40423 10929
rect 40647 11899 40681 11918
rect 40647 11827 40681 11839
rect 40647 11755 40681 11771
rect 40647 11683 40681 11703
rect 40647 11611 40681 11635
rect 40647 11539 40681 11567
rect 40647 11467 40681 11499
rect 40647 11397 40681 11431
rect 40647 11329 40681 11361
rect 40647 11261 40681 11289
rect 40647 11193 40681 11217
rect 40647 11125 40681 11145
rect 40647 11057 40681 11073
rect 40647 10989 40681 11001
rect 40647 10910 40681 10929
rect 40905 11899 40939 11918
rect 40905 11827 40939 11839
rect 40905 11755 40939 11771
rect 40905 11683 40939 11703
rect 40905 11611 40939 11635
rect 40905 11539 40939 11567
rect 40905 11467 40939 11499
rect 40905 11397 40939 11431
rect 40905 11329 40939 11361
rect 40905 11261 40939 11289
rect 40905 11193 40939 11217
rect 40905 11125 40939 11145
rect 40905 11057 40939 11073
rect 40905 10989 40939 11001
rect 40905 10910 40939 10929
rect 41163 11899 41197 11918
rect 41163 11827 41197 11839
rect 41163 11755 41197 11771
rect 41163 11683 41197 11703
rect 41163 11611 41197 11635
rect 41163 11539 41197 11567
rect 41163 11467 41197 11499
rect 41163 11397 41197 11431
rect 41163 11329 41197 11361
rect 41163 11261 41197 11289
rect 41163 11193 41197 11217
rect 41163 11125 41197 11145
rect 41163 11057 41197 11073
rect 41163 10989 41197 11001
rect 41163 10910 41197 10929
rect 41421 11899 41455 11918
rect 41421 11827 41455 11839
rect 41421 11755 41455 11771
rect 41421 11683 41455 11703
rect 41421 11611 41455 11635
rect 41421 11539 41455 11567
rect 41421 11467 41455 11499
rect 41421 11397 41455 11431
rect 41421 11329 41455 11361
rect 41421 11261 41455 11289
rect 41421 11193 41455 11217
rect 41421 11125 41455 11145
rect 41421 11057 41455 11073
rect 41421 10989 41455 11001
rect 41421 10910 41455 10929
rect 41679 11899 41713 11918
rect 41679 11827 41713 11839
rect 41679 11755 41713 11771
rect 41679 11683 41713 11703
rect 41679 11611 41713 11635
rect 41679 11539 41713 11567
rect 41679 11467 41713 11499
rect 41679 11397 41713 11431
rect 41679 11329 41713 11361
rect 41679 11261 41713 11289
rect 41679 11193 41713 11217
rect 41679 11125 41713 11145
rect 41679 11057 41713 11073
rect 41679 10989 41713 11001
rect 41679 10910 41713 10929
rect 41937 11899 41971 11918
rect 41937 11827 41971 11839
rect 41937 11755 41971 11771
rect 41937 11683 41971 11703
rect 41937 11611 41971 11635
rect 41937 11539 41971 11567
rect 41937 11467 41971 11499
rect 41937 11397 41971 11431
rect 41937 11329 41971 11361
rect 41937 11261 41971 11289
rect 41937 11193 41971 11217
rect 41937 11125 41971 11145
rect 41937 11057 41971 11073
rect 41937 10989 41971 11001
rect 41937 10910 41971 10929
rect 42203 11915 42237 11949
rect 42271 11915 42303 11949
rect 42203 11881 42303 11915
rect 42203 11847 42237 11881
rect 42271 11847 42303 11881
rect 42203 11813 42303 11847
rect 42203 11779 42237 11813
rect 42271 11779 42303 11813
rect 42203 11745 42303 11779
rect 42203 11711 42237 11745
rect 42271 11711 42303 11745
rect 42203 11677 42303 11711
rect 42203 11643 42237 11677
rect 42271 11643 42303 11677
rect 42203 11609 42303 11643
rect 42203 11575 42237 11609
rect 42271 11575 42303 11609
rect 42203 11541 42303 11575
rect 42203 11507 42237 11541
rect 42271 11507 42303 11541
rect 42203 11473 42303 11507
rect 42203 11439 42237 11473
rect 42271 11439 42303 11473
rect 42203 11405 42303 11439
rect 42203 11371 42237 11405
rect 42271 11371 42303 11405
rect 42203 11337 42303 11371
rect 42203 11303 42237 11337
rect 42271 11303 42303 11337
rect 42203 11269 42303 11303
rect 42203 11235 42237 11269
rect 42271 11235 42303 11269
rect 42203 11201 42303 11235
rect 42203 11167 42237 11201
rect 42271 11167 42303 11201
rect 42203 11133 42303 11167
rect 42203 11099 42237 11133
rect 42271 11099 42303 11133
rect 42203 11065 42303 11099
rect 42203 11031 42237 11065
rect 42271 11031 42303 11065
rect 42203 10997 42303 11031
rect 42203 10963 42237 10997
rect 42271 10963 42303 10997
rect 42203 10929 42303 10963
rect 36484 10867 36511 10901
rect 36545 10867 36576 10901
rect 42203 10895 42237 10929
rect 42271 10895 42303 10929
rect 36484 10833 36576 10867
rect 36823 10842 36870 10876
rect 36906 10842 36940 10876
rect 36976 10842 37023 10876
rect 37081 10842 37128 10876
rect 37164 10842 37198 10876
rect 37234 10842 37281 10876
rect 37339 10842 37386 10876
rect 37422 10842 37456 10876
rect 37492 10842 37539 10876
rect 37597 10842 37644 10876
rect 37680 10842 37714 10876
rect 37750 10842 37797 10876
rect 37855 10842 37902 10876
rect 37938 10842 37972 10876
rect 38008 10842 38055 10876
rect 38113 10842 38160 10876
rect 38196 10842 38230 10876
rect 38266 10842 38313 10876
rect 38371 10842 38418 10876
rect 38454 10842 38488 10876
rect 38524 10842 38571 10876
rect 38629 10842 38676 10876
rect 38712 10842 38746 10876
rect 38782 10842 38829 10876
rect 38887 10842 38934 10876
rect 38970 10842 39004 10876
rect 39040 10842 39087 10876
rect 39145 10842 39192 10876
rect 39228 10842 39262 10876
rect 39298 10842 39345 10876
rect 39403 10842 39450 10876
rect 39486 10842 39520 10876
rect 39556 10842 39603 10876
rect 39661 10842 39708 10876
rect 39744 10842 39778 10876
rect 39814 10842 39861 10876
rect 39919 10842 39966 10876
rect 40002 10842 40036 10876
rect 40072 10842 40119 10876
rect 40177 10842 40224 10876
rect 40260 10842 40294 10876
rect 40330 10842 40377 10876
rect 40435 10842 40482 10876
rect 40518 10842 40552 10876
rect 40588 10842 40635 10876
rect 40693 10842 40740 10876
rect 40776 10842 40810 10876
rect 40846 10842 40893 10876
rect 40951 10842 40998 10876
rect 41034 10842 41068 10876
rect 41104 10842 41151 10876
rect 41209 10842 41256 10876
rect 41292 10842 41326 10876
rect 41362 10842 41409 10876
rect 41467 10842 41514 10876
rect 41550 10842 41584 10876
rect 41620 10842 41667 10876
rect 41725 10842 41772 10876
rect 41808 10842 41842 10876
rect 41878 10842 41925 10876
rect 42203 10861 42303 10895
rect 36484 10799 36511 10833
rect 36545 10799 36576 10833
rect 36484 10765 36576 10799
rect 36484 10731 36511 10765
rect 36545 10731 36576 10765
rect 36484 10697 36576 10731
rect 36484 10663 36511 10697
rect 36545 10663 36576 10697
rect 36484 10629 36576 10663
rect 36484 10595 36511 10629
rect 36545 10595 36576 10629
rect 42203 10827 42237 10861
rect 42271 10827 42303 10861
rect 42203 10793 42303 10827
rect 42203 10759 42237 10793
rect 42271 10759 42303 10793
rect 42203 10725 42303 10759
rect 42203 10691 42237 10725
rect 42271 10691 42303 10725
rect 42203 10657 42303 10691
rect 42203 10623 42237 10657
rect 42271 10623 42303 10657
rect 36484 10561 36576 10595
rect 37858 10587 37905 10621
rect 37941 10587 37975 10621
rect 38011 10587 38058 10621
rect 38324 10587 38371 10621
rect 38407 10587 38441 10621
rect 38477 10587 38524 10621
rect 38582 10587 38629 10621
rect 38665 10587 38699 10621
rect 38735 10587 38782 10621
rect 38840 10587 38887 10621
rect 38923 10587 38957 10621
rect 38993 10587 39040 10621
rect 39098 10587 39145 10621
rect 39181 10587 39215 10621
rect 39251 10587 39298 10621
rect 39356 10587 39403 10621
rect 39439 10587 39473 10621
rect 39509 10587 39556 10621
rect 39614 10587 39661 10621
rect 39697 10587 39731 10621
rect 39767 10587 39814 10621
rect 39872 10587 39919 10621
rect 39955 10587 39989 10621
rect 40025 10587 40072 10621
rect 40130 10587 40177 10621
rect 40213 10587 40247 10621
rect 40283 10587 40330 10621
rect 40388 10587 40435 10621
rect 40471 10587 40505 10621
rect 40541 10587 40588 10621
rect 40646 10587 40693 10621
rect 40729 10587 40763 10621
rect 40799 10587 40846 10621
rect 42203 10589 42303 10623
rect 36484 10527 36511 10561
rect 36545 10527 36576 10561
rect 42203 10555 42237 10589
rect 42271 10555 42303 10589
rect 36484 10493 36576 10527
rect 36484 10459 36511 10493
rect 36545 10459 36576 10493
rect 36484 10425 36576 10459
rect 36484 10391 36511 10425
rect 36545 10391 36576 10425
rect 36484 10357 36576 10391
rect 36484 10323 36511 10357
rect 36545 10323 36576 10357
rect 36484 10289 36576 10323
rect 36484 10255 36511 10289
rect 36545 10255 36576 10289
rect 36484 10221 36576 10255
rect 36484 10187 36511 10221
rect 36545 10187 36576 10221
rect 36484 10153 36576 10187
rect 36484 10119 36511 10153
rect 36545 10119 36576 10153
rect 36484 10085 36576 10119
rect 36484 10051 36511 10085
rect 36545 10051 36576 10085
rect 36484 10017 36576 10051
rect 36484 9983 36511 10017
rect 36545 9983 36576 10017
rect 36484 9949 36576 9983
rect 36484 9915 36511 9949
rect 36545 9915 36576 9949
rect 36484 9881 36576 9915
rect 36484 9847 36511 9881
rect 36545 9847 36576 9881
rect 36484 9813 36576 9847
rect 36484 9779 36511 9813
rect 36545 9779 36576 9813
rect 36484 9745 36576 9779
rect 36484 9711 36511 9745
rect 36545 9711 36576 9745
rect 36484 9677 36576 9711
rect 36484 9643 36511 9677
rect 36545 9643 36576 9677
rect 36484 9609 36576 9643
rect 36484 9575 36511 9609
rect 36545 9575 36576 9609
rect 36484 9541 36576 9575
rect 37812 10534 37846 10553
rect 37812 10462 37846 10474
rect 37812 10390 37846 10406
rect 37812 10318 37846 10338
rect 37812 10246 37846 10270
rect 37812 10174 37846 10202
rect 37812 10102 37846 10134
rect 37812 10032 37846 10066
rect 37812 9964 37846 9996
rect 37812 9896 37846 9924
rect 37812 9828 37846 9852
rect 37812 9760 37846 9780
rect 37812 9692 37846 9708
rect 37812 9624 37846 9636
rect 37812 9545 37846 9564
rect 38070 10534 38104 10553
rect 38070 10462 38104 10474
rect 38070 10390 38104 10406
rect 38070 10318 38104 10338
rect 38070 10246 38104 10270
rect 38070 10174 38104 10202
rect 38070 10102 38104 10134
rect 38070 10032 38104 10066
rect 38070 9964 38104 9996
rect 38070 9896 38104 9924
rect 38070 9828 38104 9852
rect 38070 9760 38104 9780
rect 38070 9692 38104 9708
rect 38070 9624 38104 9636
rect 38070 9545 38104 9564
rect 38278 10534 38312 10553
rect 38278 10462 38312 10474
rect 38278 10390 38312 10406
rect 38278 10318 38312 10338
rect 38278 10246 38312 10270
rect 38278 10174 38312 10202
rect 38278 10102 38312 10134
rect 38278 10032 38312 10066
rect 38278 9964 38312 9996
rect 38278 9896 38312 9924
rect 38278 9828 38312 9852
rect 38278 9760 38312 9780
rect 38278 9692 38312 9708
rect 38278 9624 38312 9636
rect 38278 9545 38312 9564
rect 38536 10534 38570 10553
rect 38536 10462 38570 10474
rect 38536 10390 38570 10406
rect 38536 10318 38570 10338
rect 38536 10246 38570 10270
rect 38536 10174 38570 10202
rect 38536 10102 38570 10134
rect 38536 10032 38570 10066
rect 38536 9964 38570 9996
rect 38536 9896 38570 9924
rect 38536 9828 38570 9852
rect 38536 9760 38570 9780
rect 38536 9692 38570 9708
rect 38536 9624 38570 9636
rect 38536 9545 38570 9564
rect 38794 10534 38828 10553
rect 38794 10462 38828 10474
rect 38794 10390 38828 10406
rect 38794 10318 38828 10338
rect 38794 10246 38828 10270
rect 38794 10174 38828 10202
rect 38794 10102 38828 10134
rect 38794 10032 38828 10066
rect 38794 9964 38828 9996
rect 38794 9896 38828 9924
rect 38794 9828 38828 9852
rect 38794 9760 38828 9780
rect 38794 9692 38828 9708
rect 38794 9624 38828 9636
rect 38794 9545 38828 9564
rect 39052 10534 39086 10553
rect 39052 10462 39086 10474
rect 39052 10390 39086 10406
rect 39052 10318 39086 10338
rect 39052 10246 39086 10270
rect 39052 10174 39086 10202
rect 39052 10102 39086 10134
rect 39052 10032 39086 10066
rect 39052 9964 39086 9996
rect 39052 9896 39086 9924
rect 39052 9828 39086 9852
rect 39052 9760 39086 9780
rect 39052 9692 39086 9708
rect 39052 9624 39086 9636
rect 39052 9545 39086 9564
rect 39310 10534 39344 10553
rect 39310 10462 39344 10474
rect 39310 10390 39344 10406
rect 39310 10318 39344 10338
rect 39310 10246 39344 10270
rect 39310 10174 39344 10202
rect 39310 10102 39344 10134
rect 39310 10032 39344 10066
rect 39310 9964 39344 9996
rect 39310 9896 39344 9924
rect 39310 9828 39344 9852
rect 39310 9760 39344 9780
rect 39310 9692 39344 9708
rect 39310 9624 39344 9636
rect 39310 9545 39344 9564
rect 39568 10534 39602 10553
rect 39568 10462 39602 10474
rect 39568 10390 39602 10406
rect 39568 10318 39602 10338
rect 39568 10246 39602 10270
rect 39568 10174 39602 10202
rect 39568 10102 39602 10134
rect 39568 10032 39602 10066
rect 39568 9964 39602 9996
rect 39568 9896 39602 9924
rect 39568 9828 39602 9852
rect 39568 9760 39602 9780
rect 39568 9692 39602 9708
rect 39568 9624 39602 9636
rect 39568 9545 39602 9564
rect 39826 10534 39860 10553
rect 39826 10462 39860 10474
rect 39826 10390 39860 10406
rect 39826 10318 39860 10338
rect 39826 10246 39860 10270
rect 39826 10174 39860 10202
rect 39826 10102 39860 10134
rect 39826 10032 39860 10066
rect 39826 9964 39860 9996
rect 39826 9896 39860 9924
rect 39826 9828 39860 9852
rect 39826 9760 39860 9780
rect 39826 9692 39860 9708
rect 39826 9624 39860 9636
rect 39826 9545 39860 9564
rect 40084 10534 40118 10553
rect 40084 10462 40118 10474
rect 40084 10390 40118 10406
rect 40084 10318 40118 10338
rect 40084 10246 40118 10270
rect 40084 10174 40118 10202
rect 40084 10102 40118 10134
rect 40084 10032 40118 10066
rect 40084 9964 40118 9996
rect 40084 9896 40118 9924
rect 40084 9828 40118 9852
rect 40084 9760 40118 9780
rect 40084 9692 40118 9708
rect 40084 9624 40118 9636
rect 40084 9545 40118 9564
rect 40342 10534 40376 10553
rect 40342 10462 40376 10474
rect 40342 10390 40376 10406
rect 40342 10318 40376 10338
rect 40342 10246 40376 10270
rect 40342 10174 40376 10202
rect 40342 10102 40376 10134
rect 40342 10032 40376 10066
rect 40342 9964 40376 9996
rect 40342 9896 40376 9924
rect 40342 9828 40376 9852
rect 40342 9760 40376 9780
rect 40342 9692 40376 9708
rect 40342 9624 40376 9636
rect 40342 9545 40376 9564
rect 40600 10534 40634 10553
rect 40600 10462 40634 10474
rect 40600 10390 40634 10406
rect 40600 10318 40634 10338
rect 40600 10246 40634 10270
rect 40600 10174 40634 10202
rect 40600 10102 40634 10134
rect 40600 10032 40634 10066
rect 40600 9964 40634 9996
rect 40600 9896 40634 9924
rect 40600 9828 40634 9852
rect 40600 9760 40634 9780
rect 40600 9692 40634 9708
rect 40600 9624 40634 9636
rect 40600 9545 40634 9564
rect 40858 10534 40892 10553
rect 40858 10462 40892 10474
rect 40858 10390 40892 10406
rect 40858 10318 40892 10338
rect 40858 10246 40892 10270
rect 40858 10174 40892 10202
rect 40858 10102 40892 10134
rect 40858 10032 40892 10066
rect 40858 9964 40892 9996
rect 40858 9896 40892 9924
rect 40858 9828 40892 9852
rect 40858 9760 40892 9780
rect 40858 9692 40892 9708
rect 40858 9624 40892 9636
rect 40858 9545 40892 9564
rect 42203 10521 42303 10555
rect 42203 10487 42237 10521
rect 42271 10487 42303 10521
rect 42203 10453 42303 10487
rect 42203 10419 42237 10453
rect 42271 10419 42303 10453
rect 42203 10385 42303 10419
rect 42203 10351 42237 10385
rect 42271 10351 42303 10385
rect 42203 10317 42303 10351
rect 42203 10283 42237 10317
rect 42271 10283 42303 10317
rect 42203 10249 42303 10283
rect 42203 10215 42237 10249
rect 42271 10215 42303 10249
rect 42203 10181 42303 10215
rect 42203 10147 42237 10181
rect 42271 10147 42303 10181
rect 42203 10113 42303 10147
rect 42203 10079 42237 10113
rect 42271 10079 42303 10113
rect 42203 10045 42303 10079
rect 42203 10011 42237 10045
rect 42271 10011 42303 10045
rect 42203 9977 42303 10011
rect 42203 9943 42237 9977
rect 42271 9943 42303 9977
rect 42203 9909 42303 9943
rect 42203 9875 42237 9909
rect 42271 9875 42303 9909
rect 42203 9841 42303 9875
rect 42203 9807 42237 9841
rect 42271 9807 42303 9841
rect 42203 9773 42303 9807
rect 42203 9739 42237 9773
rect 42271 9739 42303 9773
rect 42203 9705 42303 9739
rect 42203 9671 42237 9705
rect 42271 9671 42303 9705
rect 42203 9637 42303 9671
rect 42203 9603 42237 9637
rect 42271 9603 42303 9637
rect 42203 9569 42303 9603
rect 36484 9507 36511 9541
rect 36545 9507 36576 9541
rect 42203 9535 42237 9569
rect 42271 9535 42303 9569
rect 36484 9473 36576 9507
rect 37858 9477 37905 9511
rect 37941 9477 37975 9511
rect 38011 9477 38058 9511
rect 38324 9477 38371 9511
rect 38407 9477 38441 9511
rect 38477 9477 38524 9511
rect 38582 9477 38629 9511
rect 38665 9477 38699 9511
rect 38735 9477 38782 9511
rect 38840 9477 38887 9511
rect 38923 9477 38957 9511
rect 38993 9477 39040 9511
rect 39098 9477 39145 9511
rect 39181 9477 39215 9511
rect 39251 9477 39298 9511
rect 39356 9477 39403 9511
rect 39439 9477 39473 9511
rect 39509 9477 39556 9511
rect 39614 9477 39661 9511
rect 39697 9477 39731 9511
rect 39767 9477 39814 9511
rect 39872 9477 39919 9511
rect 39955 9477 39989 9511
rect 40025 9477 40072 9511
rect 40130 9477 40177 9511
rect 40213 9477 40247 9511
rect 40283 9477 40330 9511
rect 40388 9477 40435 9511
rect 40471 9477 40505 9511
rect 40541 9477 40588 9511
rect 40646 9477 40693 9511
rect 40729 9477 40763 9511
rect 40799 9477 40846 9511
rect 42203 9501 42303 9535
rect 36484 9439 36511 9473
rect 36545 9439 36576 9473
rect 36484 9405 36576 9439
rect 36484 9371 36511 9405
rect 36545 9371 36576 9405
rect 36484 9179 36576 9371
rect 42203 9467 42237 9501
rect 42271 9467 42303 9501
rect 42203 9433 42303 9467
rect 42203 9399 42237 9433
rect 42271 9399 42303 9433
rect 42203 9365 42303 9399
rect 42203 9331 42237 9365
rect 42271 9331 42303 9365
rect 42203 9179 42303 9331
rect 36484 9149 42303 9179
rect 36484 9115 36779 9149
rect 36813 9115 36847 9149
rect 36881 9115 36915 9149
rect 36949 9115 36983 9149
rect 37017 9115 37051 9149
rect 37085 9115 37119 9149
rect 37153 9115 37187 9149
rect 37221 9115 37255 9149
rect 37289 9115 37323 9149
rect 37357 9115 37391 9149
rect 37425 9115 37459 9149
rect 37493 9115 37527 9149
rect 37561 9115 37595 9149
rect 37629 9115 37663 9149
rect 37697 9115 37731 9149
rect 37765 9115 37799 9149
rect 37833 9115 37867 9149
rect 37901 9115 37935 9149
rect 37969 9115 38003 9149
rect 38037 9115 38071 9149
rect 38105 9115 38139 9149
rect 38173 9115 38207 9149
rect 38241 9115 38275 9149
rect 38309 9115 38343 9149
rect 38377 9115 38411 9149
rect 38445 9115 38479 9149
rect 38513 9115 38547 9149
rect 38581 9115 38615 9149
rect 38649 9115 38683 9149
rect 38717 9115 38751 9149
rect 38785 9115 38819 9149
rect 38853 9115 38887 9149
rect 38921 9115 38955 9149
rect 38989 9115 39023 9149
rect 39057 9115 39091 9149
rect 39125 9115 39159 9149
rect 39193 9115 39227 9149
rect 39261 9115 39295 9149
rect 39329 9115 39363 9149
rect 39397 9115 39431 9149
rect 39465 9115 39499 9149
rect 39533 9115 39567 9149
rect 39601 9115 39635 9149
rect 39669 9115 39703 9149
rect 39737 9115 39771 9149
rect 39805 9115 39839 9149
rect 39873 9115 39907 9149
rect 39941 9115 39975 9149
rect 40009 9115 40043 9149
rect 40077 9115 40111 9149
rect 40145 9115 40179 9149
rect 40213 9115 40247 9149
rect 40281 9115 40315 9149
rect 40349 9115 40383 9149
rect 40417 9115 40451 9149
rect 40485 9115 40519 9149
rect 40553 9115 40587 9149
rect 40621 9115 40655 9149
rect 40689 9115 40723 9149
rect 40757 9115 40791 9149
rect 40825 9115 40859 9149
rect 40893 9115 40927 9149
rect 40961 9115 40995 9149
rect 41029 9115 41063 9149
rect 41097 9115 41131 9149
rect 41165 9115 41199 9149
rect 41233 9115 41267 9149
rect 41301 9115 41335 9149
rect 41369 9115 41403 9149
rect 41437 9115 41471 9149
rect 41505 9115 41539 9149
rect 41573 9115 41607 9149
rect 41641 9115 41675 9149
rect 41709 9115 41743 9149
rect 41777 9115 41811 9149
rect 41845 9115 41879 9149
rect 41913 9115 41947 9149
rect 41981 9115 42015 9149
rect 42049 9115 42303 9149
rect 36484 9087 44191 9115
rect 36484 9086 36576 9087
rect 29774 8995 29808 9029
rect 29774 8927 29808 8961
rect 29774 8859 29808 8893
rect 29774 8791 29808 8825
rect 29774 8723 29808 8757
rect 29774 8655 29808 8689
rect 29774 8587 29808 8621
rect 29774 8519 29808 8553
rect 29774 8451 29808 8485
rect 29774 8383 29808 8417
rect 29774 8315 29808 8349
rect 29774 8247 29808 8281
rect 29774 8179 29808 8213
rect 29774 8111 29808 8145
rect 29774 8043 29808 8077
rect 29774 7975 29808 8009
rect 29774 7907 29808 7941
rect 29774 7839 29808 7873
rect 29774 7771 29808 7805
rect 29774 7703 29808 7737
rect 29774 7635 29808 7669
rect 29774 7567 29808 7601
rect 29774 7499 29808 7533
rect 29774 7431 29808 7465
rect 29774 7363 29808 7397
rect 29774 7295 29808 7329
rect 29774 7227 29808 7261
rect 29774 7159 29808 7193
rect 29774 7091 29808 7125
rect 29774 7023 29808 7057
rect 29774 6955 29808 6989
rect 29774 6900 29808 6921
rect 27364 6896 27774 6898
rect 29608 6896 29808 6900
rect 27364 6887 27700 6896
rect 27364 6869 27570 6887
rect 27318 6853 27570 6869
rect 27604 6853 27700 6887
rect 27318 6835 27700 6853
rect 27318 6801 27330 6835
rect 27364 6819 27700 6835
rect 27364 6801 27570 6819
rect 27318 6785 27570 6801
rect 27604 6785 27700 6819
rect 27318 6767 27700 6785
rect 27318 6733 27330 6767
rect 27364 6751 27700 6767
rect 27364 6733 27570 6751
rect 27318 6717 27570 6733
rect 27604 6717 27700 6751
rect 27318 6699 27700 6717
rect 27318 6665 27330 6699
rect 27364 6683 27700 6699
rect 27364 6665 27570 6683
rect 27318 6649 27570 6665
rect 27604 6649 27700 6683
rect 27318 6631 27700 6649
rect 27318 6597 27330 6631
rect 27364 6615 27700 6631
rect 27364 6597 27570 6615
rect 27318 6581 27570 6597
rect 27604 6581 27700 6615
rect 27318 6563 27700 6581
rect 27318 6529 27330 6563
rect 27364 6547 27700 6563
rect 27364 6529 27570 6547
rect 27318 6513 27570 6529
rect 27604 6513 27700 6547
rect 27318 6495 27700 6513
rect 27318 6468 27330 6495
rect 26398 6427 26432 6461
rect 26398 6359 26432 6393
rect 26398 6291 26432 6325
rect 26398 6223 26432 6257
rect 26398 6155 26432 6189
rect 26398 6087 26432 6121
rect 26398 6019 26432 6053
rect 26398 5951 26432 5985
rect 26398 5883 26432 5917
rect 26398 5815 26432 5849
rect 26398 5747 26432 5781
rect 26398 5679 26432 5713
rect 26398 5611 26432 5645
rect 26398 5543 26432 5577
rect 26398 5475 26432 5509
rect 26398 5407 26432 5441
rect 26398 5339 26432 5373
rect 26398 5271 26432 5305
rect 26398 5203 26432 5237
rect 26398 5135 26432 5169
rect 26398 5067 26432 5101
rect 26398 4999 26432 5033
rect 26398 4931 26432 4965
rect 26398 4863 26432 4897
rect 26398 4795 26432 4829
rect 26398 4727 26432 4761
rect 26398 4659 26432 4693
rect 26398 4591 26432 4625
rect 26398 4523 26432 4557
rect 26398 4455 26432 4489
rect 26398 4387 26432 4421
rect 26398 4319 26432 4353
rect 26398 4251 26432 4285
rect 26398 4183 26432 4217
rect 26398 4115 26432 4149
rect 26398 4047 26432 4081
rect 26398 3979 26432 4013
rect 26398 3911 26432 3945
rect 26398 3843 26432 3877
rect 26398 3775 26432 3809
rect 26398 3707 26432 3741
rect 26398 3639 26432 3673
rect 26398 3571 26432 3605
rect 22376 3537 26398 3552
rect 22376 3514 26432 3537
rect 22376 3480 23515 3514
rect 23549 3480 23583 3514
rect 23617 3480 23651 3514
rect 23685 3480 23719 3514
rect 23753 3480 23787 3514
rect 23821 3480 23855 3514
rect 23889 3480 23923 3514
rect 23957 3480 23991 3514
rect 24025 3480 24059 3514
rect 24093 3480 24127 3514
rect 24161 3480 24195 3514
rect 24229 3480 24263 3514
rect 24297 3480 24331 3514
rect 24365 3504 24399 3514
rect 24433 3504 24467 3514
rect 24365 3480 24389 3504
rect 24433 3480 24461 3504
rect 24501 3480 24535 3514
rect 24569 3480 24603 3514
rect 24637 3480 24671 3514
rect 24705 3480 25015 3514
rect 25049 3480 25083 3514
rect 25117 3480 25151 3514
rect 25185 3480 25219 3514
rect 25253 3480 25287 3514
rect 25321 3480 25355 3514
rect 25389 3480 25423 3514
rect 25457 3480 25491 3514
rect 25525 3480 25559 3514
rect 25593 3480 25627 3514
rect 25661 3480 25695 3514
rect 25729 3480 25763 3514
rect 25797 3480 25831 3514
rect 25865 3480 25899 3514
rect 25933 3480 25967 3514
rect 26001 3480 26035 3514
rect 26069 3480 26103 3514
rect 26137 3480 26171 3514
rect 26205 3503 26432 3514
rect 27364 6479 27700 6495
rect 27364 6468 27570 6479
rect 27330 6427 27364 6461
rect 27330 6359 27364 6393
rect 27604 6468 27700 6479
rect 27770 6468 27774 6896
rect 29678 6887 29808 6896
rect 29678 6853 29774 6887
rect 29678 6819 29808 6853
rect 29678 6785 29774 6819
rect 29678 6751 29808 6785
rect 29678 6717 29774 6751
rect 29678 6683 29808 6717
rect 29678 6649 29774 6683
rect 29678 6615 29808 6649
rect 29678 6581 29774 6615
rect 29678 6547 29808 6581
rect 29678 6513 29774 6547
rect 29678 6479 29808 6513
rect 29678 6470 29774 6479
rect 27570 6368 27604 6445
rect 29774 6368 29808 6445
rect 27570 6334 27686 6368
rect 27720 6334 27754 6368
rect 27788 6334 27822 6368
rect 27856 6334 27890 6368
rect 27924 6334 27958 6368
rect 27992 6334 28026 6368
rect 28060 6334 28094 6368
rect 28128 6334 28162 6368
rect 28196 6334 28230 6368
rect 28264 6334 28298 6368
rect 28332 6334 28366 6368
rect 28400 6334 28434 6368
rect 28468 6334 28502 6368
rect 28536 6334 28570 6368
rect 28604 6334 28638 6368
rect 28672 6334 28706 6368
rect 28740 6334 28774 6368
rect 28808 6334 28842 6368
rect 28876 6334 28910 6368
rect 28944 6334 28978 6368
rect 29012 6334 29046 6368
rect 29080 6334 29114 6368
rect 29148 6334 29182 6368
rect 29216 6334 29250 6368
rect 29284 6334 29318 6368
rect 29352 6334 29386 6368
rect 29420 6334 29454 6368
rect 29488 6334 29522 6368
rect 29556 6334 29590 6368
rect 29624 6334 29658 6368
rect 29692 6334 29808 6368
rect 37608 8609 44191 9087
rect 37608 8575 37843 8609
rect 37877 8575 37911 8609
rect 37945 8575 37979 8609
rect 38013 8575 38047 8609
rect 38081 8575 38115 8609
rect 38149 8575 38183 8609
rect 38217 8575 38251 8609
rect 38285 8575 38319 8609
rect 38353 8575 38387 8609
rect 38421 8575 38455 8609
rect 38489 8575 38523 8609
rect 38557 8575 38591 8609
rect 38625 8575 38659 8609
rect 38693 8575 38727 8609
rect 38761 8575 38795 8609
rect 38829 8575 38863 8609
rect 38897 8575 38931 8609
rect 38965 8575 38999 8609
rect 39033 8575 39067 8609
rect 39101 8575 39135 8609
rect 39169 8575 39203 8609
rect 39237 8575 39271 8609
rect 39305 8575 39339 8609
rect 39373 8575 39407 8609
rect 39441 8575 39475 8609
rect 39509 8575 39543 8609
rect 39577 8575 39611 8609
rect 39645 8575 39679 8609
rect 39713 8575 39747 8609
rect 39781 8575 39815 8609
rect 39849 8575 39883 8609
rect 39917 8575 39951 8609
rect 39985 8575 40019 8609
rect 40053 8575 40087 8609
rect 40121 8575 40155 8609
rect 40189 8575 40223 8609
rect 40257 8575 40291 8609
rect 40325 8575 40359 8609
rect 40393 8575 40427 8609
rect 40461 8575 40495 8609
rect 40529 8575 40563 8609
rect 40597 8575 40631 8609
rect 40665 8575 40699 8609
rect 40733 8575 40767 8609
rect 40801 8575 40835 8609
rect 40869 8575 40903 8609
rect 40937 8575 40971 8609
rect 41005 8575 41039 8609
rect 41073 8575 41107 8609
rect 41141 8575 41175 8609
rect 41209 8575 41243 8609
rect 41277 8575 41311 8609
rect 41345 8575 41379 8609
rect 41413 8575 41447 8609
rect 41481 8575 41515 8609
rect 41549 8575 41583 8609
rect 41617 8575 41651 8609
rect 41685 8575 41719 8609
rect 41753 8575 41787 8609
rect 41821 8575 41855 8609
rect 41889 8575 41923 8609
rect 41957 8575 41991 8609
rect 42025 8575 42184 8609
rect 37608 8564 42184 8575
rect 37608 8432 37674 8564
rect 37608 8398 37624 8432
rect 37658 8398 37674 8432
rect 37608 8364 37674 8398
rect 37608 8330 37624 8364
rect 37658 8330 37674 8364
rect 42122 8444 42184 8564
rect 42122 8410 42136 8444
rect 42170 8410 42184 8444
rect 42122 8376 42184 8410
rect 37608 8296 37674 8330
rect 37858 8326 37905 8360
rect 37941 8326 37975 8360
rect 38011 8326 38058 8360
rect 38116 8326 38163 8360
rect 38199 8326 38233 8360
rect 38269 8326 38316 8360
rect 38374 8326 38421 8360
rect 38457 8326 38491 8360
rect 38527 8326 38574 8360
rect 38632 8326 38679 8360
rect 38715 8326 38749 8360
rect 38785 8326 38832 8360
rect 38890 8326 38937 8360
rect 38973 8326 39007 8360
rect 39043 8326 39090 8360
rect 39148 8326 39195 8360
rect 39231 8326 39265 8360
rect 39301 8326 39348 8360
rect 39406 8326 39453 8360
rect 39489 8326 39523 8360
rect 39559 8326 39606 8360
rect 39664 8326 39711 8360
rect 39747 8326 39781 8360
rect 39817 8326 39864 8360
rect 39922 8326 39969 8360
rect 40005 8326 40039 8360
rect 40075 8326 40122 8360
rect 40180 8326 40227 8360
rect 40263 8326 40297 8360
rect 40333 8326 40380 8360
rect 40438 8326 40485 8360
rect 40521 8326 40555 8360
rect 40591 8326 40638 8360
rect 40696 8326 40743 8360
rect 40779 8326 40813 8360
rect 40849 8326 40896 8360
rect 40954 8326 41001 8360
rect 41037 8326 41071 8360
rect 41107 8326 41154 8360
rect 41212 8326 41259 8360
rect 41295 8326 41329 8360
rect 41365 8326 41412 8360
rect 41470 8326 41517 8360
rect 41553 8326 41587 8360
rect 41623 8326 41670 8360
rect 41728 8326 41775 8360
rect 41811 8326 41845 8360
rect 41881 8326 41928 8360
rect 42122 8342 42136 8376
rect 42170 8342 42184 8376
rect 37608 8262 37624 8296
rect 37658 8262 37674 8296
rect 42122 8308 42184 8342
rect 37608 8228 37674 8262
rect 37608 8194 37624 8228
rect 37658 8194 37674 8228
rect 37608 8160 37674 8194
rect 37608 8126 37624 8160
rect 37658 8126 37674 8160
rect 37608 8092 37674 8126
rect 37608 8058 37624 8092
rect 37658 8058 37674 8092
rect 37608 8024 37674 8058
rect 37608 7990 37624 8024
rect 37658 7990 37674 8024
rect 37608 7956 37674 7990
rect 37608 7922 37624 7956
rect 37658 7922 37674 7956
rect 37608 7888 37674 7922
rect 37608 7854 37624 7888
rect 37658 7854 37674 7888
rect 37608 7820 37674 7854
rect 37608 7786 37624 7820
rect 37658 7786 37674 7820
rect 37608 7752 37674 7786
rect 37608 7718 37624 7752
rect 37658 7718 37674 7752
rect 37608 7684 37674 7718
rect 37608 7650 37624 7684
rect 37658 7650 37674 7684
rect 37608 7616 37674 7650
rect 37608 7582 37624 7616
rect 37658 7582 37674 7616
rect 37608 7548 37674 7582
rect 37608 7514 37624 7548
rect 37658 7514 37674 7548
rect 37608 7480 37674 7514
rect 37608 7446 37624 7480
rect 37658 7446 37674 7480
rect 37608 7412 37674 7446
rect 37608 7378 37624 7412
rect 37658 7378 37674 7412
rect 37608 7344 37674 7378
rect 37608 7310 37624 7344
rect 37658 7310 37674 7344
rect 37608 7276 37674 7310
rect 37608 7242 37624 7276
rect 37658 7242 37674 7276
rect 37608 7208 37674 7242
rect 37608 7174 37624 7208
rect 37658 7174 37674 7208
rect 37608 7140 37674 7174
rect 37608 7106 37624 7140
rect 37658 7106 37674 7140
rect 37608 7072 37674 7106
rect 37608 7038 37624 7072
rect 37658 7038 37674 7072
rect 37608 7004 37674 7038
rect 37608 6970 37624 7004
rect 37658 6970 37674 7004
rect 37608 6936 37674 6970
rect 37608 6902 37624 6936
rect 37658 6902 37674 6936
rect 37608 6868 37674 6902
rect 37608 6834 37624 6868
rect 37658 6834 37674 6868
rect 37608 6800 37674 6834
rect 37608 6766 37624 6800
rect 37658 6766 37674 6800
rect 37608 6732 37674 6766
rect 37608 6698 37624 6732
rect 37658 6698 37674 6732
rect 37608 6664 37674 6698
rect 37608 6636 37624 6664
rect 37608 6602 37623 6636
rect 37658 6630 37674 6664
rect 37657 6602 37674 6630
rect 37608 6596 37674 6602
rect 37608 6564 37624 6596
rect 37608 6530 37623 6564
rect 37658 6562 37674 6596
rect 37657 6530 37674 6562
rect 37608 6528 37674 6530
rect 37608 6494 37624 6528
rect 37658 6494 37674 6528
rect 37608 6492 37674 6494
rect 37608 6458 37623 6492
rect 37657 6460 37674 6492
rect 37608 6426 37624 6458
rect 37658 6426 37674 6460
rect 37608 6392 37674 6426
rect 37608 6358 37624 6392
rect 37658 6358 37674 6392
rect 27330 6291 27364 6325
rect 27330 6223 27364 6257
rect 27330 6155 27364 6189
rect 27330 6087 27364 6121
rect 27330 6019 27364 6053
rect 37608 6324 37674 6358
rect 37608 6290 37624 6324
rect 37658 6290 37674 6324
rect 37608 6256 37674 6290
rect 37812 8257 37846 8292
rect 37812 8189 37846 8207
rect 37812 8121 37846 8135
rect 37812 8053 37846 8063
rect 37812 7985 37846 7991
rect 37812 7917 37846 7919
rect 37812 7881 37846 7883
rect 37812 7809 37846 7815
rect 37812 7737 37846 7747
rect 37812 7665 37846 7679
rect 37812 7593 37846 7611
rect 37812 7521 37846 7543
rect 37812 7449 37846 7475
rect 37812 7377 37846 7407
rect 37812 7305 37846 7339
rect 37812 7237 37846 7271
rect 37812 7169 37846 7199
rect 37812 7101 37846 7127
rect 37812 7033 37846 7055
rect 37812 6965 37846 6983
rect 37812 6897 37846 6911
rect 37812 6829 37846 6839
rect 37812 6761 37846 6767
rect 37812 6693 37846 6695
rect 37812 6657 37846 6659
rect 37812 6585 37846 6591
rect 37812 6513 37846 6523
rect 37812 6441 37846 6455
rect 37812 6369 37846 6387
rect 37812 6284 37846 6319
rect 38070 8257 38104 8292
rect 38070 8189 38104 8207
rect 38070 8121 38104 8135
rect 38070 8053 38104 8063
rect 38070 7985 38104 7991
rect 38070 7917 38104 7919
rect 38070 7881 38104 7883
rect 38070 7809 38104 7815
rect 38070 7737 38104 7747
rect 38070 7665 38104 7679
rect 38070 7593 38104 7611
rect 38070 7521 38104 7543
rect 38070 7449 38104 7475
rect 38070 7377 38104 7407
rect 38070 7305 38104 7339
rect 38070 7237 38104 7271
rect 38070 7169 38104 7199
rect 38070 7101 38104 7127
rect 38070 7033 38104 7055
rect 38070 6965 38104 6983
rect 38070 6897 38104 6911
rect 38070 6829 38104 6839
rect 38070 6761 38104 6767
rect 38070 6693 38104 6695
rect 38070 6657 38104 6659
rect 38070 6585 38104 6591
rect 38070 6513 38104 6523
rect 38070 6441 38104 6455
rect 38070 6369 38104 6387
rect 38070 6284 38104 6319
rect 38328 8257 38362 8292
rect 38328 8189 38362 8207
rect 38328 8121 38362 8135
rect 38328 8053 38362 8063
rect 38328 7985 38362 7991
rect 38328 7917 38362 7919
rect 38328 7881 38362 7883
rect 38328 7809 38362 7815
rect 38328 7737 38362 7747
rect 38328 7665 38362 7679
rect 38328 7593 38362 7611
rect 38328 7521 38362 7543
rect 38328 7449 38362 7475
rect 38328 7377 38362 7407
rect 38328 7305 38362 7339
rect 38328 7237 38362 7271
rect 38328 7169 38362 7199
rect 38328 7101 38362 7127
rect 38328 7033 38362 7055
rect 38328 6965 38362 6983
rect 38328 6897 38362 6911
rect 38328 6829 38362 6839
rect 38328 6761 38362 6767
rect 38328 6693 38362 6695
rect 38328 6657 38362 6659
rect 38328 6585 38362 6591
rect 38328 6513 38362 6523
rect 38328 6441 38362 6455
rect 38328 6369 38362 6387
rect 38328 6284 38362 6319
rect 38586 8257 38620 8292
rect 38586 8189 38620 8207
rect 38586 8121 38620 8135
rect 38586 8053 38620 8063
rect 38586 7985 38620 7991
rect 38586 7917 38620 7919
rect 38586 7881 38620 7883
rect 38586 7809 38620 7815
rect 38586 7737 38620 7747
rect 38586 7665 38620 7679
rect 38586 7593 38620 7611
rect 38586 7521 38620 7543
rect 38586 7449 38620 7475
rect 38586 7377 38620 7407
rect 38586 7305 38620 7339
rect 38586 7237 38620 7271
rect 38586 7169 38620 7199
rect 38586 7101 38620 7127
rect 38586 7033 38620 7055
rect 38586 6965 38620 6983
rect 38586 6897 38620 6911
rect 38586 6829 38620 6839
rect 38586 6761 38620 6767
rect 38586 6693 38620 6695
rect 38586 6657 38620 6659
rect 38586 6585 38620 6591
rect 38586 6513 38620 6523
rect 38586 6441 38620 6455
rect 38586 6369 38620 6387
rect 38586 6284 38620 6319
rect 38844 8257 38878 8292
rect 38844 8189 38878 8207
rect 38844 8121 38878 8135
rect 38844 8053 38878 8063
rect 38844 7985 38878 7991
rect 38844 7917 38878 7919
rect 38844 7881 38878 7883
rect 38844 7809 38878 7815
rect 38844 7737 38878 7747
rect 38844 7665 38878 7679
rect 38844 7593 38878 7611
rect 38844 7521 38878 7543
rect 38844 7449 38878 7475
rect 38844 7377 38878 7407
rect 38844 7305 38878 7339
rect 38844 7237 38878 7271
rect 38844 7169 38878 7199
rect 38844 7101 38878 7127
rect 38844 7033 38878 7055
rect 38844 6965 38878 6983
rect 38844 6897 38878 6911
rect 38844 6829 38878 6839
rect 38844 6761 38878 6767
rect 38844 6693 38878 6695
rect 38844 6657 38878 6659
rect 38844 6585 38878 6591
rect 38844 6513 38878 6523
rect 38844 6441 38878 6455
rect 38844 6369 38878 6387
rect 38844 6284 38878 6319
rect 39102 8257 39136 8292
rect 39102 8189 39136 8207
rect 39102 8121 39136 8135
rect 39102 8053 39136 8063
rect 39102 7985 39136 7991
rect 39102 7917 39136 7919
rect 39102 7881 39136 7883
rect 39102 7809 39136 7815
rect 39102 7737 39136 7747
rect 39102 7665 39136 7679
rect 39102 7593 39136 7611
rect 39102 7521 39136 7543
rect 39102 7449 39136 7475
rect 39102 7377 39136 7407
rect 39102 7305 39136 7339
rect 39102 7237 39136 7271
rect 39102 7169 39136 7199
rect 39102 7101 39136 7127
rect 39102 7033 39136 7055
rect 39102 6965 39136 6983
rect 39102 6897 39136 6911
rect 39102 6829 39136 6839
rect 39102 6761 39136 6767
rect 39102 6693 39136 6695
rect 39102 6657 39136 6659
rect 39102 6585 39136 6591
rect 39102 6513 39136 6523
rect 39102 6441 39136 6455
rect 39102 6369 39136 6387
rect 39102 6284 39136 6319
rect 39360 8257 39394 8292
rect 39360 8189 39394 8207
rect 39360 8121 39394 8135
rect 39360 8053 39394 8063
rect 39360 7985 39394 7991
rect 39360 7917 39394 7919
rect 39360 7881 39394 7883
rect 39360 7809 39394 7815
rect 39360 7737 39394 7747
rect 39360 7665 39394 7679
rect 39360 7593 39394 7611
rect 39360 7521 39394 7543
rect 39360 7449 39394 7475
rect 39360 7377 39394 7407
rect 39360 7305 39394 7339
rect 39360 7237 39394 7271
rect 39360 7169 39394 7199
rect 39360 7101 39394 7127
rect 39360 7033 39394 7055
rect 39360 6965 39394 6983
rect 39360 6897 39394 6911
rect 39360 6829 39394 6839
rect 39360 6761 39394 6767
rect 39360 6693 39394 6695
rect 39360 6657 39394 6659
rect 39360 6585 39394 6591
rect 39360 6513 39394 6523
rect 39360 6441 39394 6455
rect 39360 6369 39394 6387
rect 39360 6284 39394 6319
rect 39618 8257 39652 8292
rect 39618 8189 39652 8207
rect 39618 8121 39652 8135
rect 39618 8053 39652 8063
rect 39618 7985 39652 7991
rect 39618 7917 39652 7919
rect 39618 7881 39652 7883
rect 39618 7809 39652 7815
rect 39618 7737 39652 7747
rect 39618 7665 39652 7679
rect 39618 7593 39652 7611
rect 39618 7521 39652 7543
rect 39618 7449 39652 7475
rect 39618 7377 39652 7407
rect 39618 7305 39652 7339
rect 39618 7237 39652 7271
rect 39618 7169 39652 7199
rect 39618 7101 39652 7127
rect 39618 7033 39652 7055
rect 39618 6965 39652 6983
rect 39618 6897 39652 6911
rect 39618 6829 39652 6839
rect 39618 6761 39652 6767
rect 39618 6693 39652 6695
rect 39618 6657 39652 6659
rect 39618 6585 39652 6591
rect 39618 6513 39652 6523
rect 39618 6441 39652 6455
rect 39618 6369 39652 6387
rect 39618 6284 39652 6319
rect 39876 8257 39910 8292
rect 39876 8189 39910 8207
rect 39876 8121 39910 8135
rect 39876 8053 39910 8063
rect 39876 7985 39910 7991
rect 39876 7917 39910 7919
rect 39876 7881 39910 7883
rect 39876 7809 39910 7815
rect 39876 7737 39910 7747
rect 39876 7665 39910 7679
rect 39876 7593 39910 7611
rect 39876 7521 39910 7543
rect 39876 7449 39910 7475
rect 39876 7377 39910 7407
rect 39876 7305 39910 7339
rect 39876 7237 39910 7271
rect 39876 7169 39910 7199
rect 39876 7101 39910 7127
rect 39876 7033 39910 7055
rect 39876 6965 39910 6983
rect 39876 6897 39910 6911
rect 39876 6829 39910 6839
rect 39876 6761 39910 6767
rect 39876 6693 39910 6695
rect 39876 6657 39910 6659
rect 39876 6585 39910 6591
rect 39876 6513 39910 6523
rect 39876 6441 39910 6455
rect 39876 6369 39910 6387
rect 39876 6284 39910 6319
rect 40134 8257 40168 8292
rect 40134 8189 40168 8207
rect 40134 8121 40168 8135
rect 40134 8053 40168 8063
rect 40134 7985 40168 7991
rect 40134 7917 40168 7919
rect 40134 7881 40168 7883
rect 40134 7809 40168 7815
rect 40134 7737 40168 7747
rect 40134 7665 40168 7679
rect 40134 7593 40168 7611
rect 40134 7521 40168 7543
rect 40134 7449 40168 7475
rect 40134 7377 40168 7407
rect 40134 7305 40168 7339
rect 40134 7237 40168 7271
rect 40134 7169 40168 7199
rect 40134 7101 40168 7127
rect 40134 7033 40168 7055
rect 40134 6965 40168 6983
rect 40134 6897 40168 6911
rect 40134 6829 40168 6839
rect 40134 6761 40168 6767
rect 40134 6693 40168 6695
rect 40134 6657 40168 6659
rect 40134 6585 40168 6591
rect 40134 6513 40168 6523
rect 40134 6441 40168 6455
rect 40134 6369 40168 6387
rect 40134 6284 40168 6319
rect 40392 8257 40426 8292
rect 40392 8189 40426 8207
rect 40392 8121 40426 8135
rect 40392 8053 40426 8063
rect 40392 7985 40426 7991
rect 40392 7917 40426 7919
rect 40392 7881 40426 7883
rect 40392 7809 40426 7815
rect 40392 7737 40426 7747
rect 40392 7665 40426 7679
rect 40392 7593 40426 7611
rect 40392 7521 40426 7543
rect 40392 7449 40426 7475
rect 40392 7377 40426 7407
rect 40392 7305 40426 7339
rect 40392 7237 40426 7271
rect 40392 7169 40426 7199
rect 40392 7101 40426 7127
rect 40392 7033 40426 7055
rect 40392 6965 40426 6983
rect 40392 6897 40426 6911
rect 40392 6829 40426 6839
rect 40392 6761 40426 6767
rect 40392 6693 40426 6695
rect 40392 6657 40426 6659
rect 40392 6585 40426 6591
rect 40392 6513 40426 6523
rect 40392 6441 40426 6455
rect 40392 6369 40426 6387
rect 40392 6284 40426 6319
rect 40650 8257 40684 8292
rect 40650 8189 40684 8207
rect 40650 8121 40684 8135
rect 40650 8053 40684 8063
rect 40650 7985 40684 7991
rect 40650 7917 40684 7919
rect 40650 7881 40684 7883
rect 40650 7809 40684 7815
rect 40650 7737 40684 7747
rect 40650 7665 40684 7679
rect 40650 7593 40684 7611
rect 40650 7521 40684 7543
rect 40650 7449 40684 7475
rect 40650 7377 40684 7407
rect 40650 7305 40684 7339
rect 40650 7237 40684 7271
rect 40650 7169 40684 7199
rect 40650 7101 40684 7127
rect 40650 7033 40684 7055
rect 40650 6965 40684 6983
rect 40650 6897 40684 6911
rect 40650 6829 40684 6839
rect 40650 6761 40684 6767
rect 40650 6693 40684 6695
rect 40650 6657 40684 6659
rect 40650 6585 40684 6591
rect 40650 6513 40684 6523
rect 40650 6441 40684 6455
rect 40650 6369 40684 6387
rect 40650 6284 40684 6319
rect 40908 8257 40942 8292
rect 40908 8189 40942 8207
rect 40908 8121 40942 8135
rect 40908 8053 40942 8063
rect 40908 7985 40942 7991
rect 40908 7917 40942 7919
rect 40908 7881 40942 7883
rect 40908 7809 40942 7815
rect 40908 7737 40942 7747
rect 40908 7665 40942 7679
rect 40908 7593 40942 7611
rect 40908 7521 40942 7543
rect 40908 7449 40942 7475
rect 40908 7377 40942 7407
rect 40908 7305 40942 7339
rect 40908 7237 40942 7271
rect 40908 7169 40942 7199
rect 40908 7101 40942 7127
rect 40908 7033 40942 7055
rect 40908 6965 40942 6983
rect 40908 6897 40942 6911
rect 40908 6829 40942 6839
rect 40908 6761 40942 6767
rect 40908 6693 40942 6695
rect 40908 6657 40942 6659
rect 40908 6585 40942 6591
rect 40908 6513 40942 6523
rect 40908 6441 40942 6455
rect 40908 6369 40942 6387
rect 40908 6284 40942 6319
rect 41166 8257 41200 8292
rect 41166 8189 41200 8207
rect 41166 8121 41200 8135
rect 41166 8053 41200 8063
rect 41166 7985 41200 7991
rect 41166 7917 41200 7919
rect 41166 7881 41200 7883
rect 41166 7809 41200 7815
rect 41166 7737 41200 7747
rect 41166 7665 41200 7679
rect 41166 7593 41200 7611
rect 41166 7521 41200 7543
rect 41166 7449 41200 7475
rect 41166 7377 41200 7407
rect 41166 7305 41200 7339
rect 41166 7237 41200 7271
rect 41166 7169 41200 7199
rect 41166 7101 41200 7127
rect 41166 7033 41200 7055
rect 41166 6965 41200 6983
rect 41166 6897 41200 6911
rect 41166 6829 41200 6839
rect 41166 6761 41200 6767
rect 41166 6693 41200 6695
rect 41166 6657 41200 6659
rect 41166 6585 41200 6591
rect 41166 6513 41200 6523
rect 41166 6441 41200 6455
rect 41166 6369 41200 6387
rect 41166 6284 41200 6319
rect 41424 8257 41458 8292
rect 41424 8189 41458 8207
rect 41424 8121 41458 8135
rect 41424 8053 41458 8063
rect 41424 7985 41458 7991
rect 41424 7917 41458 7919
rect 41424 7881 41458 7883
rect 41424 7809 41458 7815
rect 41424 7737 41458 7747
rect 41424 7665 41458 7679
rect 41424 7593 41458 7611
rect 41424 7521 41458 7543
rect 41424 7449 41458 7475
rect 41424 7377 41458 7407
rect 41424 7305 41458 7339
rect 41424 7237 41458 7271
rect 41424 7169 41458 7199
rect 41424 7101 41458 7127
rect 41424 7033 41458 7055
rect 41424 6965 41458 6983
rect 41424 6897 41458 6911
rect 41424 6829 41458 6839
rect 41424 6761 41458 6767
rect 41424 6693 41458 6695
rect 41424 6657 41458 6659
rect 41424 6585 41458 6591
rect 41424 6513 41458 6523
rect 41424 6441 41458 6455
rect 41424 6369 41458 6387
rect 41424 6284 41458 6319
rect 41682 8257 41716 8292
rect 41682 8189 41716 8207
rect 41682 8121 41716 8135
rect 41682 8053 41716 8063
rect 41682 7985 41716 7991
rect 41682 7917 41716 7919
rect 41682 7881 41716 7883
rect 41682 7809 41716 7815
rect 41682 7737 41716 7747
rect 41682 7665 41716 7679
rect 41682 7593 41716 7611
rect 41682 7521 41716 7543
rect 41682 7449 41716 7475
rect 41682 7377 41716 7407
rect 41682 7305 41716 7339
rect 41682 7237 41716 7271
rect 41682 7169 41716 7199
rect 41682 7101 41716 7127
rect 41682 7033 41716 7055
rect 41682 6965 41716 6983
rect 41682 6897 41716 6911
rect 41682 6829 41716 6839
rect 41682 6761 41716 6767
rect 41682 6693 41716 6695
rect 41682 6657 41716 6659
rect 41682 6585 41716 6591
rect 41682 6513 41716 6523
rect 41682 6441 41716 6455
rect 41682 6369 41716 6387
rect 41682 6284 41716 6319
rect 41940 8257 41974 8292
rect 41940 8189 41974 8207
rect 41940 8121 41974 8135
rect 41940 8053 41974 8063
rect 41940 7985 41974 7991
rect 41940 7917 41974 7919
rect 41940 7881 41974 7883
rect 41940 7809 41974 7815
rect 41940 7737 41974 7747
rect 41940 7665 41974 7679
rect 41940 7593 41974 7611
rect 41940 7521 41974 7543
rect 41940 7449 41974 7475
rect 41940 7377 41974 7407
rect 41940 7305 41974 7339
rect 41940 7237 41974 7271
rect 41940 7169 41974 7199
rect 41940 7101 41974 7127
rect 41940 7033 41974 7055
rect 41940 6965 41974 6983
rect 41940 6897 41974 6911
rect 41940 6829 41974 6839
rect 41940 6761 41974 6767
rect 41940 6693 41974 6695
rect 41940 6657 41974 6659
rect 41940 6585 41974 6591
rect 41940 6513 41974 6523
rect 41940 6441 41974 6455
rect 41940 6369 41974 6387
rect 41940 6284 41974 6319
rect 42122 8274 42136 8308
rect 42170 8274 42184 8308
rect 42122 8240 42184 8274
rect 42122 8206 42136 8240
rect 42170 8206 42184 8240
rect 42122 8172 42184 8206
rect 42122 8138 42136 8172
rect 42170 8138 42184 8172
rect 42122 8104 42184 8138
rect 42122 8070 42136 8104
rect 42170 8070 42184 8104
rect 42122 8036 42184 8070
rect 42122 8002 42136 8036
rect 42170 8002 42184 8036
rect 42122 7968 42184 8002
rect 42122 7934 42136 7968
rect 42170 7934 42184 7968
rect 42122 7900 42184 7934
rect 42122 7866 42136 7900
rect 42170 7866 42184 7900
rect 42122 7832 42184 7866
rect 42122 7798 42136 7832
rect 42170 7798 42184 7832
rect 42122 7764 42184 7798
rect 42122 7730 42136 7764
rect 42170 7730 42184 7764
rect 42122 7696 42184 7730
rect 42122 7662 42136 7696
rect 42170 7662 42184 7696
rect 42122 7628 42184 7662
rect 42122 7594 42136 7628
rect 42170 7594 42184 7628
rect 42122 7560 42184 7594
rect 42122 7526 42136 7560
rect 42170 7526 42184 7560
rect 42122 7492 42184 7526
rect 42122 7458 42136 7492
rect 42170 7458 42184 7492
rect 42122 7424 42184 7458
rect 42122 7390 42136 7424
rect 42170 7390 42184 7424
rect 42122 7356 42184 7390
rect 42122 7322 42136 7356
rect 42170 7322 42184 7356
rect 42122 7288 42184 7322
rect 42122 7254 42136 7288
rect 42170 7254 42184 7288
rect 42122 7220 42184 7254
rect 42122 7186 42136 7220
rect 42170 7186 42184 7220
rect 42122 7152 42184 7186
rect 42122 7118 42136 7152
rect 42170 7118 42184 7152
rect 42122 7084 42184 7118
rect 42122 7050 42136 7084
rect 42170 7050 42184 7084
rect 42122 7016 42184 7050
rect 42122 6982 42136 7016
rect 42170 6982 42184 7016
rect 42122 6948 42184 6982
rect 42122 6914 42136 6948
rect 42170 6914 42184 6948
rect 42122 6880 42184 6914
rect 42122 6846 42136 6880
rect 42170 6846 42184 6880
rect 42122 6812 42184 6846
rect 42122 6778 42136 6812
rect 42170 6778 42184 6812
rect 42122 6744 42184 6778
rect 42122 6710 42136 6744
rect 42170 6710 42184 6744
rect 42122 6676 42184 6710
rect 42122 6642 42136 6676
rect 42170 6642 42184 6676
rect 42122 6635 42184 6642
rect 42122 6574 42136 6635
rect 42170 6574 42184 6635
rect 42122 6563 42184 6574
rect 42122 6506 42136 6563
rect 42170 6506 42184 6563
rect 42122 6491 42184 6506
rect 42122 6438 42136 6491
rect 42170 6438 42184 6491
rect 42122 6404 42184 6438
rect 42122 6370 42136 6404
rect 42170 6370 42184 6404
rect 42122 6336 42184 6370
rect 42122 6302 42136 6336
rect 42170 6302 42184 6336
rect 37608 6222 37624 6256
rect 37658 6222 37674 6256
rect 42122 6268 42184 6302
rect 37608 6188 37674 6222
rect 37858 6216 37905 6250
rect 37941 6216 37975 6250
rect 38011 6216 38058 6250
rect 38116 6216 38163 6250
rect 38199 6216 38233 6250
rect 38269 6216 38316 6250
rect 38374 6216 38421 6250
rect 38457 6216 38491 6250
rect 38527 6216 38574 6250
rect 38632 6216 38679 6250
rect 38715 6216 38749 6250
rect 38785 6216 38832 6250
rect 38890 6216 38937 6250
rect 38973 6216 39007 6250
rect 39043 6216 39090 6250
rect 39148 6216 39195 6250
rect 39231 6216 39265 6250
rect 39301 6216 39348 6250
rect 39406 6216 39453 6250
rect 39489 6216 39523 6250
rect 39559 6216 39606 6250
rect 39664 6216 39711 6250
rect 39747 6216 39781 6250
rect 39817 6216 39864 6250
rect 39922 6216 39969 6250
rect 40005 6216 40039 6250
rect 40075 6216 40122 6250
rect 40180 6216 40227 6250
rect 40263 6216 40297 6250
rect 40333 6216 40380 6250
rect 40438 6216 40485 6250
rect 40521 6216 40555 6250
rect 40591 6216 40638 6250
rect 40696 6216 40743 6250
rect 40779 6216 40813 6250
rect 40849 6216 40896 6250
rect 40954 6216 41001 6250
rect 41037 6216 41071 6250
rect 41107 6216 41154 6250
rect 41212 6216 41259 6250
rect 41295 6216 41329 6250
rect 41365 6216 41412 6250
rect 41470 6216 41517 6250
rect 41553 6216 41587 6250
rect 41623 6216 41670 6250
rect 41728 6216 41775 6250
rect 41811 6216 41845 6250
rect 41881 6216 41928 6250
rect 42122 6234 42136 6268
rect 42170 6234 42184 6268
rect 37608 6154 37624 6188
rect 37658 6154 37674 6188
rect 37608 6042 37674 6154
rect 42122 6200 42184 6234
rect 42122 6166 42136 6200
rect 42170 6166 42184 6200
rect 42122 6042 42184 6166
rect 37608 6039 42184 6042
rect 27330 5951 27364 5985
rect 27330 5883 27364 5917
rect 27330 5815 27364 5849
rect 27330 5747 27364 5781
rect 37600 6029 42186 6039
rect 37600 5995 37819 6029
rect 37853 5995 37887 6029
rect 37921 5995 37955 6029
rect 37989 5995 38023 6029
rect 38057 5995 38091 6029
rect 38125 5995 38159 6029
rect 38193 5995 38227 6029
rect 38261 5995 38295 6029
rect 38329 5995 38363 6029
rect 38397 5995 38431 6029
rect 38465 5995 38499 6029
rect 38533 5995 38567 6029
rect 38601 5995 38635 6029
rect 38669 5995 38703 6029
rect 38737 5995 38771 6029
rect 38805 5995 38839 6029
rect 38873 5995 38907 6029
rect 38941 5995 38975 6029
rect 39009 5995 39043 6029
rect 39077 5995 39111 6029
rect 39145 5995 39179 6029
rect 39213 5995 39247 6029
rect 39281 5995 39315 6029
rect 39349 5995 39383 6029
rect 39417 5995 39451 6029
rect 39485 5995 39519 6029
rect 39553 5995 39587 6029
rect 39621 5995 39655 6029
rect 39689 5995 39723 6029
rect 39757 5995 39791 6029
rect 39825 5995 39859 6029
rect 39893 5995 39927 6029
rect 39961 5995 39995 6029
rect 40029 5995 40063 6029
rect 40097 5995 40131 6029
rect 40165 5995 40199 6029
rect 40233 5995 40267 6029
rect 40301 5995 40335 6029
rect 40369 5995 40403 6029
rect 40437 5995 40471 6029
rect 40505 5995 40539 6029
rect 40573 5995 40607 6029
rect 40641 5995 40675 6029
rect 40709 5995 40743 6029
rect 40777 5995 40811 6029
rect 40845 5995 40879 6029
rect 40913 5995 40947 6029
rect 40981 5995 41015 6029
rect 41049 5995 41083 6029
rect 41117 5995 41151 6029
rect 41185 5995 41219 6029
rect 41253 5995 41287 6029
rect 41321 5995 41355 6029
rect 41389 5995 41423 6029
rect 41457 5995 41491 6029
rect 41525 5995 41559 6029
rect 41593 5995 41627 6029
rect 41661 5995 41695 6029
rect 41729 5995 41763 6029
rect 41797 5995 41831 6029
rect 41865 5995 41899 6029
rect 41933 5995 41967 6029
rect 42001 5995 42186 6029
rect 37600 5761 42186 5995
rect 27330 5679 27364 5713
rect 27330 5611 27364 5645
rect 27330 5543 27364 5577
rect 27330 5475 27364 5509
rect 27330 5407 27364 5441
rect 27330 5339 27364 5373
rect 27330 5271 27364 5305
rect 27330 5203 27364 5237
rect 27330 5135 27364 5169
rect 27330 5067 27364 5101
rect 27330 4999 27364 5033
rect 27330 4931 27364 4965
rect 37294 4963 42586 5761
rect 27330 4863 27364 4897
rect 27330 4795 27364 4829
rect 27330 4727 27364 4761
rect 27330 4659 27364 4693
rect 27330 4591 27364 4625
rect 27330 4523 27364 4557
rect 27330 4455 27364 4489
rect 27330 4387 27364 4421
rect 27330 4319 27364 4353
rect 27330 4251 27364 4285
rect 27330 4183 27364 4217
rect 27330 4115 27364 4149
rect 27330 4047 27364 4081
rect 27330 3979 27364 4013
rect 27330 3911 27364 3945
rect 27330 3843 27364 3877
rect 27330 3775 27364 3809
rect 27330 3707 27364 3741
rect 27330 3639 27364 3673
rect 27330 3571 27364 3605
rect 26205 3480 26398 3503
rect 22376 3470 24389 3480
rect 24423 3470 24461 3480
rect 24495 3470 26398 3480
rect 22376 3469 26398 3470
rect 26432 3469 26528 3502
rect 22376 3435 26528 3469
rect 22376 3401 26398 3435
rect 26432 3401 26528 3435
rect 22376 3367 26528 3401
rect 22376 3333 26398 3367
rect 26432 3333 26528 3367
rect 22376 3299 26528 3333
rect 22376 3265 26398 3299
rect 26432 3265 26528 3299
rect 22376 3231 26528 3265
rect 22376 3197 26398 3231
rect 26432 3197 26528 3231
rect 22376 3163 26528 3197
rect 22376 3129 26398 3163
rect 26432 3129 26528 3163
rect 22376 3095 26528 3129
rect 22376 3061 26398 3095
rect 26432 3080 26528 3095
rect 27142 3082 27164 3502
rect 27330 3503 27364 3537
rect 27234 3469 27330 3502
rect 27234 3435 27364 3469
rect 27234 3401 27330 3435
rect 27234 3367 27364 3401
rect 27234 3333 27330 3367
rect 27234 3299 27364 3333
rect 27234 3265 27330 3299
rect 27234 3231 27364 3265
rect 27234 3197 27330 3231
rect 27234 3163 27364 3197
rect 27234 3129 27330 3163
rect 27234 3095 27364 3129
rect 27234 3082 27330 3095
rect 26432 3072 26582 3080
rect 22376 3052 26432 3061
rect 26398 2984 26432 3052
rect 27330 2984 27364 3061
rect 26398 2950 26524 2984
rect 26558 2950 26592 2984
rect 26626 2950 26660 2984
rect 26694 2950 26728 2984
rect 26762 2950 26796 2984
rect 26830 2950 26864 2984
rect 26898 2950 26932 2984
rect 26966 2950 27000 2984
rect 27034 2950 27068 2984
rect 27102 2950 27136 2984
rect 27170 2950 27204 2984
rect 27238 2950 27364 2984
rect -7120 -39 -6980 787
rect -5434 -39 -5286 787
rect 38472 1537 40306 4963
rect 38472 711 38612 1537
rect 40158 711 40306 1537
rect 38472 649 40306 711
rect -7120 -101 -5286 -39
<< viali >>
rect -4261 21359 -3579 22185
rect 41331 22109 42013 22935
rect 41520 19037 41770 19215
rect 43604 19093 43710 19199
rect 23273 18794 23297 18828
rect 23297 18794 23307 18828
rect 23345 18794 23365 18828
rect 23365 18794 23379 18828
rect 23417 18794 23433 18828
rect 23433 18794 23451 18828
rect 23489 18794 23501 18828
rect 23501 18794 23523 18828
rect 23561 18794 23569 18828
rect 23569 18794 23595 18828
rect 23633 18794 23637 18828
rect 23637 18794 23667 18828
rect 23705 18794 23739 18828
rect 23777 18794 23807 18828
rect 23807 18794 23811 18828
rect 23849 18794 23875 18828
rect 23875 18794 23883 18828
rect 23921 18794 23943 18828
rect 23943 18794 23955 18828
rect 23993 18794 24011 18828
rect 24011 18794 24027 18828
rect 24065 18794 24079 18828
rect 24079 18794 24099 18828
rect 24137 18794 24147 18828
rect 24147 18794 24171 18828
rect 23176 18706 23210 18732
rect 23176 18698 23210 18706
rect 23176 18638 23210 18660
rect 24234 18706 24268 18732
rect 24234 18698 24268 18706
rect 23176 18626 23210 18638
rect 23176 18570 23210 18588
rect 23176 18554 23210 18570
rect 24234 18638 24268 18660
rect 24234 18626 24268 18638
rect 24234 18570 24268 18588
rect -4072 18287 -3822 18465
rect -1988 18343 -1882 18449
rect 23176 18502 23210 18516
rect 23176 18482 23210 18502
rect 23176 18434 23210 18444
rect 23176 18410 23210 18434
rect 24234 18554 24268 18570
rect 24234 18502 24268 18516
rect 24234 18482 24268 18502
rect 24234 18434 24268 18444
rect 24234 18410 24268 18434
rect 23176 18366 23210 18372
rect 23176 18338 23210 18366
rect 23176 18298 23210 18300
rect 23176 18266 23210 18298
rect -2887 18140 -2885 18174
rect -2885 18140 -2853 18174
rect -2815 18140 -2783 18174
rect -2783 18140 -2781 18174
rect -2629 18140 -2627 18174
rect -2627 18140 -2595 18174
rect -2557 18140 -2525 18174
rect -2525 18140 -2523 18174
rect -2371 18140 -2369 18174
rect -2369 18140 -2337 18174
rect -2299 18140 -2267 18174
rect -2267 18140 -2265 18174
rect -2113 18140 -2111 18174
rect -2111 18140 -2079 18174
rect -2041 18140 -2009 18174
rect -2009 18140 -2007 18174
rect -1855 18140 -1853 18174
rect -1853 18140 -1821 18174
rect -1783 18140 -1751 18174
rect -1751 18140 -1749 18174
rect -1597 18140 -1595 18174
rect -1595 18140 -1563 18174
rect -1525 18140 -1493 18174
rect -1493 18140 -1491 18174
rect -1339 18140 -1337 18174
rect -1337 18140 -1305 18174
rect -1267 18140 -1235 18174
rect -1235 18140 -1233 18174
rect -1081 18140 -1079 18174
rect -1079 18140 -1047 18174
rect -1009 18140 -977 18174
rect -977 18140 -975 18174
rect -823 18140 -821 18174
rect -821 18140 -789 18174
rect -751 18140 -719 18174
rect -719 18140 -717 18174
rect -565 18140 -563 18174
rect -563 18140 -531 18174
rect -493 18140 -461 18174
rect -461 18140 -459 18174
rect -6239 17536 -6205 17541
rect -6167 17536 -6133 17541
rect -6239 17507 -6226 17536
rect -6226 17507 -6205 17536
rect -6167 17507 -6158 17536
rect -6158 17507 -6133 17536
rect -6355 17271 -6353 17305
rect -6353 17271 -6321 17305
rect -6283 17271 -6251 17305
rect -6251 17271 -6249 17305
rect -6097 17271 -6095 17305
rect -6095 17271 -6063 17305
rect -6025 17271 -5993 17305
rect -5993 17271 -5991 17305
rect -6448 17183 -6414 17209
rect -6448 17175 -6414 17183
rect -6448 17115 -6414 17137
rect -6448 17103 -6414 17115
rect -6448 17047 -6414 17065
rect -6448 17031 -6414 17047
rect -6448 16979 -6414 16993
rect -6448 16959 -6414 16979
rect -6448 16911 -6414 16921
rect -6448 16887 -6414 16911
rect -6448 16843 -6414 16849
rect -6448 16815 -6414 16843
rect -6448 16775 -6414 16777
rect -6448 16743 -6414 16775
rect -6448 16673 -6414 16705
rect -6448 16671 -6414 16673
rect -6448 16605 -6414 16633
rect -6448 16599 -6414 16605
rect -6448 16537 -6414 16561
rect -6448 16527 -6414 16537
rect -6448 16469 -6414 16489
rect -6448 16455 -6414 16469
rect -6448 16401 -6414 16417
rect -6448 16383 -6414 16401
rect -6448 16333 -6414 16345
rect -6448 16311 -6414 16333
rect -6448 16265 -6414 16273
rect -6448 16239 -6414 16265
rect -6190 17183 -6156 17209
rect -6190 17175 -6156 17183
rect -6190 17115 -6156 17137
rect -6190 17103 -6156 17115
rect -6190 17047 -6156 17065
rect -6190 17031 -6156 17047
rect -6190 16979 -6156 16993
rect -6190 16959 -6156 16979
rect -6190 16911 -6156 16921
rect -6190 16887 -6156 16911
rect -6190 16843 -6156 16849
rect -6190 16815 -6156 16843
rect -6190 16775 -6156 16777
rect -6190 16743 -6156 16775
rect -6190 16673 -6156 16705
rect -6190 16671 -6156 16673
rect -6190 16605 -6156 16633
rect -6190 16599 -6156 16605
rect -6190 16537 -6156 16561
rect -6190 16527 -6156 16537
rect -6190 16469 -6156 16489
rect -6190 16455 -6156 16469
rect -6190 16401 -6156 16417
rect -6190 16383 -6156 16401
rect -6190 16333 -6156 16345
rect -6190 16311 -6156 16333
rect -6190 16265 -6156 16273
rect -6190 16239 -6156 16265
rect -5932 17183 -5898 17209
rect -5932 17175 -5898 17183
rect -5932 17115 -5898 17137
rect -5932 17103 -5898 17115
rect -5932 17047 -5898 17065
rect -5932 17031 -5898 17047
rect -5932 16979 -5898 16993
rect -5932 16959 -5898 16979
rect -5932 16911 -5898 16921
rect -5932 16887 -5898 16911
rect -5932 16843 -5898 16849
rect -5932 16815 -5898 16843
rect -5932 16775 -5898 16777
rect -5932 16743 -5898 16775
rect -5932 16673 -5898 16705
rect -5932 16671 -5898 16673
rect -5932 16605 -5898 16633
rect -5932 16599 -5898 16605
rect -5932 16537 -5898 16561
rect -5932 16527 -5898 16537
rect -5932 16469 -5898 16489
rect -5932 16455 -5898 16469
rect -5932 16401 -5898 16417
rect -5932 16383 -5898 16401
rect -5932 16333 -5898 16345
rect -5932 16311 -5898 16333
rect -5932 16265 -5898 16273
rect -5932 16239 -5898 16265
rect -6355 16143 -6353 16177
rect -6353 16143 -6321 16177
rect -6283 16143 -6251 16177
rect -6251 16143 -6249 16177
rect -6097 16143 -6095 16177
rect -6095 16143 -6063 16177
rect -6025 16143 -5993 16177
rect -5993 16143 -5991 16177
rect -2980 18028 -2946 18046
rect -2980 18012 -2946 18028
rect -2980 17960 -2946 17974
rect -2980 17940 -2946 17960
rect -2980 17892 -2946 17902
rect -2980 17868 -2946 17892
rect -2980 17824 -2946 17830
rect -2980 17796 -2946 17824
rect -2980 17756 -2946 17758
rect -2980 17724 -2946 17756
rect -2980 17654 -2946 17686
rect -2980 17652 -2946 17654
rect -2980 17586 -2946 17614
rect -2980 17580 -2946 17586
rect -2980 17518 -2946 17542
rect -2980 17508 -2946 17518
rect -2980 17450 -2946 17470
rect -2980 17436 -2946 17450
rect -2980 17382 -2946 17398
rect -2980 17364 -2946 17382
rect -2980 17314 -2946 17326
rect -2980 17292 -2946 17314
rect -2980 17246 -2946 17254
rect -2980 17220 -2946 17246
rect -2980 17178 -2946 17182
rect -2980 17148 -2946 17178
rect -2980 17076 -2946 17110
rect -2980 17008 -2946 17038
rect -2980 17004 -2946 17008
rect -2980 16940 -2946 16966
rect -2980 16932 -2946 16940
rect -2980 16872 -2946 16894
rect -2980 16860 -2946 16872
rect -2980 16804 -2946 16822
rect -2980 16788 -2946 16804
rect -2980 16736 -2946 16750
rect -2980 16716 -2946 16736
rect -2980 16668 -2946 16678
rect -2980 16644 -2946 16668
rect -2980 16600 -2946 16606
rect -2980 16572 -2946 16600
rect -2980 16532 -2946 16534
rect -2980 16500 -2946 16532
rect -2980 16430 -2946 16462
rect -2980 16428 -2946 16430
rect -2980 16362 -2946 16390
rect -2980 16356 -2946 16362
rect -2980 16294 -2946 16318
rect -2980 16284 -2946 16294
rect -2980 16226 -2946 16246
rect -2980 16212 -2946 16226
rect -2980 16158 -2946 16174
rect -2980 16140 -2946 16158
rect -2722 18028 -2688 18046
rect -2722 18012 -2688 18028
rect -2722 17960 -2688 17974
rect -2722 17940 -2688 17960
rect -2722 17892 -2688 17902
rect -2722 17868 -2688 17892
rect -2722 17824 -2688 17830
rect -2722 17796 -2688 17824
rect -2722 17756 -2688 17758
rect -2722 17724 -2688 17756
rect -2722 17654 -2688 17686
rect -2722 17652 -2688 17654
rect -2722 17586 -2688 17614
rect -2722 17580 -2688 17586
rect -2722 17518 -2688 17542
rect -2722 17508 -2688 17518
rect -2722 17450 -2688 17470
rect -2722 17436 -2688 17450
rect -2722 17382 -2688 17398
rect -2722 17364 -2688 17382
rect -2722 17314 -2688 17326
rect -2722 17292 -2688 17314
rect -2722 17246 -2688 17254
rect -2722 17220 -2688 17246
rect -2722 17178 -2688 17182
rect -2722 17148 -2688 17178
rect -2722 17076 -2688 17110
rect -2722 17008 -2688 17038
rect -2722 17004 -2688 17008
rect -2722 16940 -2688 16966
rect -2722 16932 -2688 16940
rect -2722 16872 -2688 16894
rect -2722 16860 -2688 16872
rect -2722 16804 -2688 16822
rect -2722 16788 -2688 16804
rect -2722 16736 -2688 16750
rect -2722 16716 -2688 16736
rect -2722 16668 -2688 16678
rect -2722 16644 -2688 16668
rect -2722 16600 -2688 16606
rect -2722 16572 -2688 16600
rect -2722 16532 -2688 16534
rect -2722 16500 -2688 16532
rect -2722 16430 -2688 16462
rect -2722 16428 -2688 16430
rect -2722 16362 -2688 16390
rect -2722 16356 -2688 16362
rect -2722 16294 -2688 16318
rect -2722 16284 -2688 16294
rect -2722 16226 -2688 16246
rect -2722 16212 -2688 16226
rect -2722 16158 -2688 16174
rect -2722 16140 -2688 16158
rect -2464 18028 -2430 18046
rect -2464 18012 -2430 18028
rect -2464 17960 -2430 17974
rect -2464 17940 -2430 17960
rect -2464 17892 -2430 17902
rect -2464 17868 -2430 17892
rect -2464 17824 -2430 17830
rect -2464 17796 -2430 17824
rect -2464 17756 -2430 17758
rect -2464 17724 -2430 17756
rect -2464 17654 -2430 17686
rect -2464 17652 -2430 17654
rect -2464 17586 -2430 17614
rect -2464 17580 -2430 17586
rect -2464 17518 -2430 17542
rect -2464 17508 -2430 17518
rect -2464 17450 -2430 17470
rect -2464 17436 -2430 17450
rect -2464 17382 -2430 17398
rect -2464 17364 -2430 17382
rect -2464 17314 -2430 17326
rect -2464 17292 -2430 17314
rect -2464 17246 -2430 17254
rect -2464 17220 -2430 17246
rect -2464 17178 -2430 17182
rect -2464 17148 -2430 17178
rect -2464 17076 -2430 17110
rect -2464 17008 -2430 17038
rect -2464 17004 -2430 17008
rect -2464 16940 -2430 16966
rect -2464 16932 -2430 16940
rect -2464 16872 -2430 16894
rect -2464 16860 -2430 16872
rect -2464 16804 -2430 16822
rect -2464 16788 -2430 16804
rect -2464 16736 -2430 16750
rect -2464 16716 -2430 16736
rect -2464 16668 -2430 16678
rect -2464 16644 -2430 16668
rect -2464 16600 -2430 16606
rect -2464 16572 -2430 16600
rect -2464 16532 -2430 16534
rect -2464 16500 -2430 16532
rect -2464 16430 -2430 16462
rect -2464 16428 -2430 16430
rect -2464 16362 -2430 16390
rect -2464 16356 -2430 16362
rect -2464 16294 -2430 16318
rect -2464 16284 -2430 16294
rect -2464 16226 -2430 16246
rect -2464 16212 -2430 16226
rect -2464 16158 -2430 16174
rect -2464 16140 -2430 16158
rect -2206 18028 -2172 18046
rect -2206 18012 -2172 18028
rect -2206 17960 -2172 17974
rect -2206 17940 -2172 17960
rect -2206 17892 -2172 17902
rect -2206 17868 -2172 17892
rect -2206 17824 -2172 17830
rect -2206 17796 -2172 17824
rect -2206 17756 -2172 17758
rect -2206 17724 -2172 17756
rect -2206 17654 -2172 17686
rect -2206 17652 -2172 17654
rect -2206 17586 -2172 17614
rect -2206 17580 -2172 17586
rect -2206 17518 -2172 17542
rect -2206 17508 -2172 17518
rect -2206 17450 -2172 17470
rect -2206 17436 -2172 17450
rect -2206 17382 -2172 17398
rect -2206 17364 -2172 17382
rect -2206 17314 -2172 17326
rect -2206 17292 -2172 17314
rect -2206 17246 -2172 17254
rect -2206 17220 -2172 17246
rect -2206 17178 -2172 17182
rect -2206 17148 -2172 17178
rect -2206 17076 -2172 17110
rect -2206 17008 -2172 17038
rect -2206 17004 -2172 17008
rect -2206 16940 -2172 16966
rect -2206 16932 -2172 16940
rect -2206 16872 -2172 16894
rect -2206 16860 -2172 16872
rect -2206 16804 -2172 16822
rect -2206 16788 -2172 16804
rect -2206 16736 -2172 16750
rect -2206 16716 -2172 16736
rect -2206 16668 -2172 16678
rect -2206 16644 -2172 16668
rect -2206 16600 -2172 16606
rect -2206 16572 -2172 16600
rect -2206 16532 -2172 16534
rect -2206 16500 -2172 16532
rect -2206 16430 -2172 16462
rect -2206 16428 -2172 16430
rect -2206 16362 -2172 16390
rect -2206 16356 -2172 16362
rect -2206 16294 -2172 16318
rect -2206 16284 -2172 16294
rect -2206 16226 -2172 16246
rect -2206 16212 -2172 16226
rect -2206 16158 -2172 16174
rect -2206 16140 -2172 16158
rect -1948 18028 -1914 18046
rect -1948 18012 -1914 18028
rect -1948 17960 -1914 17974
rect -1948 17940 -1914 17960
rect -1948 17892 -1914 17902
rect -1948 17868 -1914 17892
rect -1948 17824 -1914 17830
rect -1948 17796 -1914 17824
rect -1948 17756 -1914 17758
rect -1948 17724 -1914 17756
rect -1948 17654 -1914 17686
rect -1948 17652 -1914 17654
rect -1948 17586 -1914 17614
rect -1948 17580 -1914 17586
rect -1948 17518 -1914 17542
rect -1948 17508 -1914 17518
rect -1948 17450 -1914 17470
rect -1948 17436 -1914 17450
rect -1948 17382 -1914 17398
rect -1948 17364 -1914 17382
rect -1948 17314 -1914 17326
rect -1948 17292 -1914 17314
rect -1948 17246 -1914 17254
rect -1948 17220 -1914 17246
rect -1948 17178 -1914 17182
rect -1948 17148 -1914 17178
rect -1948 17076 -1914 17110
rect -1948 17008 -1914 17038
rect -1948 17004 -1914 17008
rect -1948 16940 -1914 16966
rect -1948 16932 -1914 16940
rect -1948 16872 -1914 16894
rect -1948 16860 -1914 16872
rect -1948 16804 -1914 16822
rect -1948 16788 -1914 16804
rect -1948 16736 -1914 16750
rect -1948 16716 -1914 16736
rect -1948 16668 -1914 16678
rect -1948 16644 -1914 16668
rect -1948 16600 -1914 16606
rect -1948 16572 -1914 16600
rect -1948 16532 -1914 16534
rect -1948 16500 -1914 16532
rect -1948 16430 -1914 16462
rect -1948 16428 -1914 16430
rect -1948 16362 -1914 16390
rect -1948 16356 -1914 16362
rect -1948 16294 -1914 16318
rect -1948 16284 -1914 16294
rect -1948 16226 -1914 16246
rect -1948 16212 -1914 16226
rect -1948 16158 -1914 16174
rect -1948 16140 -1914 16158
rect -1690 18028 -1656 18046
rect -1690 18012 -1656 18028
rect -1690 17960 -1656 17974
rect -1690 17940 -1656 17960
rect -1690 17892 -1656 17902
rect -1690 17868 -1656 17892
rect -1690 17824 -1656 17830
rect -1690 17796 -1656 17824
rect -1690 17756 -1656 17758
rect -1690 17724 -1656 17756
rect -1690 17654 -1656 17686
rect -1690 17652 -1656 17654
rect -1690 17586 -1656 17614
rect -1690 17580 -1656 17586
rect -1690 17518 -1656 17542
rect -1690 17508 -1656 17518
rect -1690 17450 -1656 17470
rect -1690 17436 -1656 17450
rect -1690 17382 -1656 17398
rect -1690 17364 -1656 17382
rect -1690 17314 -1656 17326
rect -1690 17292 -1656 17314
rect -1690 17246 -1656 17254
rect -1690 17220 -1656 17246
rect -1690 17178 -1656 17182
rect -1690 17148 -1656 17178
rect -1690 17076 -1656 17110
rect -1690 17008 -1656 17038
rect -1690 17004 -1656 17008
rect -1690 16940 -1656 16966
rect -1690 16932 -1656 16940
rect -1690 16872 -1656 16894
rect -1690 16860 -1656 16872
rect -1690 16804 -1656 16822
rect -1690 16788 -1656 16804
rect -1690 16736 -1656 16750
rect -1690 16716 -1656 16736
rect -1690 16668 -1656 16678
rect -1690 16644 -1656 16668
rect -1690 16600 -1656 16606
rect -1690 16572 -1656 16600
rect -1690 16532 -1656 16534
rect -1690 16500 -1656 16532
rect -1690 16430 -1656 16462
rect -1690 16428 -1656 16430
rect -1690 16362 -1656 16390
rect -1690 16356 -1656 16362
rect -1690 16294 -1656 16318
rect -1690 16284 -1656 16294
rect -1690 16226 -1656 16246
rect -1690 16212 -1656 16226
rect -1690 16158 -1656 16174
rect -1690 16140 -1656 16158
rect -1432 18028 -1398 18046
rect -1432 18012 -1398 18028
rect -1432 17960 -1398 17974
rect -1432 17940 -1398 17960
rect -1432 17892 -1398 17902
rect -1432 17868 -1398 17892
rect -1432 17824 -1398 17830
rect -1432 17796 -1398 17824
rect -1432 17756 -1398 17758
rect -1432 17724 -1398 17756
rect -1432 17654 -1398 17686
rect -1432 17652 -1398 17654
rect -1432 17586 -1398 17614
rect -1432 17580 -1398 17586
rect -1432 17518 -1398 17542
rect -1432 17508 -1398 17518
rect -1432 17450 -1398 17470
rect -1432 17436 -1398 17450
rect -1432 17382 -1398 17398
rect -1432 17364 -1398 17382
rect -1432 17314 -1398 17326
rect -1432 17292 -1398 17314
rect -1432 17246 -1398 17254
rect -1432 17220 -1398 17246
rect -1432 17178 -1398 17182
rect -1432 17148 -1398 17178
rect -1432 17076 -1398 17110
rect -1432 17008 -1398 17038
rect -1432 17004 -1398 17008
rect -1432 16940 -1398 16966
rect -1432 16932 -1398 16940
rect -1432 16872 -1398 16894
rect -1432 16860 -1398 16872
rect -1432 16804 -1398 16822
rect -1432 16788 -1398 16804
rect -1432 16736 -1398 16750
rect -1432 16716 -1398 16736
rect -1432 16668 -1398 16678
rect -1432 16644 -1398 16668
rect -1432 16600 -1398 16606
rect -1432 16572 -1398 16600
rect -1432 16532 -1398 16534
rect -1432 16500 -1398 16532
rect -1432 16430 -1398 16462
rect -1432 16428 -1398 16430
rect -1432 16362 -1398 16390
rect -1432 16356 -1398 16362
rect -1432 16294 -1398 16318
rect -1432 16284 -1398 16294
rect -1432 16226 -1398 16246
rect -1432 16212 -1398 16226
rect -1432 16158 -1398 16174
rect -1432 16140 -1398 16158
rect -1174 18028 -1140 18046
rect -1174 18012 -1140 18028
rect -1174 17960 -1140 17974
rect -1174 17940 -1140 17960
rect -1174 17892 -1140 17902
rect -1174 17868 -1140 17892
rect -1174 17824 -1140 17830
rect -1174 17796 -1140 17824
rect -1174 17756 -1140 17758
rect -1174 17724 -1140 17756
rect -1174 17654 -1140 17686
rect -1174 17652 -1140 17654
rect -1174 17586 -1140 17614
rect -1174 17580 -1140 17586
rect -1174 17518 -1140 17542
rect -1174 17508 -1140 17518
rect -1174 17450 -1140 17470
rect -1174 17436 -1140 17450
rect -1174 17382 -1140 17398
rect -1174 17364 -1140 17382
rect -1174 17314 -1140 17326
rect -1174 17292 -1140 17314
rect -1174 17246 -1140 17254
rect -1174 17220 -1140 17246
rect -1174 17178 -1140 17182
rect -1174 17148 -1140 17178
rect -1174 17076 -1140 17110
rect -1174 17008 -1140 17038
rect -1174 17004 -1140 17008
rect -1174 16940 -1140 16966
rect -1174 16932 -1140 16940
rect -1174 16872 -1140 16894
rect -1174 16860 -1140 16872
rect -1174 16804 -1140 16822
rect -1174 16788 -1140 16804
rect -1174 16736 -1140 16750
rect -1174 16716 -1140 16736
rect -1174 16668 -1140 16678
rect -1174 16644 -1140 16668
rect -1174 16600 -1140 16606
rect -1174 16572 -1140 16600
rect -1174 16532 -1140 16534
rect -1174 16500 -1140 16532
rect -1174 16430 -1140 16462
rect -1174 16428 -1140 16430
rect -1174 16362 -1140 16390
rect -1174 16356 -1140 16362
rect -1174 16294 -1140 16318
rect -1174 16284 -1140 16294
rect -1174 16226 -1140 16246
rect -1174 16212 -1140 16226
rect -1174 16158 -1140 16174
rect -1174 16140 -1140 16158
rect -916 18028 -882 18046
rect -916 18012 -882 18028
rect -916 17960 -882 17974
rect -916 17940 -882 17960
rect -916 17892 -882 17902
rect -916 17868 -882 17892
rect -916 17824 -882 17830
rect -916 17796 -882 17824
rect -916 17756 -882 17758
rect -916 17724 -882 17756
rect -916 17654 -882 17686
rect -916 17652 -882 17654
rect -916 17586 -882 17614
rect -916 17580 -882 17586
rect -916 17518 -882 17542
rect -916 17508 -882 17518
rect -916 17450 -882 17470
rect -916 17436 -882 17450
rect -916 17382 -882 17398
rect -916 17364 -882 17382
rect -916 17314 -882 17326
rect -916 17292 -882 17314
rect -916 17246 -882 17254
rect -916 17220 -882 17246
rect -916 17178 -882 17182
rect -916 17148 -882 17178
rect -916 17076 -882 17110
rect -916 17008 -882 17038
rect -916 17004 -882 17008
rect -916 16940 -882 16966
rect -916 16932 -882 16940
rect -916 16872 -882 16894
rect -916 16860 -882 16872
rect -916 16804 -882 16822
rect -916 16788 -882 16804
rect -916 16736 -882 16750
rect -916 16716 -882 16736
rect -916 16668 -882 16678
rect -916 16644 -882 16668
rect -916 16600 -882 16606
rect -916 16572 -882 16600
rect -916 16532 -882 16534
rect -916 16500 -882 16532
rect -916 16430 -882 16462
rect -916 16428 -882 16430
rect -916 16362 -882 16390
rect -916 16356 -882 16362
rect -916 16294 -882 16318
rect -916 16284 -882 16294
rect -916 16226 -882 16246
rect -916 16212 -882 16226
rect -916 16158 -882 16174
rect -916 16140 -882 16158
rect -658 18028 -624 18046
rect -658 18012 -624 18028
rect -658 17960 -624 17974
rect -658 17940 -624 17960
rect -658 17892 -624 17902
rect -658 17868 -624 17892
rect -658 17824 -624 17830
rect -658 17796 -624 17824
rect -658 17756 -624 17758
rect -658 17724 -624 17756
rect -658 17654 -624 17686
rect -658 17652 -624 17654
rect -658 17586 -624 17614
rect -658 17580 -624 17586
rect -658 17518 -624 17542
rect -658 17508 -624 17518
rect -658 17450 -624 17470
rect -658 17436 -624 17450
rect -658 17382 -624 17398
rect -658 17364 -624 17382
rect -658 17314 -624 17326
rect -658 17292 -624 17314
rect -658 17246 -624 17254
rect -658 17220 -624 17246
rect -658 17178 -624 17182
rect -658 17148 -624 17178
rect -658 17076 -624 17110
rect -658 17008 -624 17038
rect -658 17004 -624 17008
rect -658 16940 -624 16966
rect -658 16932 -624 16940
rect -658 16872 -624 16894
rect -658 16860 -624 16872
rect -658 16804 -624 16822
rect -658 16788 -624 16804
rect -658 16736 -624 16750
rect -658 16716 -624 16736
rect -658 16668 -624 16678
rect -658 16644 -624 16668
rect -658 16600 -624 16606
rect -658 16572 -624 16600
rect -658 16532 -624 16534
rect -658 16500 -624 16532
rect -658 16430 -624 16462
rect -658 16428 -624 16430
rect -658 16362 -624 16390
rect -658 16356 -624 16362
rect -658 16294 -624 16318
rect -658 16284 -624 16294
rect -658 16226 -624 16246
rect -658 16212 -624 16226
rect -658 16158 -624 16174
rect -658 16140 -624 16158
rect -400 18028 -366 18046
rect -400 18012 -366 18028
rect -400 17960 -366 17974
rect -400 17940 -366 17960
rect -400 17892 -366 17902
rect -400 17868 -366 17892
rect -400 17824 -366 17830
rect -400 17796 -366 17824
rect -400 17756 -366 17758
rect -400 17724 -366 17756
rect -400 17654 -366 17686
rect -400 17652 -366 17654
rect -400 17586 -366 17614
rect -400 17580 -366 17586
rect -400 17518 -366 17542
rect -400 17508 -366 17518
rect -400 17450 -366 17470
rect -400 17436 -366 17450
rect -400 17382 -366 17398
rect -400 17364 -366 17382
rect -400 17314 -366 17326
rect -400 17292 -366 17314
rect -400 17246 -366 17254
rect -400 17220 -366 17246
rect -400 17178 -366 17182
rect -400 17148 -366 17178
rect -400 17076 -366 17110
rect -400 17008 -366 17038
rect -400 17004 -366 17008
rect -400 16940 -366 16966
rect -400 16932 -366 16940
rect -400 16872 -366 16894
rect -400 16860 -366 16872
rect -400 16804 -366 16822
rect -400 16788 -366 16804
rect -400 16736 -366 16750
rect -400 16716 -366 16736
rect -400 16668 -366 16678
rect -400 16644 -366 16668
rect -400 16600 -366 16606
rect -400 16572 -366 16600
rect -400 16532 -366 16534
rect -400 16500 -366 16532
rect -400 16430 -366 16462
rect -400 16428 -366 16430
rect -400 16362 -366 16390
rect -400 16356 -366 16362
rect -400 16294 -366 16318
rect -400 16284 -366 16294
rect -400 16226 -366 16246
rect -400 16212 -366 16226
rect -400 16158 -366 16174
rect -400 16140 -366 16158
rect 23176 18196 23210 18228
rect 23176 18194 23210 18196
rect 23176 18128 23210 18156
rect 23176 18122 23210 18128
rect 23176 18060 23210 18084
rect 23176 18050 23210 18060
rect 24234 18366 24268 18372
rect 24234 18338 24268 18366
rect 24234 18298 24268 18300
rect 24234 18266 24268 18298
rect 24234 18196 24268 18228
rect 24234 18194 24268 18196
rect 24234 18128 24268 18156
rect 24234 18122 24268 18128
rect 24234 18060 24268 18084
rect 24234 18050 24268 18060
rect 23176 17992 23210 18012
rect 23176 17978 23210 17992
rect 23176 17924 23210 17940
rect 23176 17906 23210 17924
rect 23176 17856 23210 17868
rect 23176 17834 23210 17856
rect 23176 17788 23210 17796
rect 23176 17762 23210 17788
rect 24234 17992 24268 18012
rect 24234 17978 24268 17992
rect 24234 17924 24268 17940
rect 24234 17906 24268 17924
rect 24234 17856 24268 17868
rect 24234 17834 24268 17856
rect 24234 17788 24268 17796
rect 24234 17762 24268 17788
rect 24789 18794 24813 18828
rect 24813 18794 24823 18828
rect 24861 18794 24881 18828
rect 24881 18794 24895 18828
rect 24933 18794 24949 18828
rect 24949 18794 24967 18828
rect 25005 18794 25017 18828
rect 25017 18794 25039 18828
rect 25077 18794 25085 18828
rect 25085 18794 25111 18828
rect 25149 18794 25153 18828
rect 25153 18794 25183 18828
rect 25221 18794 25255 18828
rect 25293 18794 25323 18828
rect 25323 18794 25327 18828
rect 25365 18794 25391 18828
rect 25391 18794 25399 18828
rect 25437 18794 25459 18828
rect 25459 18794 25471 18828
rect 25509 18794 25527 18828
rect 25527 18794 25543 18828
rect 25581 18794 25595 18828
rect 25595 18794 25615 18828
rect 25653 18794 25663 18828
rect 25663 18794 25687 18828
rect 25847 18794 25871 18828
rect 25871 18794 25881 18828
rect 25919 18794 25939 18828
rect 25939 18794 25953 18828
rect 25991 18794 26007 18828
rect 26007 18794 26025 18828
rect 26063 18794 26075 18828
rect 26075 18794 26097 18828
rect 26135 18794 26143 18828
rect 26143 18794 26169 18828
rect 26207 18794 26211 18828
rect 26211 18794 26241 18828
rect 26279 18794 26313 18828
rect 26351 18794 26381 18828
rect 26381 18794 26385 18828
rect 26423 18794 26449 18828
rect 26449 18794 26457 18828
rect 26495 18794 26517 18828
rect 26517 18794 26529 18828
rect 26567 18794 26585 18828
rect 26585 18794 26601 18828
rect 26639 18794 26653 18828
rect 26653 18794 26673 18828
rect 26711 18794 26721 18828
rect 26721 18794 26745 18828
rect 26905 18794 26929 18828
rect 26929 18794 26939 18828
rect 26977 18794 26997 18828
rect 26997 18794 27011 18828
rect 27049 18794 27065 18828
rect 27065 18794 27083 18828
rect 27121 18794 27133 18828
rect 27133 18794 27155 18828
rect 27193 18794 27201 18828
rect 27201 18794 27227 18828
rect 27265 18794 27269 18828
rect 27269 18794 27299 18828
rect 27337 18794 27371 18828
rect 27409 18794 27439 18828
rect 27439 18794 27443 18828
rect 27481 18794 27507 18828
rect 27507 18794 27515 18828
rect 27553 18794 27575 18828
rect 27575 18794 27587 18828
rect 27625 18794 27643 18828
rect 27643 18794 27659 18828
rect 27697 18794 27711 18828
rect 27711 18794 27731 18828
rect 27769 18794 27779 18828
rect 27779 18794 27803 18828
rect 24692 18712 24726 18720
rect 24692 18686 24726 18712
rect 24692 18644 24726 18648
rect 24692 18614 24726 18644
rect 24692 18542 24726 18576
rect 25750 18712 25784 18720
rect 25750 18686 25784 18712
rect 25750 18644 25784 18648
rect 25750 18614 25784 18644
rect 24692 18474 24726 18504
rect 24692 18470 24726 18474
rect 24692 18406 24726 18432
rect 24692 18398 24726 18406
rect 23273 17666 23297 17700
rect 23297 17666 23307 17700
rect 23345 17666 23365 17700
rect 23365 17666 23379 17700
rect 23417 17666 23433 17700
rect 23433 17666 23451 17700
rect 23489 17666 23501 17700
rect 23501 17666 23523 17700
rect 23561 17666 23569 17700
rect 23569 17666 23595 17700
rect 23633 17666 23637 17700
rect 23637 17666 23667 17700
rect 23705 17666 23739 17700
rect 23777 17666 23807 17700
rect 23807 17666 23811 17700
rect 23849 17666 23875 17700
rect 23875 17666 23883 17700
rect 23921 17666 23943 17700
rect 23943 17666 23955 17700
rect 23993 17666 24011 17700
rect 24011 17666 24027 17700
rect 24065 17666 24079 17700
rect 24079 17666 24099 17700
rect 24137 17666 24147 17700
rect 24147 17666 24171 17700
rect -2887 16012 -2885 16046
rect -2885 16012 -2853 16046
rect -2815 16012 -2783 16046
rect -2783 16012 -2781 16046
rect -2629 16012 -2627 16046
rect -2627 16012 -2595 16046
rect -2557 16012 -2525 16046
rect -2525 16012 -2523 16046
rect -2371 16012 -2369 16046
rect -2369 16012 -2337 16046
rect -2299 16012 -2267 16046
rect -2267 16012 -2265 16046
rect -2113 16012 -2111 16046
rect -2111 16012 -2079 16046
rect -2041 16012 -2009 16046
rect -2009 16012 -2007 16046
rect -1855 16012 -1853 16046
rect -1853 16012 -1821 16046
rect -1783 16012 -1751 16046
rect -1751 16012 -1749 16046
rect -1597 16012 -1595 16046
rect -1595 16012 -1563 16046
rect -1525 16012 -1493 16046
rect -1493 16012 -1491 16046
rect -1339 16012 -1337 16046
rect -1337 16012 -1305 16046
rect -1267 16012 -1235 16046
rect -1235 16012 -1233 16046
rect -1081 16012 -1079 16046
rect -1079 16012 -1047 16046
rect -1009 16012 -977 16046
rect -977 16012 -975 16046
rect -823 16012 -821 16046
rect -821 16012 -789 16046
rect -751 16012 -719 16046
rect -719 16012 -717 16046
rect -565 16012 -563 16046
rect -563 16012 -531 16046
rect -493 16012 -461 16046
rect -461 16012 -459 16046
rect -7075 15057 -6825 15163
rect -6059 15056 -5737 15162
rect -5006 15137 -4972 15171
rect -5006 15065 -4972 15099
rect -7459 14770 -7425 14788
rect -7459 14754 -7425 14770
rect -7459 14702 -7425 14716
rect -7459 14682 -7425 14702
rect -7459 14634 -7425 14644
rect -7459 14610 -7425 14634
rect -7459 14566 -7425 14572
rect -7459 14538 -7425 14566
rect -7459 14498 -7425 14500
rect -7459 14466 -7425 14498
rect -7459 14396 -7425 14428
rect -7459 14394 -7425 14396
rect -7459 14328 -7425 14356
rect -7459 14322 -7425 14328
rect -7459 14260 -7425 14284
rect -7459 14250 -7425 14260
rect -7459 14192 -7425 14212
rect -7459 14178 -7425 14192
rect -7459 14124 -7425 14140
rect -7459 14106 -7425 14124
rect -7459 14056 -7425 14068
rect -7459 14034 -7425 14056
rect -7459 13988 -7425 13996
rect -7459 13962 -7425 13988
rect -7459 13920 -7425 13924
rect -7459 13890 -7425 13920
rect -7459 13818 -7425 13852
rect -7459 13750 -7425 13780
rect -7459 13746 -7425 13750
rect -7459 13682 -7425 13708
rect -7459 13674 -7425 13682
rect -7459 13614 -7425 13636
rect -7459 13602 -7425 13614
rect -7459 13546 -7425 13564
rect -7459 13530 -7425 13546
rect -7459 13478 -7425 13492
rect -7459 13458 -7425 13478
rect -7459 13410 -7425 13420
rect -7459 13386 -7425 13410
rect -7459 13342 -7425 13348
rect -7459 13314 -7425 13342
rect -7459 13274 -7425 13276
rect -7459 13242 -7425 13274
rect -7459 13172 -7425 13204
rect -7459 13170 -7425 13172
rect -7459 13104 -7425 13132
rect -7459 13098 -7425 13104
rect -7459 13036 -7425 13060
rect -7459 13026 -7425 13036
rect -7459 12968 -7425 12988
rect -7459 12954 -7425 12968
rect -7459 12900 -7425 12916
rect -7459 12882 -7425 12900
rect -7201 14770 -7167 14788
rect -7201 14754 -7167 14770
rect -7201 14702 -7167 14716
rect -7201 14682 -7167 14702
rect -7201 14634 -7167 14644
rect -7201 14610 -7167 14634
rect -7201 14566 -7167 14572
rect -7201 14538 -7167 14566
rect -7201 14498 -7167 14500
rect -7201 14466 -7167 14498
rect -7201 14396 -7167 14428
rect -7201 14394 -7167 14396
rect -7201 14328 -7167 14356
rect -7201 14322 -7167 14328
rect -7201 14260 -7167 14284
rect -7201 14250 -7167 14260
rect -7201 14192 -7167 14212
rect -7201 14178 -7167 14192
rect -7201 14124 -7167 14140
rect -7201 14106 -7167 14124
rect -7201 14056 -7167 14068
rect -7201 14034 -7167 14056
rect -7201 13988 -7167 13996
rect -7201 13962 -7167 13988
rect -7201 13920 -7167 13924
rect -7201 13890 -7167 13920
rect -7201 13818 -7167 13852
rect -7201 13750 -7167 13780
rect -7201 13746 -7167 13750
rect -7201 13682 -7167 13708
rect -7201 13674 -7167 13682
rect -7201 13614 -7167 13636
rect -7201 13602 -7167 13614
rect -7201 13546 -7167 13564
rect -7201 13530 -7167 13546
rect -7201 13478 -7167 13492
rect -7201 13458 -7167 13478
rect -7201 13410 -7167 13420
rect -7201 13386 -7167 13410
rect -7201 13342 -7167 13348
rect -7201 13314 -7167 13342
rect -7201 13274 -7167 13276
rect -7201 13242 -7167 13274
rect -7201 13172 -7167 13204
rect -7201 13170 -7167 13172
rect -7201 13104 -7167 13132
rect -7201 13098 -7167 13104
rect -7201 13036 -7167 13060
rect -7201 13026 -7167 13036
rect -7201 12968 -7167 12988
rect -7201 12954 -7167 12968
rect -7201 12900 -7167 12916
rect -7201 12882 -7167 12900
rect -6943 14770 -6909 14788
rect -6943 14754 -6909 14770
rect -6943 14702 -6909 14716
rect -6943 14682 -6909 14702
rect -6943 14634 -6909 14644
rect -6943 14610 -6909 14634
rect -6943 14566 -6909 14572
rect -6943 14538 -6909 14566
rect -6943 14498 -6909 14500
rect -6943 14466 -6909 14498
rect -6943 14396 -6909 14428
rect -6943 14394 -6909 14396
rect -6943 14328 -6909 14356
rect -6943 14322 -6909 14328
rect -6943 14260 -6909 14284
rect -6943 14250 -6909 14260
rect -6943 14192 -6909 14212
rect -6943 14178 -6909 14192
rect -6943 14124 -6909 14140
rect -6943 14106 -6909 14124
rect -6943 14056 -6909 14068
rect -6943 14034 -6909 14056
rect -6943 13988 -6909 13996
rect -6943 13962 -6909 13988
rect -6943 13920 -6909 13924
rect -6943 13890 -6909 13920
rect -6943 13818 -6909 13852
rect -6943 13750 -6909 13780
rect -6943 13746 -6909 13750
rect -6943 13682 -6909 13708
rect -6943 13674 -6909 13682
rect -6943 13614 -6909 13636
rect -6943 13602 -6909 13614
rect -6943 13546 -6909 13564
rect -6943 13530 -6909 13546
rect -6943 13478 -6909 13492
rect -6943 13458 -6909 13478
rect -6943 13410 -6909 13420
rect -6943 13386 -6909 13410
rect -6943 13342 -6909 13348
rect -6943 13314 -6909 13342
rect -6943 13274 -6909 13276
rect -6943 13242 -6909 13274
rect -6943 13172 -6909 13204
rect -6943 13170 -6909 13172
rect -6943 13104 -6909 13132
rect -6943 13098 -6909 13104
rect -6943 13036 -6909 13060
rect -6943 13026 -6909 13036
rect -6943 12968 -6909 12988
rect -6943 12954 -6909 12968
rect -6943 12900 -6909 12916
rect -6943 12882 -6909 12900
rect -6685 14770 -6651 14788
rect -6685 14754 -6651 14770
rect -6685 14702 -6651 14716
rect -6685 14682 -6651 14702
rect -6685 14634 -6651 14644
rect -6685 14610 -6651 14634
rect -6685 14566 -6651 14572
rect -6685 14538 -6651 14566
rect -6685 14498 -6651 14500
rect -6685 14466 -6651 14498
rect -6685 14396 -6651 14428
rect -6685 14394 -6651 14396
rect -6685 14328 -6651 14356
rect -6685 14322 -6651 14328
rect -6685 14260 -6651 14284
rect -6685 14250 -6651 14260
rect -6685 14192 -6651 14212
rect -6685 14178 -6651 14192
rect -6685 14124 -6651 14140
rect -6685 14106 -6651 14124
rect -6685 14056 -6651 14068
rect -6685 14034 -6651 14056
rect -6685 13988 -6651 13996
rect -6685 13962 -6651 13988
rect -6685 13920 -6651 13924
rect -6685 13890 -6651 13920
rect -6685 13818 -6651 13852
rect -6685 13750 -6651 13780
rect -6685 13746 -6651 13750
rect -6685 13682 -6651 13708
rect -6685 13674 -6651 13682
rect -6685 13614 -6651 13636
rect -6685 13602 -6651 13614
rect -6685 13546 -6651 13564
rect -6685 13530 -6651 13546
rect -6685 13478 -6651 13492
rect -6685 13458 -6651 13478
rect -6685 13410 -6651 13420
rect -6685 13386 -6651 13410
rect -6685 13342 -6651 13348
rect -6685 13314 -6651 13342
rect -6685 13274 -6651 13276
rect -6685 13242 -6651 13274
rect -6685 13172 -6651 13204
rect -6685 13170 -6651 13172
rect -6685 13104 -6651 13132
rect -6685 13098 -6651 13104
rect -6685 13036 -6651 13060
rect -6685 13026 -6651 13036
rect -6685 12968 -6651 12988
rect -6685 12954 -6651 12968
rect -6685 12900 -6651 12916
rect -6685 12882 -6651 12900
rect -6427 14770 -6393 14788
rect -6427 14754 -6393 14770
rect -6427 14702 -6393 14716
rect -6427 14682 -6393 14702
rect -6427 14634 -6393 14644
rect -6427 14610 -6393 14634
rect -6427 14566 -6393 14572
rect -6427 14538 -6393 14566
rect -6427 14498 -6393 14500
rect -6427 14466 -6393 14498
rect -6427 14396 -6393 14428
rect -6427 14394 -6393 14396
rect -6427 14328 -6393 14356
rect -6427 14322 -6393 14328
rect -6427 14260 -6393 14284
rect -6427 14250 -6393 14260
rect -6427 14192 -6393 14212
rect -6427 14178 -6393 14192
rect -6427 14124 -6393 14140
rect -6427 14106 -6393 14124
rect -6427 14056 -6393 14068
rect -6427 14034 -6393 14056
rect -6427 13988 -6393 13996
rect -6427 13962 -6393 13988
rect -6427 13920 -6393 13924
rect -6427 13890 -6393 13920
rect -6427 13818 -6393 13852
rect -6427 13750 -6393 13780
rect -6427 13746 -6393 13750
rect -6427 13682 -6393 13708
rect -6427 13674 -6393 13682
rect -6427 13614 -6393 13636
rect -6427 13602 -6393 13614
rect -6427 13546 -6393 13564
rect -6427 13530 -6393 13546
rect -6427 13478 -6393 13492
rect -6427 13458 -6393 13478
rect -6427 13410 -6393 13420
rect -6427 13386 -6393 13410
rect -6427 13342 -6393 13348
rect -6427 13314 -6393 13342
rect -6427 13274 -6393 13276
rect -6427 13242 -6393 13274
rect -6427 13172 -6393 13204
rect -6427 13170 -6393 13172
rect -6427 13104 -6393 13132
rect -6427 13098 -6393 13104
rect -6427 13036 -6393 13060
rect -6427 13026 -6393 13036
rect -6427 12968 -6393 12988
rect -6427 12954 -6393 12968
rect -6427 12900 -6393 12916
rect -6427 12882 -6393 12900
rect -6169 14770 -6135 14788
rect -6169 14754 -6135 14770
rect -6169 14702 -6135 14716
rect -6169 14682 -6135 14702
rect -6169 14634 -6135 14644
rect -6169 14610 -6135 14634
rect -6169 14566 -6135 14572
rect -6169 14538 -6135 14566
rect -6169 14498 -6135 14500
rect -6169 14466 -6135 14498
rect -6169 14396 -6135 14428
rect -6169 14394 -6135 14396
rect -6169 14328 -6135 14356
rect -6169 14322 -6135 14328
rect -6169 14260 -6135 14284
rect -6169 14250 -6135 14260
rect -6169 14192 -6135 14212
rect -6169 14178 -6135 14192
rect -6169 14124 -6135 14140
rect -6169 14106 -6135 14124
rect -6169 14056 -6135 14068
rect -6169 14034 -6135 14056
rect -6169 13988 -6135 13996
rect -6169 13962 -6135 13988
rect -6169 13920 -6135 13924
rect -6169 13890 -6135 13920
rect -6169 13818 -6135 13852
rect -6169 13750 -6135 13780
rect -6169 13746 -6135 13750
rect -6169 13682 -6135 13708
rect -6169 13674 -6135 13682
rect -6169 13614 -6135 13636
rect -6169 13602 -6135 13614
rect -6169 13546 -6135 13564
rect -6169 13530 -6135 13546
rect -6169 13478 -6135 13492
rect -6169 13458 -6135 13478
rect -6169 13410 -6135 13420
rect -6169 13386 -6135 13410
rect -6169 13342 -6135 13348
rect -6169 13314 -6135 13342
rect -6169 13274 -6135 13276
rect -6169 13242 -6135 13274
rect -6169 13172 -6135 13204
rect -6169 13170 -6135 13172
rect -6169 13104 -6135 13132
rect -6169 13098 -6135 13104
rect -6169 13036 -6135 13060
rect -6169 13026 -6135 13036
rect -6169 12968 -6135 12988
rect -6169 12954 -6135 12968
rect -6169 12900 -6135 12916
rect -6169 12882 -6135 12900
rect -6840 12724 -6806 12758
rect -6768 12724 -6734 12758
rect -5911 14770 -5877 14788
rect -5911 14754 -5877 14770
rect -5911 14702 -5877 14716
rect -5911 14682 -5877 14702
rect -5911 14634 -5877 14644
rect -5911 14610 -5877 14634
rect -5911 14566 -5877 14572
rect -5911 14538 -5877 14566
rect -5911 14498 -5877 14500
rect -5911 14466 -5877 14498
rect -5911 14396 -5877 14428
rect -5911 14394 -5877 14396
rect -5911 14328 -5877 14356
rect -5911 14322 -5877 14328
rect -5911 14260 -5877 14284
rect -5911 14250 -5877 14260
rect -5911 14192 -5877 14212
rect -5911 14178 -5877 14192
rect -5911 14124 -5877 14140
rect -5911 14106 -5877 14124
rect -5911 14056 -5877 14068
rect -5911 14034 -5877 14056
rect -5911 13988 -5877 13996
rect -5911 13962 -5877 13988
rect -5911 13920 -5877 13924
rect -5911 13890 -5877 13920
rect -5911 13818 -5877 13852
rect -5911 13750 -5877 13780
rect -5911 13746 -5877 13750
rect -5911 13682 -5877 13708
rect -5911 13674 -5877 13682
rect -5911 13614 -5877 13636
rect -5911 13602 -5877 13614
rect -5911 13546 -5877 13564
rect -5911 13530 -5877 13546
rect -5911 13478 -5877 13492
rect -5911 13458 -5877 13478
rect -5911 13410 -5877 13420
rect -5911 13386 -5877 13410
rect -5911 13342 -5877 13348
rect -5911 13314 -5877 13342
rect -5911 13274 -5877 13276
rect -5911 13242 -5877 13274
rect -5911 13172 -5877 13204
rect -5911 13170 -5877 13172
rect -5911 13104 -5877 13132
rect -5911 13098 -5877 13104
rect -5911 13036 -5877 13060
rect -5911 13026 -5877 13036
rect -5911 12968 -5877 12988
rect -5911 12954 -5877 12968
rect -5911 12900 -5877 12916
rect -5911 12882 -5877 12900
rect -5436 14901 -5402 14935
rect -5364 14901 -5330 14935
rect -5292 14901 -5258 14935
rect -5653 14770 -5619 14788
rect -5653 14754 -5619 14770
rect -5653 14702 -5619 14716
rect -5653 14682 -5619 14702
rect -5653 14634 -5619 14644
rect -5653 14610 -5619 14634
rect -5653 14566 -5619 14572
rect -5653 14538 -5619 14566
rect -5653 14498 -5619 14500
rect -5653 14466 -5619 14498
rect -5653 14396 -5619 14428
rect -5653 14394 -5619 14396
rect -5653 14328 -5619 14356
rect -5653 14322 -5619 14328
rect -5653 14260 -5619 14284
rect -5653 14250 -5619 14260
rect -5653 14192 -5619 14212
rect -5653 14178 -5619 14192
rect -5653 14124 -5619 14140
rect -5653 14106 -5619 14124
rect -5653 14056 -5619 14068
rect -5653 14034 -5619 14056
rect -5653 13988 -5619 13996
rect -5653 13962 -5619 13988
rect -5653 13920 -5619 13924
rect -5653 13890 -5619 13920
rect -5653 13818 -5619 13852
rect -5653 13750 -5619 13780
rect -5653 13746 -5619 13750
rect -5653 13682 -5619 13708
rect -5653 13674 -5619 13682
rect -5653 13614 -5619 13636
rect -5653 13602 -5619 13614
rect -5653 13546 -5619 13564
rect -5653 13530 -5619 13546
rect -5653 13478 -5619 13492
rect -5653 13458 -5619 13478
rect -5653 13410 -5619 13420
rect -5653 13386 -5619 13410
rect -5653 13342 -5619 13348
rect -5653 13314 -5619 13342
rect -5653 13274 -5619 13276
rect -5653 13242 -5619 13274
rect -5653 13172 -5619 13204
rect -5653 13170 -5619 13172
rect -5653 13104 -5619 13132
rect -5653 13098 -5619 13104
rect -5653 13036 -5619 13060
rect -5653 13026 -5619 13036
rect -5653 12968 -5619 12988
rect -5653 12954 -5619 12968
rect -5653 12900 -5619 12916
rect -5653 12882 -5619 12900
rect -5395 14770 -5361 14788
rect -5395 14754 -5361 14770
rect -5395 14702 -5361 14716
rect -5395 14682 -5361 14702
rect -5395 14634 -5361 14644
rect -5395 14610 -5361 14634
rect -5395 14566 -5361 14572
rect -5395 14538 -5361 14566
rect -5395 14498 -5361 14500
rect -5395 14466 -5361 14498
rect -5395 14396 -5361 14428
rect -5395 14394 -5361 14396
rect -5395 14328 -5361 14356
rect -5395 14322 -5361 14328
rect -5395 14260 -5361 14284
rect -5395 14250 -5361 14260
rect -5395 14192 -5361 14212
rect -5395 14178 -5361 14192
rect -5395 14124 -5361 14140
rect -5395 14106 -5361 14124
rect -5395 14056 -5361 14068
rect -5395 14034 -5361 14056
rect -5395 13988 -5361 13996
rect -5395 13962 -5361 13988
rect -5395 13920 -5361 13924
rect -5395 13890 -5361 13920
rect -5395 13818 -5361 13852
rect -5395 13750 -5361 13780
rect -5395 13746 -5361 13750
rect -5395 13682 -5361 13708
rect -5395 13674 -5361 13682
rect -5395 13614 -5361 13636
rect -5395 13602 -5361 13614
rect -5395 13546 -5361 13564
rect -5395 13530 -5361 13546
rect -5395 13478 -5361 13492
rect -5395 13458 -5361 13478
rect -5395 13410 -5361 13420
rect -5395 13386 -5361 13410
rect -5395 13342 -5361 13348
rect -5395 13314 -5361 13342
rect -5395 13274 -5361 13276
rect -5395 13242 -5361 13274
rect -5395 13172 -5361 13204
rect -5395 13170 -5361 13172
rect -5395 13104 -5361 13132
rect -5395 13098 -5361 13104
rect -5395 13036 -5361 13060
rect -5395 13026 -5361 13036
rect -5395 12968 -5361 12988
rect -5395 12954 -5361 12968
rect -5395 12900 -5361 12916
rect -5395 12882 -5361 12900
rect -5137 14770 -5103 14788
rect -5137 14754 -5103 14770
rect -5137 14702 -5103 14716
rect -5137 14682 -5103 14702
rect -5137 14634 -5103 14644
rect -5137 14610 -5103 14634
rect -5137 14566 -5103 14572
rect -5137 14538 -5103 14566
rect -5137 14498 -5103 14500
rect -5137 14466 -5103 14498
rect -5137 14396 -5103 14428
rect -5137 14394 -5103 14396
rect -5137 14328 -5103 14356
rect -5137 14322 -5103 14328
rect -5137 14260 -5103 14284
rect -5137 14250 -5103 14260
rect -5137 14192 -5103 14212
rect -5137 14178 -5103 14192
rect -5137 14124 -5103 14140
rect -5137 14106 -5103 14124
rect -5137 14056 -5103 14068
rect -5137 14034 -5103 14056
rect -5137 13988 -5103 13996
rect -5137 13962 -5103 13988
rect -5137 13920 -5103 13924
rect -5137 13890 -5103 13920
rect -5137 13818 -5103 13852
rect -5137 13750 -5103 13780
rect -5137 13746 -5103 13750
rect -5137 13682 -5103 13708
rect -5137 13674 -5103 13682
rect -5137 13614 -5103 13636
rect -5137 13602 -5103 13614
rect -5137 13546 -5103 13564
rect -5137 13530 -5103 13546
rect -5137 13478 -5103 13492
rect -5137 13458 -5103 13478
rect -5137 13410 -5103 13420
rect -5137 13386 -5103 13410
rect -5137 13342 -5103 13348
rect -5137 13314 -5103 13342
rect -5137 13274 -5103 13276
rect -5137 13242 -5103 13274
rect -5137 13172 -5103 13204
rect -5137 13170 -5103 13172
rect -5137 13104 -5103 13132
rect -5137 13098 -5103 13104
rect -5137 13036 -5103 13060
rect -5137 13026 -5103 13036
rect -5137 12968 -5103 12988
rect -5137 12954 -5103 12968
rect -5137 12900 -5103 12916
rect -5137 12882 -5103 12900
rect -4879 14770 -4845 14788
rect -4879 14754 -4845 14770
rect -4879 14702 -4845 14716
rect -4879 14682 -4845 14702
rect -4879 14634 -4845 14644
rect -4879 14610 -4845 14634
rect -4879 14566 -4845 14572
rect -4879 14538 -4845 14566
rect -4879 14498 -4845 14500
rect -4879 14466 -4845 14498
rect -4879 14396 -4845 14428
rect -4879 14394 -4845 14396
rect -4879 14328 -4845 14356
rect -4879 14322 -4845 14328
rect -4879 14260 -4845 14284
rect -4879 14250 -4845 14260
rect -4879 14192 -4845 14212
rect -4879 14178 -4845 14192
rect -4879 14124 -4845 14140
rect -4879 14106 -4845 14124
rect -4879 14056 -4845 14068
rect -4879 14034 -4845 14056
rect -4879 13988 -4845 13996
rect -4879 13962 -4845 13988
rect -4879 13920 -4845 13924
rect -4879 13890 -4845 13920
rect -4879 13818 -4845 13852
rect -4879 13750 -4845 13780
rect -4879 13746 -4845 13750
rect -4879 13682 -4845 13708
rect -4879 13674 -4845 13682
rect -4879 13614 -4845 13636
rect -4879 13602 -4845 13614
rect -4879 13546 -4845 13564
rect -4879 13530 -4845 13546
rect -4879 13478 -4845 13492
rect -4879 13458 -4845 13478
rect -4879 13410 -4845 13420
rect -4879 13386 -4845 13410
rect -4879 13342 -4845 13348
rect -4879 13314 -4845 13342
rect -4879 13274 -4845 13276
rect -4879 13242 -4845 13274
rect -4879 13172 -4845 13204
rect -4879 13170 -4845 13172
rect -4879 13104 -4845 13132
rect -4879 13098 -4845 13104
rect -4879 13036 -4845 13060
rect -4879 13026 -4845 13036
rect -4879 12968 -4845 12988
rect -4879 12954 -4845 12968
rect -4879 12900 -4845 12916
rect -4879 12882 -4845 12900
rect -7339 12518 -7305 12552
rect -7339 12446 -7305 12480
rect -6550 12526 -6516 12560
rect -6550 12454 -6516 12488
rect -6310 12528 -6276 12562
rect -6310 12456 -6276 12490
rect -5531 12523 -5497 12557
rect -5531 12451 -5497 12485
rect -5262 12536 -5228 12570
rect -5262 12464 -5228 12498
rect 10358 15011 11256 17061
rect 23247 17174 23271 17208
rect 23271 17174 23281 17208
rect 23319 17174 23339 17208
rect 23339 17174 23353 17208
rect 23391 17174 23407 17208
rect 23407 17174 23425 17208
rect 23463 17174 23475 17208
rect 23475 17174 23497 17208
rect 23535 17174 23543 17208
rect 23543 17174 23569 17208
rect 23607 17174 23611 17208
rect 23611 17174 23641 17208
rect 23679 17174 23713 17208
rect 23751 17174 23781 17208
rect 23781 17174 23785 17208
rect 23823 17174 23849 17208
rect 23849 17174 23857 17208
rect 23895 17174 23917 17208
rect 23917 17174 23929 17208
rect 23967 17174 23985 17208
rect 23985 17174 24001 17208
rect 24039 17174 24053 17208
rect 24053 17174 24073 17208
rect 24111 17174 24121 17208
rect 24121 17174 24145 17208
rect 23150 17095 23184 17121
rect 23150 17087 23184 17095
rect 23150 17027 23184 17049
rect 23150 17015 23184 17027
rect 24208 17095 24242 17121
rect 24208 17087 24242 17095
rect 24208 17027 24242 17049
rect 24208 17015 24242 17027
rect 23150 16959 23184 16977
rect 23150 16943 23184 16959
rect 23150 16891 23184 16905
rect 23150 16871 23184 16891
rect 24208 16959 24242 16977
rect 24208 16943 24242 16959
rect 24208 16891 24242 16905
rect 24208 16871 24242 16891
rect 23150 16823 23184 16833
rect 23150 16799 23184 16823
rect 23150 16755 23184 16761
rect 23150 16727 23184 16755
rect 23150 16687 23184 16689
rect 23150 16655 23184 16687
rect 23150 16585 23184 16617
rect 23150 16583 23184 16585
rect 23150 16517 23184 16545
rect 24208 16823 24242 16833
rect 24208 16799 24242 16823
rect 24208 16755 24242 16761
rect 24208 16727 24242 16755
rect 25750 18542 25784 18576
rect 25750 18474 25784 18504
rect 25750 18470 25784 18474
rect 25750 18406 25784 18432
rect 25750 18398 25784 18406
rect 24692 18338 24726 18360
rect 24692 18326 24726 18338
rect 24692 18270 24726 18288
rect 24692 18254 24726 18270
rect 24692 18202 24726 18216
rect 24692 18182 24726 18202
rect 24692 18134 24726 18144
rect 24692 18110 24726 18134
rect 24692 18066 24726 18072
rect 24692 18038 24726 18066
rect 24692 17998 24726 18000
rect 24692 17966 24726 17998
rect 24692 17896 24726 17928
rect 24692 17894 24726 17896
rect 24692 17828 24726 17856
rect 24692 17822 24726 17828
rect 24692 17760 24726 17784
rect 24692 17750 24726 17760
rect 24692 17692 24726 17712
rect 24692 17678 24726 17692
rect 24692 17624 24726 17640
rect 24692 17606 24726 17624
rect 24692 17556 24726 17568
rect 24692 17534 24726 17556
rect 24692 17488 24726 17496
rect 24692 17462 24726 17488
rect 24692 17420 24726 17424
rect 24692 17390 24726 17420
rect 24692 17318 24726 17352
rect 24692 17250 24726 17280
rect 24692 17246 24726 17250
rect 24692 17182 24726 17208
rect 24692 17174 24726 17182
rect 25750 18338 25784 18360
rect 25750 18326 25784 18338
rect 25750 18270 25784 18288
rect 25750 18254 25784 18270
rect 25750 18202 25784 18216
rect 25750 18182 25784 18202
rect 25750 18134 25784 18144
rect 25750 18110 25784 18134
rect 25750 18066 25784 18072
rect 25750 18038 25784 18066
rect 25750 17998 25784 18000
rect 25750 17966 25784 17998
rect 25750 17896 25784 17928
rect 25750 17894 25784 17896
rect 25750 17828 25784 17856
rect 25750 17822 25784 17828
rect 25750 17760 25784 17784
rect 25750 17750 25784 17760
rect 25750 17692 25784 17712
rect 25750 17678 25784 17692
rect 25750 17624 25784 17640
rect 25750 17606 25784 17624
rect 25750 17556 25784 17568
rect 25750 17534 25784 17556
rect 25750 17488 25784 17496
rect 25750 17462 25784 17488
rect 25750 17420 25784 17424
rect 25750 17390 25784 17420
rect 25750 17318 25784 17352
rect 25750 17250 25784 17280
rect 25750 17246 25784 17250
rect 25750 17182 25784 17208
rect 25750 17174 25784 17182
rect 26808 18712 26842 18720
rect 26808 18686 26842 18712
rect 26808 18644 26842 18648
rect 26808 18614 26842 18644
rect 26808 18542 26842 18576
rect 26808 18474 26842 18504
rect 26808 18470 26842 18474
rect 26808 18406 26842 18432
rect 26808 18398 26842 18406
rect 26808 18338 26842 18360
rect 26808 18326 26842 18338
rect 26808 18270 26842 18288
rect 26808 18254 26842 18270
rect 26808 18202 26842 18216
rect 26808 18182 26842 18202
rect 26808 18134 26842 18144
rect 26808 18110 26842 18134
rect 26808 18066 26842 18072
rect 26808 18038 26842 18066
rect 26808 17998 26842 18000
rect 26808 17966 26842 17998
rect 26808 17896 26842 17928
rect 26808 17894 26842 17896
rect 26808 17828 26842 17856
rect 26808 17822 26842 17828
rect 26808 17760 26842 17784
rect 26808 17750 26842 17760
rect 26808 17692 26842 17712
rect 26808 17678 26842 17692
rect 26808 17624 26842 17640
rect 26808 17606 26842 17624
rect 26808 17556 26842 17568
rect 26808 17534 26842 17556
rect 26808 17488 26842 17496
rect 26808 17462 26842 17488
rect 26808 17420 26842 17424
rect 26808 17390 26842 17420
rect 26808 17318 26842 17352
rect 26808 17250 26842 17280
rect 26808 17246 26842 17250
rect 26808 17182 26842 17208
rect 26808 17174 26842 17182
rect 27866 18712 27900 18720
rect 27866 18686 27900 18712
rect 27866 18644 27900 18648
rect 27866 18614 27900 18644
rect 27866 18542 27900 18576
rect 27866 18474 27900 18504
rect 27866 18470 27900 18474
rect 27866 18406 27900 18432
rect 27866 18398 27900 18406
rect 27866 18338 27900 18360
rect 27866 18326 27900 18338
rect 27866 18270 27900 18288
rect 27866 18254 27900 18270
rect 27866 18202 27900 18216
rect 27866 18182 27900 18202
rect 27866 18134 27900 18144
rect 27866 18110 27900 18134
rect 27866 18066 27900 18072
rect 27866 18038 27900 18066
rect 27866 17998 27900 18000
rect 27866 17966 27900 17998
rect 27866 17896 27900 17928
rect 27866 17894 27900 17896
rect 27866 17828 27900 17856
rect 27866 17822 27900 17828
rect 27866 17760 27900 17784
rect 27866 17750 27900 17760
rect 27866 17692 27900 17712
rect 27866 17678 27900 17692
rect 27866 17624 27900 17640
rect 27866 17606 27900 17624
rect 27866 17556 27900 17568
rect 27866 17534 27900 17556
rect 27866 17488 27900 17496
rect 27866 17462 27900 17488
rect 27866 17420 27900 17424
rect 27866 17390 27900 17420
rect 27866 17318 27900 17352
rect 27866 17250 27900 17280
rect 27866 17246 27900 17250
rect 27866 17182 27900 17208
rect 27866 17174 27900 17182
rect 42705 18890 42707 18924
rect 42707 18890 42739 18924
rect 42777 18890 42809 18924
rect 42809 18890 42811 18924
rect 42963 18890 42965 18924
rect 42965 18890 42997 18924
rect 43035 18890 43067 18924
rect 43067 18890 43069 18924
rect 43221 18890 43223 18924
rect 43223 18890 43255 18924
rect 43293 18890 43325 18924
rect 43325 18890 43327 18924
rect 43479 18890 43481 18924
rect 43481 18890 43513 18924
rect 43551 18890 43583 18924
rect 43583 18890 43585 18924
rect 43737 18890 43739 18924
rect 43739 18890 43771 18924
rect 43809 18890 43841 18924
rect 43841 18890 43843 18924
rect 43995 18890 43997 18924
rect 43997 18890 44029 18924
rect 44067 18890 44099 18924
rect 44099 18890 44101 18924
rect 44253 18890 44255 18924
rect 44255 18890 44287 18924
rect 44325 18890 44357 18924
rect 44357 18890 44359 18924
rect 44511 18890 44513 18924
rect 44513 18890 44545 18924
rect 44583 18890 44615 18924
rect 44615 18890 44617 18924
rect 44769 18890 44771 18924
rect 44771 18890 44803 18924
rect 44841 18890 44873 18924
rect 44873 18890 44875 18924
rect 45027 18890 45029 18924
rect 45029 18890 45061 18924
rect 45099 18890 45131 18924
rect 45131 18890 45133 18924
rect 39353 18286 39387 18291
rect 39425 18286 39459 18291
rect 39353 18257 39366 18286
rect 39366 18257 39387 18286
rect 39425 18257 39434 18286
rect 39434 18257 39459 18286
rect 24789 17066 24813 17100
rect 24813 17066 24823 17100
rect 24861 17066 24881 17100
rect 24881 17066 24895 17100
rect 24933 17066 24949 17100
rect 24949 17066 24967 17100
rect 25005 17066 25017 17100
rect 25017 17066 25039 17100
rect 25077 17066 25085 17100
rect 25085 17066 25111 17100
rect 25149 17066 25153 17100
rect 25153 17066 25183 17100
rect 25221 17066 25255 17100
rect 25293 17066 25323 17100
rect 25323 17066 25327 17100
rect 25365 17066 25391 17100
rect 25391 17066 25399 17100
rect 25437 17066 25459 17100
rect 25459 17066 25471 17100
rect 25509 17066 25527 17100
rect 25527 17066 25543 17100
rect 25581 17066 25595 17100
rect 25595 17066 25615 17100
rect 25653 17066 25663 17100
rect 25663 17066 25687 17100
rect 25847 17066 25871 17100
rect 25871 17066 25881 17100
rect 25919 17066 25939 17100
rect 25939 17066 25953 17100
rect 25991 17066 26007 17100
rect 26007 17066 26025 17100
rect 26063 17066 26075 17100
rect 26075 17066 26097 17100
rect 26135 17066 26143 17100
rect 26143 17066 26169 17100
rect 26207 17066 26211 17100
rect 26211 17066 26241 17100
rect 26279 17066 26313 17100
rect 26351 17066 26381 17100
rect 26381 17066 26385 17100
rect 26423 17066 26449 17100
rect 26449 17066 26457 17100
rect 26495 17066 26517 17100
rect 26517 17066 26529 17100
rect 26567 17066 26585 17100
rect 26585 17066 26601 17100
rect 26639 17066 26653 17100
rect 26653 17066 26673 17100
rect 26711 17066 26721 17100
rect 26721 17066 26745 17100
rect 26905 17066 26929 17100
rect 26929 17066 26939 17100
rect 26977 17066 26997 17100
rect 26997 17066 27011 17100
rect 27049 17066 27065 17100
rect 27065 17066 27083 17100
rect 27121 17066 27133 17100
rect 27133 17066 27155 17100
rect 27193 17066 27201 17100
rect 27201 17066 27227 17100
rect 27265 17066 27269 17100
rect 27269 17066 27299 17100
rect 27337 17066 27371 17100
rect 27409 17066 27439 17100
rect 27439 17066 27443 17100
rect 27481 17066 27507 17100
rect 27507 17066 27515 17100
rect 27553 17066 27575 17100
rect 27575 17066 27587 17100
rect 27625 17066 27643 17100
rect 27643 17066 27659 17100
rect 27697 17066 27711 17100
rect 27711 17066 27731 17100
rect 27769 17066 27779 17100
rect 27779 17066 27803 17100
rect 39237 18021 39239 18055
rect 39239 18021 39271 18055
rect 39309 18021 39341 18055
rect 39341 18021 39343 18055
rect 39495 18021 39497 18055
rect 39497 18021 39529 18055
rect 39567 18021 39599 18055
rect 39599 18021 39601 18055
rect 39144 17933 39178 17959
rect 39144 17925 39178 17933
rect 39144 17865 39178 17887
rect 39144 17853 39178 17865
rect 39144 17797 39178 17815
rect 39144 17781 39178 17797
rect 39144 17729 39178 17743
rect 39144 17709 39178 17729
rect 39144 17661 39178 17671
rect 39144 17637 39178 17661
rect 39144 17593 39178 17599
rect 39144 17565 39178 17593
rect 39144 17525 39178 17527
rect 39144 17493 39178 17525
rect 39144 17423 39178 17455
rect 39144 17421 39178 17423
rect 39144 17355 39178 17383
rect 39144 17349 39178 17355
rect 39144 17287 39178 17311
rect 39144 17277 39178 17287
rect 39144 17219 39178 17239
rect 39144 17205 39178 17219
rect 39144 17151 39178 17167
rect 39144 17133 39178 17151
rect 39144 17083 39178 17095
rect 39144 17061 39178 17083
rect 39144 17015 39178 17023
rect 39144 16989 39178 17015
rect 39402 17933 39436 17959
rect 39402 17925 39436 17933
rect 39402 17865 39436 17887
rect 39402 17853 39436 17865
rect 39402 17797 39436 17815
rect 39402 17781 39436 17797
rect 39402 17729 39436 17743
rect 39402 17709 39436 17729
rect 39402 17661 39436 17671
rect 39402 17637 39436 17661
rect 39402 17593 39436 17599
rect 39402 17565 39436 17593
rect 39402 17525 39436 17527
rect 39402 17493 39436 17525
rect 39402 17423 39436 17455
rect 39402 17421 39436 17423
rect 39402 17355 39436 17383
rect 39402 17349 39436 17355
rect 39402 17287 39436 17311
rect 39402 17277 39436 17287
rect 39402 17219 39436 17239
rect 39402 17205 39436 17219
rect 39402 17151 39436 17167
rect 39402 17133 39436 17151
rect 39402 17083 39436 17095
rect 39402 17061 39436 17083
rect 39402 17015 39436 17023
rect 39402 16989 39436 17015
rect 39660 17933 39694 17959
rect 39660 17925 39694 17933
rect 39660 17865 39694 17887
rect 39660 17853 39694 17865
rect 39660 17797 39694 17815
rect 39660 17781 39694 17797
rect 39660 17729 39694 17743
rect 39660 17709 39694 17729
rect 39660 17661 39694 17671
rect 39660 17637 39694 17661
rect 39660 17593 39694 17599
rect 39660 17565 39694 17593
rect 39660 17525 39694 17527
rect 39660 17493 39694 17525
rect 39660 17423 39694 17455
rect 39660 17421 39694 17423
rect 39660 17355 39694 17383
rect 39660 17349 39694 17355
rect 39660 17287 39694 17311
rect 39660 17277 39694 17287
rect 39660 17219 39694 17239
rect 39660 17205 39694 17219
rect 39660 17151 39694 17167
rect 39660 17133 39694 17151
rect 39660 17083 39694 17095
rect 39660 17061 39694 17083
rect 39660 17015 39694 17023
rect 39660 16989 39694 17015
rect 24208 16687 24242 16689
rect 24208 16655 24242 16687
rect 24208 16585 24242 16617
rect 24208 16583 24242 16585
rect 39237 16893 39239 16927
rect 39239 16893 39271 16927
rect 39309 16893 39341 16927
rect 39341 16893 39343 16927
rect 39495 16893 39497 16927
rect 39497 16893 39529 16927
rect 39567 16893 39599 16927
rect 39599 16893 39601 16927
rect 23150 16511 23184 16517
rect 23150 16449 23184 16473
rect 23150 16439 23184 16449
rect 23150 16381 23184 16401
rect 24208 16517 24242 16545
rect 24208 16511 24242 16517
rect 24208 16449 24242 16473
rect 24208 16439 24242 16449
rect 23150 16367 23184 16381
rect 23150 16313 23184 16329
rect 23150 16295 23184 16313
rect 23150 16245 23184 16257
rect 23150 16223 23184 16245
rect 23150 16177 23184 16185
rect 23150 16151 23184 16177
rect 24208 16381 24242 16401
rect 24208 16367 24242 16381
rect 24208 16313 24242 16329
rect 24208 16295 24242 16313
rect 24208 16245 24242 16257
rect 24208 16223 24242 16245
rect 24208 16177 24242 16185
rect 24208 16151 24242 16177
rect 23247 16064 23271 16098
rect 23271 16064 23281 16098
rect 23319 16064 23339 16098
rect 23339 16064 23353 16098
rect 23391 16064 23407 16098
rect 23407 16064 23425 16098
rect 23463 16064 23475 16098
rect 23475 16064 23497 16098
rect 23535 16064 23543 16098
rect 23543 16064 23569 16098
rect 23607 16064 23611 16098
rect 23611 16064 23641 16098
rect 23679 16064 23713 16098
rect 23751 16064 23781 16098
rect 23781 16064 23785 16098
rect 23823 16064 23849 16098
rect 23849 16064 23857 16098
rect 23895 16064 23917 16098
rect 23917 16064 23929 16098
rect 23967 16064 23985 16098
rect 23985 16064 24001 16098
rect 24039 16064 24053 16098
rect 24053 16064 24073 16098
rect 24111 16064 24121 16098
rect 24121 16064 24145 16098
rect 24609 16568 24643 16602
rect 24681 16568 24715 16602
rect 24753 16568 24787 16602
rect 24825 16568 24859 16602
rect 24897 16568 24931 16602
rect 24969 16568 25003 16602
rect 27140 16568 27174 16602
rect 27212 16568 27246 16602
rect 27284 16568 27318 16602
rect 27356 16568 27390 16602
rect 27428 16568 27462 16602
rect 27500 16568 27534 16602
rect 42612 18778 42646 18796
rect 42612 18762 42646 18778
rect 42612 18710 42646 18724
rect 42612 18690 42646 18710
rect 42612 18642 42646 18652
rect 42612 18618 42646 18642
rect 42612 18574 42646 18580
rect 42612 18546 42646 18574
rect 42612 18506 42646 18508
rect 42612 18474 42646 18506
rect 42612 18404 42646 18436
rect 42612 18402 42646 18404
rect 42612 18336 42646 18364
rect 42612 18330 42646 18336
rect 42612 18268 42646 18292
rect 42612 18258 42646 18268
rect 42612 18200 42646 18220
rect 42612 18186 42646 18200
rect 42612 18132 42646 18148
rect 42612 18114 42646 18132
rect 42612 18064 42646 18076
rect 42612 18042 42646 18064
rect 42612 17996 42646 18004
rect 42612 17970 42646 17996
rect 42612 17928 42646 17932
rect 42612 17898 42646 17928
rect 42612 17826 42646 17860
rect 42612 17758 42646 17788
rect 42612 17754 42646 17758
rect 42612 17690 42646 17716
rect 42612 17682 42646 17690
rect 42612 17622 42646 17644
rect 42612 17610 42646 17622
rect 42612 17554 42646 17572
rect 42612 17538 42646 17554
rect 42612 17486 42646 17500
rect 42612 17466 42646 17486
rect 42612 17418 42646 17428
rect 42612 17394 42646 17418
rect 42612 17350 42646 17356
rect 42612 17322 42646 17350
rect 42612 17282 42646 17284
rect 42612 17250 42646 17282
rect 42612 17180 42646 17212
rect 42612 17178 42646 17180
rect 42612 17112 42646 17140
rect 42612 17106 42646 17112
rect 42612 17044 42646 17068
rect 42612 17034 42646 17044
rect 42612 16976 42646 16996
rect 42612 16962 42646 16976
rect 42612 16908 42646 16924
rect 42612 16890 42646 16908
rect 42870 18778 42904 18796
rect 42870 18762 42904 18778
rect 42870 18710 42904 18724
rect 42870 18690 42904 18710
rect 42870 18642 42904 18652
rect 42870 18618 42904 18642
rect 42870 18574 42904 18580
rect 42870 18546 42904 18574
rect 42870 18506 42904 18508
rect 42870 18474 42904 18506
rect 42870 18404 42904 18436
rect 42870 18402 42904 18404
rect 42870 18336 42904 18364
rect 42870 18330 42904 18336
rect 42870 18268 42904 18292
rect 42870 18258 42904 18268
rect 42870 18200 42904 18220
rect 42870 18186 42904 18200
rect 42870 18132 42904 18148
rect 42870 18114 42904 18132
rect 42870 18064 42904 18076
rect 42870 18042 42904 18064
rect 42870 17996 42904 18004
rect 42870 17970 42904 17996
rect 42870 17928 42904 17932
rect 42870 17898 42904 17928
rect 42870 17826 42904 17860
rect 42870 17758 42904 17788
rect 42870 17754 42904 17758
rect 42870 17690 42904 17716
rect 42870 17682 42904 17690
rect 42870 17622 42904 17644
rect 42870 17610 42904 17622
rect 42870 17554 42904 17572
rect 42870 17538 42904 17554
rect 42870 17486 42904 17500
rect 42870 17466 42904 17486
rect 42870 17418 42904 17428
rect 42870 17394 42904 17418
rect 42870 17350 42904 17356
rect 42870 17322 42904 17350
rect 42870 17282 42904 17284
rect 42870 17250 42904 17282
rect 42870 17180 42904 17212
rect 42870 17178 42904 17180
rect 42870 17112 42904 17140
rect 42870 17106 42904 17112
rect 42870 17044 42904 17068
rect 42870 17034 42904 17044
rect 42870 16976 42904 16996
rect 42870 16962 42904 16976
rect 42870 16908 42904 16924
rect 42870 16890 42904 16908
rect 43128 18778 43162 18796
rect 43128 18762 43162 18778
rect 43128 18710 43162 18724
rect 43128 18690 43162 18710
rect 43128 18642 43162 18652
rect 43128 18618 43162 18642
rect 43128 18574 43162 18580
rect 43128 18546 43162 18574
rect 43128 18506 43162 18508
rect 43128 18474 43162 18506
rect 43128 18404 43162 18436
rect 43128 18402 43162 18404
rect 43128 18336 43162 18364
rect 43128 18330 43162 18336
rect 43128 18268 43162 18292
rect 43128 18258 43162 18268
rect 43128 18200 43162 18220
rect 43128 18186 43162 18200
rect 43128 18132 43162 18148
rect 43128 18114 43162 18132
rect 43128 18064 43162 18076
rect 43128 18042 43162 18064
rect 43128 17996 43162 18004
rect 43128 17970 43162 17996
rect 43128 17928 43162 17932
rect 43128 17898 43162 17928
rect 43128 17826 43162 17860
rect 43128 17758 43162 17788
rect 43128 17754 43162 17758
rect 43128 17690 43162 17716
rect 43128 17682 43162 17690
rect 43128 17622 43162 17644
rect 43128 17610 43162 17622
rect 43128 17554 43162 17572
rect 43128 17538 43162 17554
rect 43128 17486 43162 17500
rect 43128 17466 43162 17486
rect 43128 17418 43162 17428
rect 43128 17394 43162 17418
rect 43128 17350 43162 17356
rect 43128 17322 43162 17350
rect 43128 17282 43162 17284
rect 43128 17250 43162 17282
rect 43128 17180 43162 17212
rect 43128 17178 43162 17180
rect 43128 17112 43162 17140
rect 43128 17106 43162 17112
rect 43128 17044 43162 17068
rect 43128 17034 43162 17044
rect 43128 16976 43162 16996
rect 43128 16962 43162 16976
rect 43128 16908 43162 16924
rect 43128 16890 43162 16908
rect 43386 18778 43420 18796
rect 43386 18762 43420 18778
rect 43386 18710 43420 18724
rect 43386 18690 43420 18710
rect 43386 18642 43420 18652
rect 43386 18618 43420 18642
rect 43386 18574 43420 18580
rect 43386 18546 43420 18574
rect 43386 18506 43420 18508
rect 43386 18474 43420 18506
rect 43386 18404 43420 18436
rect 43386 18402 43420 18404
rect 43386 18336 43420 18364
rect 43386 18330 43420 18336
rect 43386 18268 43420 18292
rect 43386 18258 43420 18268
rect 43386 18200 43420 18220
rect 43386 18186 43420 18200
rect 43386 18132 43420 18148
rect 43386 18114 43420 18132
rect 43386 18064 43420 18076
rect 43386 18042 43420 18064
rect 43386 17996 43420 18004
rect 43386 17970 43420 17996
rect 43386 17928 43420 17932
rect 43386 17898 43420 17928
rect 43386 17826 43420 17860
rect 43386 17758 43420 17788
rect 43386 17754 43420 17758
rect 43386 17690 43420 17716
rect 43386 17682 43420 17690
rect 43386 17622 43420 17644
rect 43386 17610 43420 17622
rect 43386 17554 43420 17572
rect 43386 17538 43420 17554
rect 43386 17486 43420 17500
rect 43386 17466 43420 17486
rect 43386 17418 43420 17428
rect 43386 17394 43420 17418
rect 43386 17350 43420 17356
rect 43386 17322 43420 17350
rect 43386 17282 43420 17284
rect 43386 17250 43420 17282
rect 43386 17180 43420 17212
rect 43386 17178 43420 17180
rect 43386 17112 43420 17140
rect 43386 17106 43420 17112
rect 43386 17044 43420 17068
rect 43386 17034 43420 17044
rect 43386 16976 43420 16996
rect 43386 16962 43420 16976
rect 43386 16908 43420 16924
rect 43386 16890 43420 16908
rect 43644 18778 43678 18796
rect 43644 18762 43678 18778
rect 43644 18710 43678 18724
rect 43644 18690 43678 18710
rect 43644 18642 43678 18652
rect 43644 18618 43678 18642
rect 43644 18574 43678 18580
rect 43644 18546 43678 18574
rect 43644 18506 43678 18508
rect 43644 18474 43678 18506
rect 43644 18404 43678 18436
rect 43644 18402 43678 18404
rect 43644 18336 43678 18364
rect 43644 18330 43678 18336
rect 43644 18268 43678 18292
rect 43644 18258 43678 18268
rect 43644 18200 43678 18220
rect 43644 18186 43678 18200
rect 43644 18132 43678 18148
rect 43644 18114 43678 18132
rect 43644 18064 43678 18076
rect 43644 18042 43678 18064
rect 43644 17996 43678 18004
rect 43644 17970 43678 17996
rect 43644 17928 43678 17932
rect 43644 17898 43678 17928
rect 43644 17826 43678 17860
rect 43644 17758 43678 17788
rect 43644 17754 43678 17758
rect 43644 17690 43678 17716
rect 43644 17682 43678 17690
rect 43644 17622 43678 17644
rect 43644 17610 43678 17622
rect 43644 17554 43678 17572
rect 43644 17538 43678 17554
rect 43644 17486 43678 17500
rect 43644 17466 43678 17486
rect 43644 17418 43678 17428
rect 43644 17394 43678 17418
rect 43644 17350 43678 17356
rect 43644 17322 43678 17350
rect 43644 17282 43678 17284
rect 43644 17250 43678 17282
rect 43644 17180 43678 17212
rect 43644 17178 43678 17180
rect 43644 17112 43678 17140
rect 43644 17106 43678 17112
rect 43644 17044 43678 17068
rect 43644 17034 43678 17044
rect 43644 16976 43678 16996
rect 43644 16962 43678 16976
rect 43644 16908 43678 16924
rect 43644 16890 43678 16908
rect 43902 18778 43936 18796
rect 43902 18762 43936 18778
rect 43902 18710 43936 18724
rect 43902 18690 43936 18710
rect 43902 18642 43936 18652
rect 43902 18618 43936 18642
rect 43902 18574 43936 18580
rect 43902 18546 43936 18574
rect 43902 18506 43936 18508
rect 43902 18474 43936 18506
rect 43902 18404 43936 18436
rect 43902 18402 43936 18404
rect 43902 18336 43936 18364
rect 43902 18330 43936 18336
rect 43902 18268 43936 18292
rect 43902 18258 43936 18268
rect 43902 18200 43936 18220
rect 43902 18186 43936 18200
rect 43902 18132 43936 18148
rect 43902 18114 43936 18132
rect 43902 18064 43936 18076
rect 43902 18042 43936 18064
rect 43902 17996 43936 18004
rect 43902 17970 43936 17996
rect 43902 17928 43936 17932
rect 43902 17898 43936 17928
rect 43902 17826 43936 17860
rect 43902 17758 43936 17788
rect 43902 17754 43936 17758
rect 43902 17690 43936 17716
rect 43902 17682 43936 17690
rect 43902 17622 43936 17644
rect 43902 17610 43936 17622
rect 43902 17554 43936 17572
rect 43902 17538 43936 17554
rect 43902 17486 43936 17500
rect 43902 17466 43936 17486
rect 43902 17418 43936 17428
rect 43902 17394 43936 17418
rect 43902 17350 43936 17356
rect 43902 17322 43936 17350
rect 43902 17282 43936 17284
rect 43902 17250 43936 17282
rect 43902 17180 43936 17212
rect 43902 17178 43936 17180
rect 43902 17112 43936 17140
rect 43902 17106 43936 17112
rect 43902 17044 43936 17068
rect 43902 17034 43936 17044
rect 43902 16976 43936 16996
rect 43902 16962 43936 16976
rect 43902 16908 43936 16924
rect 43902 16890 43936 16908
rect 44160 18778 44194 18796
rect 44160 18762 44194 18778
rect 44160 18710 44194 18724
rect 44160 18690 44194 18710
rect 44160 18642 44194 18652
rect 44160 18618 44194 18642
rect 44160 18574 44194 18580
rect 44160 18546 44194 18574
rect 44160 18506 44194 18508
rect 44160 18474 44194 18506
rect 44160 18404 44194 18436
rect 44160 18402 44194 18404
rect 44160 18336 44194 18364
rect 44160 18330 44194 18336
rect 44160 18268 44194 18292
rect 44160 18258 44194 18268
rect 44160 18200 44194 18220
rect 44160 18186 44194 18200
rect 44160 18132 44194 18148
rect 44160 18114 44194 18132
rect 44160 18064 44194 18076
rect 44160 18042 44194 18064
rect 44160 17996 44194 18004
rect 44160 17970 44194 17996
rect 44160 17928 44194 17932
rect 44160 17898 44194 17928
rect 44160 17826 44194 17860
rect 44160 17758 44194 17788
rect 44160 17754 44194 17758
rect 44160 17690 44194 17716
rect 44160 17682 44194 17690
rect 44160 17622 44194 17644
rect 44160 17610 44194 17622
rect 44160 17554 44194 17572
rect 44160 17538 44194 17554
rect 44160 17486 44194 17500
rect 44160 17466 44194 17486
rect 44160 17418 44194 17428
rect 44160 17394 44194 17418
rect 44160 17350 44194 17356
rect 44160 17322 44194 17350
rect 44160 17282 44194 17284
rect 44160 17250 44194 17282
rect 44160 17180 44194 17212
rect 44160 17178 44194 17180
rect 44160 17112 44194 17140
rect 44160 17106 44194 17112
rect 44160 17044 44194 17068
rect 44160 17034 44194 17044
rect 44160 16976 44194 16996
rect 44160 16962 44194 16976
rect 44160 16908 44194 16924
rect 44160 16890 44194 16908
rect 44418 18778 44452 18796
rect 44418 18762 44452 18778
rect 44418 18710 44452 18724
rect 44418 18690 44452 18710
rect 44418 18642 44452 18652
rect 44418 18618 44452 18642
rect 44418 18574 44452 18580
rect 44418 18546 44452 18574
rect 44418 18506 44452 18508
rect 44418 18474 44452 18506
rect 44418 18404 44452 18436
rect 44418 18402 44452 18404
rect 44418 18336 44452 18364
rect 44418 18330 44452 18336
rect 44418 18268 44452 18292
rect 44418 18258 44452 18268
rect 44418 18200 44452 18220
rect 44418 18186 44452 18200
rect 44418 18132 44452 18148
rect 44418 18114 44452 18132
rect 44418 18064 44452 18076
rect 44418 18042 44452 18064
rect 44418 17996 44452 18004
rect 44418 17970 44452 17996
rect 44418 17928 44452 17932
rect 44418 17898 44452 17928
rect 44418 17826 44452 17860
rect 44418 17758 44452 17788
rect 44418 17754 44452 17758
rect 44418 17690 44452 17716
rect 44418 17682 44452 17690
rect 44418 17622 44452 17644
rect 44418 17610 44452 17622
rect 44418 17554 44452 17572
rect 44418 17538 44452 17554
rect 44418 17486 44452 17500
rect 44418 17466 44452 17486
rect 44418 17418 44452 17428
rect 44418 17394 44452 17418
rect 44418 17350 44452 17356
rect 44418 17322 44452 17350
rect 44418 17282 44452 17284
rect 44418 17250 44452 17282
rect 44418 17180 44452 17212
rect 44418 17178 44452 17180
rect 44418 17112 44452 17140
rect 44418 17106 44452 17112
rect 44418 17044 44452 17068
rect 44418 17034 44452 17044
rect 44418 16976 44452 16996
rect 44418 16962 44452 16976
rect 44418 16908 44452 16924
rect 44418 16890 44452 16908
rect 44676 18778 44710 18796
rect 44676 18762 44710 18778
rect 44676 18710 44710 18724
rect 44676 18690 44710 18710
rect 44676 18642 44710 18652
rect 44676 18618 44710 18642
rect 44676 18574 44710 18580
rect 44676 18546 44710 18574
rect 44676 18506 44710 18508
rect 44676 18474 44710 18506
rect 44676 18404 44710 18436
rect 44676 18402 44710 18404
rect 44676 18336 44710 18364
rect 44676 18330 44710 18336
rect 44676 18268 44710 18292
rect 44676 18258 44710 18268
rect 44676 18200 44710 18220
rect 44676 18186 44710 18200
rect 44676 18132 44710 18148
rect 44676 18114 44710 18132
rect 44676 18064 44710 18076
rect 44676 18042 44710 18064
rect 44676 17996 44710 18004
rect 44676 17970 44710 17996
rect 44676 17928 44710 17932
rect 44676 17898 44710 17928
rect 44676 17826 44710 17860
rect 44676 17758 44710 17788
rect 44676 17754 44710 17758
rect 44676 17690 44710 17716
rect 44676 17682 44710 17690
rect 44676 17622 44710 17644
rect 44676 17610 44710 17622
rect 44676 17554 44710 17572
rect 44676 17538 44710 17554
rect 44676 17486 44710 17500
rect 44676 17466 44710 17486
rect 44676 17418 44710 17428
rect 44676 17394 44710 17418
rect 44676 17350 44710 17356
rect 44676 17322 44710 17350
rect 44676 17282 44710 17284
rect 44676 17250 44710 17282
rect 44676 17180 44710 17212
rect 44676 17178 44710 17180
rect 44676 17112 44710 17140
rect 44676 17106 44710 17112
rect 44676 17044 44710 17068
rect 44676 17034 44710 17044
rect 44676 16976 44710 16996
rect 44676 16962 44710 16976
rect 44676 16908 44710 16924
rect 44676 16890 44710 16908
rect 44934 18778 44968 18796
rect 44934 18762 44968 18778
rect 44934 18710 44968 18724
rect 44934 18690 44968 18710
rect 44934 18642 44968 18652
rect 44934 18618 44968 18642
rect 44934 18574 44968 18580
rect 44934 18546 44968 18574
rect 44934 18506 44968 18508
rect 44934 18474 44968 18506
rect 44934 18404 44968 18436
rect 44934 18402 44968 18404
rect 44934 18336 44968 18364
rect 44934 18330 44968 18336
rect 44934 18268 44968 18292
rect 44934 18258 44968 18268
rect 44934 18200 44968 18220
rect 44934 18186 44968 18200
rect 44934 18132 44968 18148
rect 44934 18114 44968 18132
rect 44934 18064 44968 18076
rect 44934 18042 44968 18064
rect 44934 17996 44968 18004
rect 44934 17970 44968 17996
rect 44934 17928 44968 17932
rect 44934 17898 44968 17928
rect 44934 17826 44968 17860
rect 44934 17758 44968 17788
rect 44934 17754 44968 17758
rect 44934 17690 44968 17716
rect 44934 17682 44968 17690
rect 44934 17622 44968 17644
rect 44934 17610 44968 17622
rect 44934 17554 44968 17572
rect 44934 17538 44968 17554
rect 44934 17486 44968 17500
rect 44934 17466 44968 17486
rect 44934 17418 44968 17428
rect 44934 17394 44968 17418
rect 44934 17350 44968 17356
rect 44934 17322 44968 17350
rect 44934 17282 44968 17284
rect 44934 17250 44968 17282
rect 44934 17180 44968 17212
rect 44934 17178 44968 17180
rect 44934 17112 44968 17140
rect 44934 17106 44968 17112
rect 44934 17044 44968 17068
rect 44934 17034 44968 17044
rect 44934 16976 44968 16996
rect 44934 16962 44968 16976
rect 44934 16908 44968 16924
rect 44934 16890 44968 16908
rect 45192 18778 45226 18796
rect 45192 18762 45226 18778
rect 45192 18710 45226 18724
rect 45192 18690 45226 18710
rect 45192 18642 45226 18652
rect 45192 18618 45226 18642
rect 45192 18574 45226 18580
rect 45192 18546 45226 18574
rect 45192 18506 45226 18508
rect 45192 18474 45226 18506
rect 45192 18404 45226 18436
rect 45192 18402 45226 18404
rect 45192 18336 45226 18364
rect 45192 18330 45226 18336
rect 45192 18268 45226 18292
rect 45192 18258 45226 18268
rect 45192 18200 45226 18220
rect 45192 18186 45226 18200
rect 45192 18132 45226 18148
rect 45192 18114 45226 18132
rect 45192 18064 45226 18076
rect 45192 18042 45226 18064
rect 45192 17996 45226 18004
rect 45192 17970 45226 17996
rect 45192 17928 45226 17932
rect 45192 17898 45226 17928
rect 45192 17826 45226 17860
rect 45192 17758 45226 17788
rect 45192 17754 45226 17758
rect 45192 17690 45226 17716
rect 45192 17682 45226 17690
rect 45192 17622 45226 17644
rect 45192 17610 45226 17622
rect 45192 17554 45226 17572
rect 45192 17538 45226 17554
rect 45192 17486 45226 17500
rect 45192 17466 45226 17486
rect 45192 17418 45226 17428
rect 45192 17394 45226 17418
rect 45192 17350 45226 17356
rect 45192 17322 45226 17350
rect 45192 17282 45226 17284
rect 45192 17250 45226 17282
rect 45192 17180 45226 17212
rect 45192 17178 45226 17180
rect 45192 17112 45226 17140
rect 45192 17106 45226 17112
rect 45192 17044 45226 17068
rect 45192 17034 45226 17044
rect 45192 16976 45226 16996
rect 45192 16962 45226 16976
rect 45192 16908 45226 16924
rect 45192 16890 45226 16908
rect 42705 16762 42707 16796
rect 42707 16762 42739 16796
rect 42777 16762 42809 16796
rect 42809 16762 42811 16796
rect 42963 16762 42965 16796
rect 42965 16762 42997 16796
rect 43035 16762 43067 16796
rect 43067 16762 43069 16796
rect 43221 16762 43223 16796
rect 43223 16762 43255 16796
rect 43293 16762 43325 16796
rect 43325 16762 43327 16796
rect 43479 16762 43481 16796
rect 43481 16762 43513 16796
rect 43551 16762 43583 16796
rect 43583 16762 43585 16796
rect 43737 16762 43739 16796
rect 43739 16762 43771 16796
rect 43809 16762 43841 16796
rect 43841 16762 43843 16796
rect 43995 16762 43997 16796
rect 43997 16762 44029 16796
rect 44067 16762 44099 16796
rect 44099 16762 44101 16796
rect 44253 16762 44255 16796
rect 44255 16762 44287 16796
rect 44325 16762 44357 16796
rect 44357 16762 44359 16796
rect 44511 16762 44513 16796
rect 44513 16762 44545 16796
rect 44583 16762 44615 16796
rect 44615 16762 44617 16796
rect 44769 16762 44771 16796
rect 44771 16762 44803 16796
rect 44841 16762 44873 16796
rect 44873 16762 44875 16796
rect 45027 16762 45029 16796
rect 45029 16762 45061 16796
rect 45099 16762 45131 16796
rect 45131 16762 45133 16796
rect 24609 16250 24643 16284
rect 24681 16250 24715 16284
rect 24753 16250 24787 16284
rect 24825 16250 24859 16284
rect 24897 16250 24931 16284
rect 24969 16250 25003 16284
rect 27140 16250 27174 16284
rect 27212 16250 27246 16284
rect 27284 16250 27318 16284
rect 27356 16250 27390 16284
rect 27428 16250 27462 16284
rect 27500 16250 27534 16284
rect 24609 15932 24643 15966
rect 24681 15932 24715 15966
rect 24753 15932 24787 15966
rect 24825 15932 24859 15966
rect 24897 15932 24931 15966
rect 24969 15932 25003 15966
rect 27140 15932 27174 15966
rect 27212 15932 27246 15966
rect 27284 15932 27318 15966
rect 27356 15932 27390 15966
rect 27428 15932 27462 15966
rect 27500 15932 27534 15966
rect -3862 14851 -3828 14885
rect -3862 14779 -3828 14813
rect -3862 14707 -3828 14741
rect -3862 14635 -3828 14669
rect -3862 14563 -3828 14597
rect -3862 14491 -3828 14525
rect -3862 12820 -3828 12854
rect -3862 12748 -3828 12782
rect -3862 12676 -3828 12710
rect -3862 12604 -3828 12638
rect -3862 12532 -3828 12566
rect -3862 12460 -3828 12494
rect 13091 14814 13115 14848
rect 13115 14814 13125 14848
rect 13163 14814 13183 14848
rect 13183 14814 13197 14848
rect 13235 14814 13251 14848
rect 13251 14814 13269 14848
rect 13307 14814 13319 14848
rect 13319 14814 13341 14848
rect 13379 14814 13387 14848
rect 13387 14814 13413 14848
rect 13451 14814 13455 14848
rect 13455 14814 13485 14848
rect 13523 14814 13557 14848
rect 13595 14814 13625 14848
rect 13625 14814 13629 14848
rect 13667 14814 13693 14848
rect 13693 14814 13701 14848
rect 13739 14814 13761 14848
rect 13761 14814 13773 14848
rect 13811 14814 13829 14848
rect 13829 14814 13845 14848
rect 13883 14814 13897 14848
rect 13897 14814 13917 14848
rect 13955 14814 13965 14848
rect 13965 14814 13989 14848
rect 14149 14814 14173 14848
rect 14173 14814 14183 14848
rect 14221 14814 14241 14848
rect 14241 14814 14255 14848
rect 14293 14814 14309 14848
rect 14309 14814 14327 14848
rect 14365 14814 14377 14848
rect 14377 14814 14399 14848
rect 14437 14814 14445 14848
rect 14445 14814 14471 14848
rect 14509 14814 14513 14848
rect 14513 14814 14543 14848
rect 14581 14814 14615 14848
rect 14653 14814 14683 14848
rect 14683 14814 14687 14848
rect 14725 14814 14751 14848
rect 14751 14814 14759 14848
rect 14797 14814 14819 14848
rect 14819 14814 14831 14848
rect 14869 14814 14887 14848
rect 14887 14814 14903 14848
rect 14941 14814 14955 14848
rect 14955 14814 14975 14848
rect 15013 14814 15023 14848
rect 15023 14814 15047 14848
rect 12994 14712 13028 14724
rect 12994 14690 13028 14712
rect 12994 14644 13028 14652
rect 12994 14618 13028 14644
rect 12994 14576 13028 14580
rect 12994 14546 13028 14576
rect 12994 14474 13028 14508
rect 12994 14406 13028 14436
rect 12994 14402 13028 14406
rect 12994 14338 13028 14364
rect 12994 14330 13028 14338
rect 12994 14270 13028 14292
rect 12994 14258 13028 14270
rect 12994 14202 13028 14220
rect 12994 14186 13028 14202
rect 12994 14134 13028 14148
rect 12994 14114 13028 14134
rect 12994 14066 13028 14076
rect 12994 14042 13028 14066
rect 12994 13998 13028 14004
rect 12994 13970 13028 13998
rect 12994 13930 13028 13932
rect 12994 13898 13028 13930
rect 12994 13828 13028 13860
rect 12994 13826 13028 13828
rect 12994 13760 13028 13788
rect 12994 13754 13028 13760
rect 12994 13692 13028 13716
rect 12994 13682 13028 13692
rect 12994 13624 13028 13644
rect 12994 13610 13028 13624
rect 12994 13556 13028 13572
rect 12994 13538 13028 13556
rect 12994 13488 13028 13500
rect 12994 13466 13028 13488
rect 12994 13420 13028 13428
rect 12994 13394 13028 13420
rect 12994 13352 13028 13356
rect 12994 13322 13028 13352
rect 12994 13250 13028 13284
rect 12994 13182 13028 13212
rect 12994 13178 13028 13182
rect 12994 13114 13028 13140
rect 12994 13106 13028 13114
rect 12994 13046 13028 13068
rect 12994 13034 13028 13046
rect 12994 12978 13028 12996
rect 12994 12962 13028 12978
rect 12994 12910 13028 12924
rect 12994 12890 13028 12910
rect 12994 12842 13028 12852
rect 12994 12818 13028 12842
rect 12994 12774 13028 12780
rect 12994 12746 13028 12774
rect 12994 12706 13028 12708
rect 12994 12674 13028 12706
rect 12994 12604 13028 12636
rect 12994 12602 13028 12604
rect 12994 12536 13028 12564
rect 12994 12530 13028 12536
rect 12994 12468 13028 12492
rect 12994 12458 13028 12468
rect 12994 12400 13028 12420
rect 12994 12386 13028 12400
rect 12994 12332 13028 12348
rect 12994 12314 13028 12332
rect 12994 12264 13028 12276
rect 12994 12242 13028 12264
rect 12994 12196 13028 12204
rect 12994 12170 13028 12196
rect 12994 12128 13028 12132
rect 12994 12098 13028 12128
rect 12994 12026 13028 12060
rect 12994 11958 13028 11988
rect 12994 11954 13028 11958
rect 12994 11890 13028 11916
rect 12994 11882 13028 11890
rect 12994 11822 13028 11844
rect 12994 11810 13028 11822
rect 14052 14712 14086 14724
rect 14052 14690 14086 14712
rect 14052 14644 14086 14652
rect 14052 14618 14086 14644
rect 14052 14576 14086 14580
rect 14052 14546 14086 14576
rect 14052 14474 14086 14508
rect 14052 14406 14086 14436
rect 14052 14402 14086 14406
rect 14052 14338 14086 14364
rect 14052 14330 14086 14338
rect 14052 14270 14086 14292
rect 14052 14258 14086 14270
rect 14052 14202 14086 14220
rect 14052 14186 14086 14202
rect 14052 14134 14086 14148
rect 14052 14114 14086 14134
rect 14052 14066 14086 14076
rect 14052 14042 14086 14066
rect 14052 13998 14086 14004
rect 14052 13970 14086 13998
rect 14052 13930 14086 13932
rect 14052 13898 14086 13930
rect 14052 13828 14086 13860
rect 14052 13826 14086 13828
rect 14052 13760 14086 13788
rect 14052 13754 14086 13760
rect 14052 13692 14086 13716
rect 14052 13682 14086 13692
rect 14052 13624 14086 13644
rect 14052 13610 14086 13624
rect 14052 13556 14086 13572
rect 14052 13538 14086 13556
rect 14052 13488 14086 13500
rect 14052 13466 14086 13488
rect 14052 13420 14086 13428
rect 14052 13394 14086 13420
rect 14052 13352 14086 13356
rect 14052 13322 14086 13352
rect 14052 13250 14086 13284
rect 14052 13182 14086 13212
rect 14052 13178 14086 13182
rect 14052 13114 14086 13140
rect 14052 13106 14086 13114
rect 14052 13046 14086 13068
rect 14052 13034 14086 13046
rect 14052 12978 14086 12996
rect 14052 12962 14086 12978
rect 14052 12910 14086 12924
rect 14052 12890 14086 12910
rect 14052 12842 14086 12852
rect 14052 12818 14086 12842
rect 14052 12774 14086 12780
rect 14052 12746 14086 12774
rect 14052 12706 14086 12708
rect 14052 12674 14086 12706
rect 14052 12604 14086 12636
rect 14052 12602 14086 12604
rect 14052 12536 14086 12564
rect 14052 12530 14086 12536
rect 14052 12468 14086 12492
rect 14052 12458 14086 12468
rect 14052 12400 14086 12420
rect 14052 12386 14086 12400
rect 14052 12332 14086 12348
rect 14052 12314 14086 12332
rect 14052 12264 14086 12276
rect 14052 12242 14086 12264
rect 14052 12196 14086 12204
rect 14052 12170 14086 12196
rect 14052 12128 14086 12132
rect 14052 12098 14086 12128
rect 14052 12026 14086 12060
rect 14052 11958 14086 11988
rect 14052 11954 14086 11958
rect 14052 11890 14086 11916
rect 14052 11882 14086 11890
rect 14052 11822 14086 11844
rect 14052 11810 14086 11822
rect 15110 14712 15144 14724
rect 15110 14690 15144 14712
rect 15110 14644 15144 14652
rect 15110 14618 15144 14644
rect 15110 14576 15144 14580
rect 15110 14546 15144 14576
rect 15110 14474 15144 14508
rect 15110 14406 15144 14436
rect 15110 14402 15144 14406
rect 15110 14338 15144 14364
rect 15110 14330 15144 14338
rect 15110 14270 15144 14292
rect 15110 14258 15144 14270
rect 15110 14202 15144 14220
rect 15110 14186 15144 14202
rect 15110 14134 15144 14148
rect 15110 14114 15144 14134
rect 15110 14066 15144 14076
rect 15110 14042 15144 14066
rect 15110 13998 15144 14004
rect 15110 13970 15144 13998
rect 15110 13930 15144 13932
rect 15110 13898 15144 13930
rect 15110 13828 15144 13860
rect 15110 13826 15144 13828
rect 15110 13760 15144 13788
rect 15110 13754 15144 13760
rect 15110 13692 15144 13716
rect 15110 13682 15144 13692
rect 15110 13624 15144 13644
rect 15110 13610 15144 13624
rect 15110 13556 15144 13572
rect 15110 13538 15144 13556
rect 15110 13488 15144 13500
rect 15110 13466 15144 13488
rect 15110 13420 15144 13428
rect 15110 13394 15144 13420
rect 15110 13352 15144 13356
rect 15110 13322 15144 13352
rect 15110 13250 15144 13284
rect 15110 13182 15144 13212
rect 15110 13178 15144 13182
rect 15110 13114 15144 13140
rect 15110 13106 15144 13114
rect 15110 13046 15144 13068
rect 15110 13034 15144 13046
rect 15110 12978 15144 12996
rect 15110 12962 15144 12978
rect 15110 12910 15144 12924
rect 15110 12890 15144 12910
rect 15110 12842 15144 12852
rect 15110 12818 15144 12842
rect 15110 12774 15144 12780
rect 15110 12746 15144 12774
rect 15110 12706 15144 12708
rect 15110 12674 15144 12706
rect 15110 12604 15144 12636
rect 15110 12602 15144 12604
rect 15110 12536 15144 12564
rect 15110 12530 15144 12536
rect 15110 12468 15144 12492
rect 15110 12458 15144 12468
rect 15110 12400 15144 12420
rect 15110 12386 15144 12400
rect 15110 12332 15144 12348
rect 15110 12314 15144 12332
rect 15110 12264 15144 12276
rect 15110 12242 15144 12264
rect 15110 12196 15144 12204
rect 15110 12170 15144 12196
rect 15110 12128 15144 12132
rect 15110 12098 15144 12128
rect 15110 12026 15144 12060
rect 15110 11958 15144 11988
rect 15110 11954 15144 11958
rect 15110 11890 15144 11916
rect 15110 11882 15144 11890
rect 15110 11822 15144 11844
rect 15110 11810 15144 11822
rect 13091 11686 13115 11720
rect 13115 11686 13125 11720
rect 13163 11686 13183 11720
rect 13183 11686 13197 11720
rect 13235 11686 13251 11720
rect 13251 11686 13269 11720
rect 13307 11686 13319 11720
rect 13319 11686 13341 11720
rect 13379 11686 13387 11720
rect 13387 11686 13413 11720
rect 13451 11686 13455 11720
rect 13455 11686 13485 11720
rect 13523 11686 13557 11720
rect 13595 11686 13625 11720
rect 13625 11686 13629 11720
rect 13667 11686 13693 11720
rect 13693 11686 13701 11720
rect 13739 11686 13761 11720
rect 13761 11686 13773 11720
rect 13811 11686 13829 11720
rect 13829 11686 13845 11720
rect 13883 11686 13897 11720
rect 13897 11686 13917 11720
rect 13955 11686 13965 11720
rect 13965 11686 13989 11720
rect 14149 11686 14173 11720
rect 14173 11686 14183 11720
rect 14221 11686 14241 11720
rect 14241 11686 14255 11720
rect 14293 11686 14309 11720
rect 14309 11686 14327 11720
rect 14365 11686 14377 11720
rect 14377 11686 14399 11720
rect 14437 11686 14445 11720
rect 14445 11686 14471 11720
rect 14509 11686 14513 11720
rect 14513 11686 14543 11720
rect 14581 11686 14615 11720
rect 14653 11686 14683 11720
rect 14683 11686 14687 11720
rect 14725 11686 14751 11720
rect 14751 11686 14759 11720
rect 14797 11686 14819 11720
rect 14819 11686 14831 11720
rect 14869 11686 14887 11720
rect 14887 11686 14903 11720
rect 14941 11686 14955 11720
rect 14955 11686 14975 11720
rect 15013 11686 15023 11720
rect 15023 11686 15047 11720
rect 15661 14814 15685 14848
rect 15685 14814 15695 14848
rect 15733 14814 15753 14848
rect 15753 14814 15767 14848
rect 15805 14814 15821 14848
rect 15821 14814 15839 14848
rect 15877 14814 15889 14848
rect 15889 14814 15911 14848
rect 15949 14814 15957 14848
rect 15957 14814 15983 14848
rect 16021 14814 16025 14848
rect 16025 14814 16055 14848
rect 16093 14814 16127 14848
rect 16165 14814 16195 14848
rect 16195 14814 16199 14848
rect 16237 14814 16263 14848
rect 16263 14814 16271 14848
rect 16309 14814 16331 14848
rect 16331 14814 16343 14848
rect 16381 14814 16399 14848
rect 16399 14814 16415 14848
rect 16453 14814 16467 14848
rect 16467 14814 16487 14848
rect 16525 14814 16535 14848
rect 16535 14814 16559 14848
rect 15564 14712 15598 14724
rect 15564 14690 15598 14712
rect 16622 14712 16656 14724
rect 15564 14644 15598 14652
rect 15564 14618 15598 14644
rect 15564 14576 15598 14580
rect 15564 14546 15598 14576
rect 15564 14474 15598 14508
rect 15564 14406 15598 14436
rect 16622 14690 16656 14712
rect 16622 14644 16656 14652
rect 16622 14618 16656 14644
rect 16622 14576 16656 14580
rect 16622 14546 16656 14576
rect 16622 14474 16656 14508
rect 15564 14402 15598 14406
rect 15564 14338 15598 14364
rect 15564 14330 15598 14338
rect 15564 14270 15598 14292
rect 15564 14258 15598 14270
rect 15564 14202 15598 14220
rect 15564 14186 15598 14202
rect 15564 14134 15598 14148
rect 15564 14114 15598 14134
rect 15564 14066 15598 14076
rect 15564 14042 15598 14066
rect 15564 13998 15598 14004
rect 15564 13970 15598 13998
rect 15564 13930 15598 13932
rect 15564 13898 15598 13930
rect 15564 13828 15598 13860
rect 15564 13826 15598 13828
rect 15564 13760 15598 13788
rect 15564 13754 15598 13760
rect 15564 13692 15598 13716
rect 15564 13682 15598 13692
rect 15564 13624 15598 13644
rect 15564 13610 15598 13624
rect 15564 13556 15598 13572
rect 15564 13538 15598 13556
rect 15564 13488 15598 13500
rect 15564 13466 15598 13488
rect 15564 13420 15598 13428
rect 15564 13394 15598 13420
rect 15564 13352 15598 13356
rect 15564 13322 15598 13352
rect 15564 13250 15598 13284
rect 15564 13182 15598 13212
rect 15564 13178 15598 13182
rect 15564 13114 15598 13140
rect 15564 13106 15598 13114
rect 15564 13046 15598 13068
rect 15564 13034 15598 13046
rect 15564 12978 15598 12996
rect 15564 12962 15598 12978
rect 15564 12910 15598 12924
rect 15564 12890 15598 12910
rect 15564 12842 15598 12852
rect 15564 12818 15598 12842
rect 15564 12774 15598 12780
rect 15564 12746 15598 12774
rect 15564 12706 15598 12708
rect 15564 12674 15598 12706
rect 15564 12604 15598 12636
rect 15564 12602 15598 12604
rect 15564 12536 15598 12564
rect 15564 12530 15598 12536
rect 15564 12468 15598 12492
rect 15564 12458 15598 12468
rect 15564 12400 15598 12420
rect 15564 12386 15598 12400
rect 15564 12332 15598 12348
rect 15564 12314 15598 12332
rect 15564 12264 15598 12276
rect 15564 12242 15598 12264
rect 15564 12196 15598 12204
rect 15564 12170 15598 12196
rect 15564 12128 15598 12132
rect 15564 12098 15598 12128
rect 15564 12026 15598 12060
rect 15564 11958 15598 11988
rect 15564 11954 15598 11958
rect 15564 11890 15598 11916
rect 15564 11882 15598 11890
rect 15564 11822 15598 11844
rect 15564 11810 15598 11822
rect 16622 14406 16656 14436
rect 16622 14402 16656 14406
rect 16622 14338 16656 14364
rect 16622 14330 16656 14338
rect 16622 14270 16656 14292
rect 16622 14258 16656 14270
rect 16622 14202 16656 14220
rect 16622 14186 16656 14202
rect 16622 14134 16656 14148
rect 16622 14114 16656 14134
rect 16622 14066 16656 14076
rect 16622 14042 16656 14066
rect 16622 13998 16656 14004
rect 16622 13970 16656 13998
rect 16622 13930 16656 13932
rect 16622 13898 16656 13930
rect 16622 13828 16656 13860
rect 16622 13826 16656 13828
rect 16622 13760 16656 13788
rect 16622 13754 16656 13760
rect 16622 13692 16656 13716
rect 16622 13682 16656 13692
rect 16622 13624 16656 13644
rect 16622 13610 16656 13624
rect 16622 13556 16656 13572
rect 16622 13538 16656 13556
rect 16622 13488 16656 13500
rect 16622 13466 16656 13488
rect 16622 13420 16656 13428
rect 16622 13394 16656 13420
rect 16622 13352 16656 13356
rect 16622 13322 16656 13352
rect 16622 13250 16656 13284
rect 16622 13182 16656 13212
rect 16622 13178 16656 13182
rect 16622 13114 16656 13140
rect 16622 13106 16656 13114
rect 16622 13046 16656 13068
rect 16622 13034 16656 13046
rect 16622 12978 16656 12996
rect 16622 12962 16656 12978
rect 16622 12910 16656 12924
rect 16622 12890 16656 12910
rect 16622 12842 16656 12852
rect 16622 12818 16656 12842
rect 16622 12774 16656 12780
rect 16622 12746 16656 12774
rect 16622 12706 16656 12708
rect 16622 12674 16656 12706
rect 16622 12604 16656 12636
rect 16622 12602 16656 12604
rect 16622 12536 16656 12564
rect 16622 12530 16656 12536
rect 16622 12468 16656 12492
rect 16622 12458 16656 12468
rect 16622 12400 16656 12420
rect 16622 12386 16656 12400
rect 16622 12332 16656 12348
rect 16622 12314 16656 12332
rect 16622 12264 16656 12276
rect 16622 12242 16656 12264
rect 16622 12196 16656 12204
rect 16622 12170 16656 12196
rect 16622 12128 16656 12132
rect 16622 12098 16656 12128
rect 16622 12026 16656 12060
rect 16622 11958 16656 11988
rect 16622 11954 16656 11958
rect 16622 11890 16656 11916
rect 16622 11882 16656 11890
rect 16622 11822 16656 11844
rect 16622 11810 16656 11822
rect 15661 11686 15685 11720
rect 15685 11686 15695 11720
rect 15733 11686 15753 11720
rect 15753 11686 15767 11720
rect 15805 11686 15821 11720
rect 15821 11686 15839 11720
rect 15877 11686 15889 11720
rect 15889 11686 15911 11720
rect 15949 11686 15957 11720
rect 15957 11686 15983 11720
rect 16021 11686 16025 11720
rect 16025 11686 16055 11720
rect 16093 11686 16127 11720
rect 16165 11686 16195 11720
rect 16195 11686 16199 11720
rect 16237 11686 16263 11720
rect 16263 11686 16271 11720
rect 16309 11686 16331 11720
rect 16331 11686 16343 11720
rect 16381 11686 16399 11720
rect 16399 11686 16415 11720
rect 16453 11686 16467 11720
rect 16467 11686 16487 11720
rect 16525 11686 16535 11720
rect 16535 11686 16559 11720
rect 17171 14824 17195 14858
rect 17195 14824 17205 14858
rect 17243 14824 17263 14858
rect 17263 14824 17277 14858
rect 17315 14824 17331 14858
rect 17331 14824 17349 14858
rect 17387 14824 17399 14858
rect 17399 14824 17421 14858
rect 17459 14824 17467 14858
rect 17467 14824 17493 14858
rect 17531 14824 17535 14858
rect 17535 14824 17565 14858
rect 17603 14824 17637 14858
rect 17675 14824 17705 14858
rect 17705 14824 17709 14858
rect 17747 14824 17773 14858
rect 17773 14824 17781 14858
rect 17819 14824 17841 14858
rect 17841 14824 17853 14858
rect 17891 14824 17909 14858
rect 17909 14824 17925 14858
rect 17963 14824 17977 14858
rect 17977 14824 17997 14858
rect 18035 14824 18045 14858
rect 18045 14824 18069 14858
rect 18635 14808 18659 14842
rect 18659 14808 18669 14842
rect 18707 14808 18727 14842
rect 18727 14808 18741 14842
rect 18779 14808 18795 14842
rect 18795 14808 18813 14842
rect 18851 14808 18863 14842
rect 18863 14808 18885 14842
rect 18923 14808 18931 14842
rect 18931 14808 18957 14842
rect 18995 14808 18999 14842
rect 18999 14808 19029 14842
rect 19067 14808 19101 14842
rect 19139 14808 19169 14842
rect 19169 14808 19173 14842
rect 19211 14808 19237 14842
rect 19237 14808 19245 14842
rect 19283 14808 19305 14842
rect 19305 14808 19317 14842
rect 19355 14808 19373 14842
rect 19373 14808 19389 14842
rect 19427 14808 19441 14842
rect 19441 14808 19461 14842
rect 19499 14808 19509 14842
rect 19509 14808 19533 14842
rect 17074 14722 17108 14734
rect 17074 14700 17108 14722
rect 17074 14654 17108 14662
rect 17074 14628 17108 14654
rect 17074 14586 17108 14590
rect 17074 14556 17108 14586
rect 17074 14484 17108 14518
rect 17074 14416 17108 14446
rect 17074 14412 17108 14416
rect 17074 14348 17108 14374
rect 17074 14340 17108 14348
rect 17074 14280 17108 14302
rect 17074 14268 17108 14280
rect 18132 14722 18166 14734
rect 18132 14700 18166 14722
rect 18132 14654 18166 14662
rect 18132 14628 18166 14654
rect 18132 14586 18166 14590
rect 18132 14556 18166 14586
rect 18132 14484 18166 14518
rect 18132 14416 18166 14446
rect 18132 14412 18166 14416
rect 18132 14348 18166 14374
rect 18132 14340 18166 14348
rect 18132 14280 18166 14302
rect 18132 14268 18166 14280
rect 17074 14212 17108 14230
rect 17074 14196 17108 14212
rect 17074 14144 17108 14158
rect 17074 14124 17108 14144
rect 17074 14076 17108 14086
rect 17074 14052 17108 14076
rect 17074 14008 17108 14014
rect 17074 13980 17108 14008
rect 17074 13940 17108 13942
rect 17074 13908 17108 13940
rect 17074 13838 17108 13870
rect 17074 13836 17108 13838
rect 17074 13770 17108 13798
rect 17074 13764 17108 13770
rect 17074 13702 17108 13726
rect 17074 13692 17108 13702
rect 17074 13634 17108 13654
rect 17074 13620 17108 13634
rect 17074 13566 17108 13582
rect 17074 13548 17108 13566
rect 17074 13498 17108 13510
rect 17074 13476 17108 13498
rect 17074 13430 17108 13438
rect 17074 13404 17108 13430
rect 17074 13362 17108 13366
rect 17074 13332 17108 13362
rect 17074 13260 17108 13294
rect 17074 13192 17108 13222
rect 17074 13188 17108 13192
rect 17074 13124 17108 13150
rect 17074 13116 17108 13124
rect 17074 13056 17108 13078
rect 17074 13044 17108 13056
rect 17074 12988 17108 13006
rect 17074 12972 17108 12988
rect 17074 12920 17108 12934
rect 17074 12900 17108 12920
rect 17074 12852 17108 12862
rect 17074 12828 17108 12852
rect 17074 12784 17108 12790
rect 17074 12756 17108 12784
rect 17074 12716 17108 12718
rect 17074 12684 17108 12716
rect 17074 12614 17108 12646
rect 17074 12612 17108 12614
rect 17074 12546 17108 12574
rect 17074 12540 17108 12546
rect 17074 12478 17108 12502
rect 17074 12468 17108 12478
rect 17074 12410 17108 12430
rect 17074 12396 17108 12410
rect 17074 12342 17108 12358
rect 17074 12324 17108 12342
rect 17074 12274 17108 12286
rect 17074 12252 17108 12274
rect 17074 12206 17108 12214
rect 17074 12180 17108 12206
rect 17074 12138 17108 12142
rect 17074 12108 17108 12138
rect 17074 12036 17108 12070
rect 17074 11968 17108 11998
rect 17074 11964 17108 11968
rect 17074 11900 17108 11926
rect 17074 11892 17108 11900
rect 17074 11832 17108 11854
rect 17074 11820 17108 11832
rect 18132 14212 18166 14230
rect 18132 14196 18166 14212
rect 18132 14144 18166 14158
rect 18132 14124 18166 14144
rect 18132 14076 18166 14086
rect 18132 14052 18166 14076
rect 18132 14008 18166 14014
rect 18132 13980 18166 14008
rect 18132 13940 18166 13942
rect 18132 13908 18166 13940
rect 18132 13838 18166 13870
rect 18132 13836 18166 13838
rect 18132 13770 18166 13798
rect 18132 13764 18166 13770
rect 18132 13702 18166 13726
rect 18132 13692 18166 13702
rect 18132 13634 18166 13654
rect 18132 13620 18166 13634
rect 18132 13566 18166 13582
rect 18132 13548 18166 13566
rect 18132 13498 18166 13510
rect 18132 13476 18166 13498
rect 18132 13430 18166 13438
rect 18132 13404 18166 13430
rect 18132 13362 18166 13366
rect 18132 13332 18166 13362
rect 18132 13260 18166 13294
rect 18132 13192 18166 13222
rect 18132 13188 18166 13192
rect 18132 13124 18166 13150
rect 18132 13116 18166 13124
rect 18132 13056 18166 13078
rect 18132 13044 18166 13056
rect 18132 12988 18166 13006
rect 18132 12972 18166 12988
rect 18132 12920 18166 12934
rect 18132 12900 18166 12920
rect 18132 12852 18166 12862
rect 18132 12828 18166 12852
rect 18132 12784 18166 12790
rect 18132 12756 18166 12784
rect 18132 12716 18166 12718
rect 18132 12684 18166 12716
rect 18132 12614 18166 12646
rect 18132 12612 18166 12614
rect 18132 12546 18166 12574
rect 18132 12540 18166 12546
rect 18132 12478 18166 12502
rect 18132 12468 18166 12478
rect 18132 12410 18166 12430
rect 18132 12396 18166 12410
rect 18132 12342 18166 12358
rect 18132 12324 18166 12342
rect 18132 12274 18166 12286
rect 18132 12252 18166 12274
rect 18132 12206 18166 12214
rect 18132 12180 18166 12206
rect 18132 12138 18166 12142
rect 18132 12108 18166 12138
rect 18132 12036 18166 12070
rect 18132 11968 18166 11998
rect 18132 11964 18166 11968
rect 18132 11900 18166 11926
rect 18132 11892 18166 11900
rect 18132 11832 18166 11854
rect 18132 11820 18166 11832
rect 17171 11696 17195 11730
rect 17195 11696 17205 11730
rect 17243 11696 17263 11730
rect 17263 11696 17277 11730
rect 17315 11696 17331 11730
rect 17331 11696 17349 11730
rect 17387 11696 17399 11730
rect 17399 11696 17421 11730
rect 17459 11696 17467 11730
rect 17467 11696 17493 11730
rect 17531 11696 17535 11730
rect 17535 11696 17565 11730
rect 17603 11696 17637 11730
rect 17675 11696 17705 11730
rect 17705 11696 17709 11730
rect 17747 11696 17773 11730
rect 17773 11696 17781 11730
rect 17819 11696 17841 11730
rect 17841 11696 17853 11730
rect 17891 11696 17909 11730
rect 17909 11696 17925 11730
rect 17963 11696 17977 11730
rect 17977 11696 17997 11730
rect 18035 11696 18045 11730
rect 18045 11696 18069 11730
rect 18538 14706 18572 14718
rect 18538 14684 18572 14706
rect 18538 14638 18572 14646
rect 18538 14612 18572 14638
rect 18538 14570 18572 14574
rect 18538 14540 18572 14570
rect 18538 14468 18572 14502
rect 18538 14400 18572 14430
rect 18538 14396 18572 14400
rect 18538 14332 18572 14358
rect 18538 14324 18572 14332
rect 18538 14264 18572 14286
rect 18538 14252 18572 14264
rect 19596 14706 19630 14718
rect 19596 14684 19630 14706
rect 19596 14638 19630 14646
rect 19596 14612 19630 14638
rect 19596 14570 19630 14574
rect 19596 14540 19630 14570
rect 19596 14468 19630 14502
rect 19596 14400 19630 14430
rect 19596 14396 19630 14400
rect 19596 14332 19630 14358
rect 19596 14324 19630 14332
rect 19596 14264 19630 14286
rect 19596 14252 19630 14264
rect 18538 14196 18572 14214
rect 18538 14180 18572 14196
rect 18538 14128 18572 14142
rect 18538 14108 18572 14128
rect 18538 14060 18572 14070
rect 18538 14036 18572 14060
rect 18538 13992 18572 13998
rect 18538 13964 18572 13992
rect 18538 13924 18572 13926
rect 18538 13892 18572 13924
rect 18538 13822 18572 13854
rect 18538 13820 18572 13822
rect 18538 13754 18572 13782
rect 18538 13748 18572 13754
rect 18538 13686 18572 13710
rect 18538 13676 18572 13686
rect 18538 13618 18572 13638
rect 18538 13604 18572 13618
rect 18538 13550 18572 13566
rect 18538 13532 18572 13550
rect 18538 13482 18572 13494
rect 18538 13460 18572 13482
rect 18538 13414 18572 13422
rect 18538 13388 18572 13414
rect 18538 13346 18572 13350
rect 18538 13316 18572 13346
rect 18538 13244 18572 13278
rect 18538 13176 18572 13206
rect 18538 13172 18572 13176
rect 18538 13108 18572 13134
rect 18538 13100 18572 13108
rect 18538 13040 18572 13062
rect 18538 13028 18572 13040
rect 18538 12972 18572 12990
rect 18538 12956 18572 12972
rect 18538 12904 18572 12918
rect 18538 12884 18572 12904
rect 18538 12836 18572 12846
rect 18538 12812 18572 12836
rect 18538 12768 18572 12774
rect 18538 12740 18572 12768
rect 18538 12700 18572 12702
rect 18538 12668 18572 12700
rect 18538 12598 18572 12630
rect 18538 12596 18572 12598
rect 18538 12530 18572 12558
rect 18538 12524 18572 12530
rect 18538 12462 18572 12486
rect 18538 12452 18572 12462
rect 18538 12394 18572 12414
rect 18538 12380 18572 12394
rect 18538 12326 18572 12342
rect 18538 12308 18572 12326
rect 18538 12258 18572 12270
rect 18538 12236 18572 12258
rect 18538 12190 18572 12198
rect 18538 12164 18572 12190
rect 18538 12122 18572 12126
rect 18538 12092 18572 12122
rect 18538 12020 18572 12054
rect 18538 11952 18572 11982
rect 18538 11948 18572 11952
rect 18538 11884 18572 11910
rect 18538 11876 18572 11884
rect 18538 11816 18572 11838
rect 18538 11804 18572 11816
rect 19596 14196 19630 14214
rect 19596 14180 19630 14196
rect 19596 14128 19630 14142
rect 19596 14108 19630 14128
rect 19596 14060 19630 14070
rect 19596 14036 19630 14060
rect 19596 13992 19630 13998
rect 19596 13964 19630 13992
rect 19596 13924 19630 13926
rect 19596 13892 19630 13924
rect 19596 13822 19630 13854
rect 19596 13820 19630 13822
rect 19596 13754 19630 13782
rect 19596 13748 19630 13754
rect 19596 13686 19630 13710
rect 19596 13676 19630 13686
rect 19596 13618 19630 13638
rect 19596 13604 19630 13618
rect 19596 13550 19630 13566
rect 19596 13532 19630 13550
rect 19596 13482 19630 13494
rect 19596 13460 19630 13482
rect 19596 13414 19630 13422
rect 19596 13388 19630 13414
rect 19596 13346 19630 13350
rect 19596 13316 19630 13346
rect 19596 13244 19630 13278
rect 19596 13176 19630 13206
rect 19596 13172 19630 13176
rect 19596 13108 19630 13134
rect 19596 13100 19630 13108
rect 19596 13040 19630 13062
rect 19596 13028 19630 13040
rect 19596 12972 19630 12990
rect 19596 12956 19630 12972
rect 19596 12904 19630 12918
rect 19596 12884 19630 12904
rect 19596 12836 19630 12846
rect 19596 12812 19630 12836
rect 19596 12768 19630 12774
rect 19596 12740 19630 12768
rect 19596 12700 19630 12702
rect 19596 12668 19630 12700
rect 19596 12598 19630 12630
rect 19596 12596 19630 12598
rect 19596 12530 19630 12558
rect 19596 12524 19630 12530
rect 19596 12462 19630 12486
rect 19596 12452 19630 12462
rect 19596 12394 19630 12414
rect 19596 12380 19630 12394
rect 19596 12326 19630 12342
rect 19596 12308 19630 12326
rect 19596 12258 19630 12270
rect 19596 12236 19630 12258
rect 19596 12190 19630 12198
rect 19596 12164 19630 12190
rect 19596 12122 19630 12126
rect 19596 12092 19630 12122
rect 19596 12020 19630 12054
rect 19596 11952 19630 11982
rect 19596 11948 19630 11952
rect 19596 11884 19630 11910
rect 19596 11876 19630 11884
rect 19596 11816 19630 11838
rect 19596 11804 19630 11816
rect 20530 14416 20564 14450
rect 20530 14344 20564 14378
rect 20530 14272 20564 14306
rect 20530 14200 20564 14234
rect 20530 14128 20564 14162
rect 18635 11680 18659 11714
rect 18659 11680 18669 11714
rect 18707 11680 18727 11714
rect 18727 11680 18741 11714
rect 18779 11680 18795 11714
rect 18795 11680 18813 11714
rect 18851 11680 18863 11714
rect 18863 11680 18885 11714
rect 18923 11680 18931 11714
rect 18931 11680 18957 11714
rect 18995 11680 18999 11714
rect 18999 11680 19029 11714
rect 19067 11680 19101 11714
rect 19139 11680 19169 11714
rect 19169 11680 19173 11714
rect 19211 11680 19237 11714
rect 19237 11680 19245 11714
rect 19283 11680 19305 11714
rect 19305 11680 19317 11714
rect 19355 11680 19373 11714
rect 19373 11680 19389 11714
rect 19427 11680 19441 11714
rect 19441 11680 19461 11714
rect 19499 11680 19509 11714
rect 19509 11680 19533 11714
rect 20530 14056 20564 14090
rect 20848 14416 20882 14450
rect 20848 14344 20882 14378
rect 20848 14272 20882 14306
rect 20848 14200 20882 14234
rect 20848 14128 20882 14162
rect 20848 14056 20882 14090
rect 21166 14416 21200 14450
rect 21166 14344 21200 14378
rect 21166 14272 21200 14306
rect 21166 14200 21200 14234
rect 21166 14128 21200 14162
rect 21166 14056 21200 14090
rect 21484 14416 21518 14450
rect 21484 14344 21518 14378
rect 21484 14272 21518 14306
rect 21484 14200 21518 14234
rect 21484 14128 21518 14162
rect 21484 14056 21518 14090
rect -8722 11202 -8720 11236
rect -8720 11202 -8688 11236
rect -8650 11202 -8618 11236
rect -8618 11202 -8616 11236
rect -8464 11202 -8462 11236
rect -8462 11202 -8430 11236
rect -8392 11202 -8360 11236
rect -8360 11202 -8358 11236
rect -8206 11202 -8204 11236
rect -8204 11202 -8172 11236
rect -8134 11202 -8102 11236
rect -8102 11202 -8100 11236
rect -7948 11202 -7946 11236
rect -7946 11202 -7914 11236
rect -7876 11202 -7844 11236
rect -7844 11202 -7842 11236
rect -7690 11202 -7688 11236
rect -7688 11202 -7656 11236
rect -7618 11202 -7586 11236
rect -7586 11202 -7584 11236
rect -7432 11202 -7430 11236
rect -7430 11202 -7398 11236
rect -7360 11202 -7328 11236
rect -7328 11202 -7326 11236
rect -7174 11202 -7172 11236
rect -7172 11202 -7140 11236
rect -7102 11202 -7070 11236
rect -7070 11202 -7068 11236
rect -6916 11202 -6914 11236
rect -6914 11202 -6882 11236
rect -6844 11202 -6812 11236
rect -6812 11202 -6810 11236
rect -6658 11202 -6656 11236
rect -6656 11202 -6624 11236
rect -6586 11202 -6554 11236
rect -6554 11202 -6552 11236
rect -6400 11202 -6398 11236
rect -6398 11202 -6366 11236
rect -6328 11202 -6296 11236
rect -6296 11202 -6294 11236
rect -6142 11202 -6140 11236
rect -6140 11202 -6108 11236
rect -6070 11202 -6038 11236
rect -6038 11202 -6036 11236
rect -5884 11202 -5882 11236
rect -5882 11202 -5850 11236
rect -5812 11202 -5780 11236
rect -5780 11202 -5778 11236
rect -5626 11202 -5624 11236
rect -5624 11202 -5592 11236
rect -5554 11202 -5522 11236
rect -5522 11202 -5520 11236
rect -5368 11202 -5366 11236
rect -5366 11202 -5334 11236
rect -5296 11202 -5264 11236
rect -5264 11202 -5262 11236
rect -5110 11202 -5108 11236
rect -5108 11202 -5076 11236
rect -5038 11202 -5006 11236
rect -5006 11202 -5004 11236
rect -4852 11202 -4850 11236
rect -4850 11202 -4818 11236
rect -4780 11202 -4748 11236
rect -4748 11202 -4746 11236
rect -4594 11202 -4592 11236
rect -4592 11202 -4560 11236
rect -4522 11202 -4490 11236
rect -4490 11202 -4488 11236
rect -4336 11202 -4334 11236
rect -4334 11202 -4302 11236
rect -4264 11202 -4232 11236
rect -4232 11202 -4230 11236
rect -4078 11202 -4076 11236
rect -4076 11202 -4044 11236
rect -4006 11202 -3974 11236
rect -3974 11202 -3972 11236
rect -3820 11202 -3818 11236
rect -3818 11202 -3786 11236
rect -3748 11202 -3716 11236
rect -3716 11202 -3714 11236
rect -8815 11123 -8781 11149
rect -8815 11115 -8781 11123
rect -8815 11055 -8781 11077
rect -8815 11043 -8781 11055
rect -8815 10987 -8781 11005
rect -8815 10971 -8781 10987
rect -8815 10919 -8781 10933
rect -8815 10899 -8781 10919
rect -8815 10851 -8781 10861
rect -8815 10827 -8781 10851
rect -8815 10783 -8781 10789
rect -8815 10755 -8781 10783
rect -8815 10715 -8781 10717
rect -8815 10683 -8781 10715
rect -8815 10613 -8781 10645
rect -8815 10611 -8781 10613
rect -8815 10545 -8781 10573
rect -8815 10539 -8781 10545
rect -8815 10477 -8781 10501
rect -8815 10467 -8781 10477
rect -8815 10409 -8781 10429
rect -8815 10395 -8781 10409
rect -8815 10341 -8781 10357
rect -8815 10323 -8781 10341
rect -8815 10273 -8781 10285
rect -8815 10251 -8781 10273
rect -8815 10205 -8781 10213
rect -8815 10179 -8781 10205
rect -8557 11123 -8523 11149
rect -8557 11115 -8523 11123
rect -8557 11055 -8523 11077
rect -8557 11043 -8523 11055
rect -8557 10987 -8523 11005
rect -8557 10971 -8523 10987
rect -8557 10919 -8523 10933
rect -8557 10899 -8523 10919
rect -8557 10851 -8523 10861
rect -8557 10827 -8523 10851
rect -8557 10783 -8523 10789
rect -8557 10755 -8523 10783
rect -8557 10715 -8523 10717
rect -8557 10683 -8523 10715
rect -8557 10613 -8523 10645
rect -8557 10611 -8523 10613
rect -8557 10545 -8523 10573
rect -8557 10539 -8523 10545
rect -8557 10477 -8523 10501
rect -8557 10467 -8523 10477
rect -8557 10409 -8523 10429
rect -8557 10395 -8523 10409
rect -8557 10341 -8523 10357
rect -8557 10323 -8523 10341
rect -8557 10273 -8523 10285
rect -8557 10251 -8523 10273
rect -8557 10205 -8523 10213
rect -8557 10179 -8523 10205
rect -8299 11123 -8265 11149
rect -8299 11115 -8265 11123
rect -8299 11055 -8265 11077
rect -8299 11043 -8265 11055
rect -8299 10987 -8265 11005
rect -8299 10971 -8265 10987
rect -8299 10919 -8265 10933
rect -8299 10899 -8265 10919
rect -8299 10851 -8265 10861
rect -8299 10827 -8265 10851
rect -8299 10783 -8265 10789
rect -8299 10755 -8265 10783
rect -8299 10715 -8265 10717
rect -8299 10683 -8265 10715
rect -8299 10613 -8265 10645
rect -8299 10611 -8265 10613
rect -8299 10545 -8265 10573
rect -8299 10539 -8265 10545
rect -8299 10477 -8265 10501
rect -8299 10467 -8265 10477
rect -8299 10409 -8265 10429
rect -8299 10395 -8265 10409
rect -8299 10341 -8265 10357
rect -8299 10323 -8265 10341
rect -8299 10273 -8265 10285
rect -8299 10251 -8265 10273
rect -8299 10205 -8265 10213
rect -8299 10179 -8265 10205
rect -8041 11123 -8007 11149
rect -8041 11115 -8007 11123
rect -8041 11055 -8007 11077
rect -8041 11043 -8007 11055
rect -8041 10987 -8007 11005
rect -8041 10971 -8007 10987
rect -8041 10919 -8007 10933
rect -8041 10899 -8007 10919
rect -8041 10851 -8007 10861
rect -8041 10827 -8007 10851
rect -8041 10783 -8007 10789
rect -8041 10755 -8007 10783
rect -8041 10715 -8007 10717
rect -8041 10683 -8007 10715
rect -8041 10613 -8007 10645
rect -8041 10611 -8007 10613
rect -8041 10545 -8007 10573
rect -8041 10539 -8007 10545
rect -8041 10477 -8007 10501
rect -8041 10467 -8007 10477
rect -8041 10409 -8007 10429
rect -8041 10395 -8007 10409
rect -8041 10341 -8007 10357
rect -8041 10323 -8007 10341
rect -8041 10273 -8007 10285
rect -8041 10251 -8007 10273
rect -8041 10205 -8007 10213
rect -8041 10179 -8007 10205
rect -7783 11123 -7749 11149
rect -7783 11115 -7749 11123
rect -7783 11055 -7749 11077
rect -7783 11043 -7749 11055
rect -7783 10987 -7749 11005
rect -7783 10971 -7749 10987
rect -7783 10919 -7749 10933
rect -7783 10899 -7749 10919
rect -7783 10851 -7749 10861
rect -7783 10827 -7749 10851
rect -7783 10783 -7749 10789
rect -7783 10755 -7749 10783
rect -7783 10715 -7749 10717
rect -7783 10683 -7749 10715
rect -7783 10613 -7749 10645
rect -7783 10611 -7749 10613
rect -7783 10545 -7749 10573
rect -7783 10539 -7749 10545
rect -7783 10477 -7749 10501
rect -7783 10467 -7749 10477
rect -7783 10409 -7749 10429
rect -7783 10395 -7749 10409
rect -7783 10341 -7749 10357
rect -7783 10323 -7749 10341
rect -7783 10273 -7749 10285
rect -7783 10251 -7749 10273
rect -7783 10205 -7749 10213
rect -7783 10179 -7749 10205
rect -7525 11123 -7491 11149
rect -7525 11115 -7491 11123
rect -7525 11055 -7491 11077
rect -7525 11043 -7491 11055
rect -7525 10987 -7491 11005
rect -7525 10971 -7491 10987
rect -7525 10919 -7491 10933
rect -7525 10899 -7491 10919
rect -7525 10851 -7491 10861
rect -7525 10827 -7491 10851
rect -7525 10783 -7491 10789
rect -7525 10755 -7491 10783
rect -7525 10715 -7491 10717
rect -7525 10683 -7491 10715
rect -7525 10613 -7491 10645
rect -7525 10611 -7491 10613
rect -7525 10545 -7491 10573
rect -7525 10539 -7491 10545
rect -7525 10477 -7491 10501
rect -7525 10467 -7491 10477
rect -7525 10409 -7491 10429
rect -7525 10395 -7491 10409
rect -7525 10341 -7491 10357
rect -7525 10323 -7491 10341
rect -7525 10273 -7491 10285
rect -7525 10251 -7491 10273
rect -7525 10205 -7491 10213
rect -7525 10179 -7491 10205
rect -7267 11123 -7233 11149
rect -7267 11115 -7233 11123
rect -7267 11055 -7233 11077
rect -7267 11043 -7233 11055
rect -7267 10987 -7233 11005
rect -7267 10971 -7233 10987
rect -7267 10919 -7233 10933
rect -7267 10899 -7233 10919
rect -7267 10851 -7233 10861
rect -7267 10827 -7233 10851
rect -7267 10783 -7233 10789
rect -7267 10755 -7233 10783
rect -7267 10715 -7233 10717
rect -7267 10683 -7233 10715
rect -7267 10613 -7233 10645
rect -7267 10611 -7233 10613
rect -7267 10545 -7233 10573
rect -7267 10539 -7233 10545
rect -7267 10477 -7233 10501
rect -7267 10467 -7233 10477
rect -7267 10409 -7233 10429
rect -7267 10395 -7233 10409
rect -7267 10341 -7233 10357
rect -7267 10323 -7233 10341
rect -7267 10273 -7233 10285
rect -7267 10251 -7233 10273
rect -7267 10205 -7233 10213
rect -7267 10179 -7233 10205
rect -7009 11123 -6975 11149
rect -7009 11115 -6975 11123
rect -7009 11055 -6975 11077
rect -7009 11043 -6975 11055
rect -7009 10987 -6975 11005
rect -7009 10971 -6975 10987
rect -7009 10919 -6975 10933
rect -7009 10899 -6975 10919
rect -7009 10851 -6975 10861
rect -7009 10827 -6975 10851
rect -7009 10783 -6975 10789
rect -7009 10755 -6975 10783
rect -7009 10715 -6975 10717
rect -7009 10683 -6975 10715
rect -7009 10613 -6975 10645
rect -7009 10611 -6975 10613
rect -7009 10545 -6975 10573
rect -7009 10539 -6975 10545
rect -7009 10477 -6975 10501
rect -7009 10467 -6975 10477
rect -7009 10409 -6975 10429
rect -7009 10395 -6975 10409
rect -7009 10341 -6975 10357
rect -7009 10323 -6975 10341
rect -7009 10273 -6975 10285
rect -7009 10251 -6975 10273
rect -7009 10205 -6975 10213
rect -7009 10179 -6975 10205
rect -6751 11123 -6717 11149
rect -6751 11115 -6717 11123
rect -6751 11055 -6717 11077
rect -6751 11043 -6717 11055
rect -6751 10987 -6717 11005
rect -6751 10971 -6717 10987
rect -6751 10919 -6717 10933
rect -6751 10899 -6717 10919
rect -6751 10851 -6717 10861
rect -6751 10827 -6717 10851
rect -6751 10783 -6717 10789
rect -6751 10755 -6717 10783
rect -6751 10715 -6717 10717
rect -6751 10683 -6717 10715
rect -6751 10613 -6717 10645
rect -6751 10611 -6717 10613
rect -6751 10545 -6717 10573
rect -6751 10539 -6717 10545
rect -6751 10477 -6717 10501
rect -6751 10467 -6717 10477
rect -6751 10409 -6717 10429
rect -6751 10395 -6717 10409
rect -6751 10341 -6717 10357
rect -6751 10323 -6717 10341
rect -6751 10273 -6717 10285
rect -6751 10251 -6717 10273
rect -6751 10205 -6717 10213
rect -6751 10179 -6717 10205
rect -6493 11123 -6459 11149
rect -6493 11115 -6459 11123
rect -6493 11055 -6459 11077
rect -6493 11043 -6459 11055
rect -6493 10987 -6459 11005
rect -6493 10971 -6459 10987
rect -6493 10919 -6459 10933
rect -6493 10899 -6459 10919
rect -6493 10851 -6459 10861
rect -6493 10827 -6459 10851
rect -6493 10783 -6459 10789
rect -6493 10755 -6459 10783
rect -6493 10715 -6459 10717
rect -6493 10683 -6459 10715
rect -6493 10613 -6459 10645
rect -6493 10611 -6459 10613
rect -6493 10545 -6459 10573
rect -6493 10539 -6459 10545
rect -6493 10477 -6459 10501
rect -6493 10467 -6459 10477
rect -6493 10409 -6459 10429
rect -6493 10395 -6459 10409
rect -6493 10341 -6459 10357
rect -6493 10323 -6459 10341
rect -6493 10273 -6459 10285
rect -6493 10251 -6459 10273
rect -6493 10205 -6459 10213
rect -6493 10179 -6459 10205
rect -6235 11123 -6201 11149
rect -6235 11115 -6201 11123
rect -6235 11055 -6201 11077
rect -6235 11043 -6201 11055
rect -6235 10987 -6201 11005
rect -6235 10971 -6201 10987
rect -6235 10919 -6201 10933
rect -6235 10899 -6201 10919
rect -6235 10851 -6201 10861
rect -6235 10827 -6201 10851
rect -6235 10783 -6201 10789
rect -6235 10755 -6201 10783
rect -6235 10715 -6201 10717
rect -6235 10683 -6201 10715
rect -6235 10613 -6201 10645
rect -6235 10611 -6201 10613
rect -6235 10545 -6201 10573
rect -6235 10539 -6201 10545
rect -6235 10477 -6201 10501
rect -6235 10467 -6201 10477
rect -6235 10409 -6201 10429
rect -6235 10395 -6201 10409
rect -6235 10341 -6201 10357
rect -6235 10323 -6201 10341
rect -6235 10273 -6201 10285
rect -6235 10251 -6201 10273
rect -6235 10205 -6201 10213
rect -6235 10179 -6201 10205
rect -5977 11123 -5943 11149
rect -5977 11115 -5943 11123
rect -5977 11055 -5943 11077
rect -5977 11043 -5943 11055
rect -5977 10987 -5943 11005
rect -5977 10971 -5943 10987
rect -5977 10919 -5943 10933
rect -5977 10899 -5943 10919
rect -5977 10851 -5943 10861
rect -5977 10827 -5943 10851
rect -5977 10783 -5943 10789
rect -5977 10755 -5943 10783
rect -5977 10715 -5943 10717
rect -5977 10683 -5943 10715
rect -5977 10613 -5943 10645
rect -5977 10611 -5943 10613
rect -5977 10545 -5943 10573
rect -5977 10539 -5943 10545
rect -5977 10477 -5943 10501
rect -5977 10467 -5943 10477
rect -5977 10409 -5943 10429
rect -5977 10395 -5943 10409
rect -5977 10341 -5943 10357
rect -5977 10323 -5943 10341
rect -5977 10273 -5943 10285
rect -5977 10251 -5943 10273
rect -5977 10205 -5943 10213
rect -5977 10179 -5943 10205
rect -5719 11123 -5685 11149
rect -5719 11115 -5685 11123
rect -5719 11055 -5685 11077
rect -5719 11043 -5685 11055
rect -5719 10987 -5685 11005
rect -5719 10971 -5685 10987
rect -5719 10919 -5685 10933
rect -5719 10899 -5685 10919
rect -5719 10851 -5685 10861
rect -5719 10827 -5685 10851
rect -5719 10783 -5685 10789
rect -5719 10755 -5685 10783
rect -5719 10715 -5685 10717
rect -5719 10683 -5685 10715
rect -5719 10613 -5685 10645
rect -5719 10611 -5685 10613
rect -5719 10545 -5685 10573
rect -5719 10539 -5685 10545
rect -5719 10477 -5685 10501
rect -5719 10467 -5685 10477
rect -5719 10409 -5685 10429
rect -5719 10395 -5685 10409
rect -5719 10341 -5685 10357
rect -5719 10323 -5685 10341
rect -5719 10273 -5685 10285
rect -5719 10251 -5685 10273
rect -5719 10205 -5685 10213
rect -5719 10179 -5685 10205
rect -5461 11123 -5427 11149
rect -5461 11115 -5427 11123
rect -5461 11055 -5427 11077
rect -5461 11043 -5427 11055
rect -5461 10987 -5427 11005
rect -5461 10971 -5427 10987
rect -5461 10919 -5427 10933
rect -5461 10899 -5427 10919
rect -5461 10851 -5427 10861
rect -5461 10827 -5427 10851
rect -5461 10783 -5427 10789
rect -5461 10755 -5427 10783
rect -5461 10715 -5427 10717
rect -5461 10683 -5427 10715
rect -5461 10613 -5427 10645
rect -5461 10611 -5427 10613
rect -5461 10545 -5427 10573
rect -5461 10539 -5427 10545
rect -5461 10477 -5427 10501
rect -5461 10467 -5427 10477
rect -5461 10409 -5427 10429
rect -5461 10395 -5427 10409
rect -5461 10341 -5427 10357
rect -5461 10323 -5427 10341
rect -5461 10273 -5427 10285
rect -5461 10251 -5427 10273
rect -5461 10205 -5427 10213
rect -5461 10179 -5427 10205
rect -5203 11123 -5169 11149
rect -5203 11115 -5169 11123
rect -5203 11055 -5169 11077
rect -5203 11043 -5169 11055
rect -5203 10987 -5169 11005
rect -5203 10971 -5169 10987
rect -5203 10919 -5169 10933
rect -5203 10899 -5169 10919
rect -5203 10851 -5169 10861
rect -5203 10827 -5169 10851
rect -5203 10783 -5169 10789
rect -5203 10755 -5169 10783
rect -5203 10715 -5169 10717
rect -5203 10683 -5169 10715
rect -5203 10613 -5169 10645
rect -5203 10611 -5169 10613
rect -5203 10545 -5169 10573
rect -5203 10539 -5169 10545
rect -5203 10477 -5169 10501
rect -5203 10467 -5169 10477
rect -5203 10409 -5169 10429
rect -5203 10395 -5169 10409
rect -5203 10341 -5169 10357
rect -5203 10323 -5169 10341
rect -5203 10273 -5169 10285
rect -5203 10251 -5169 10273
rect -5203 10205 -5169 10213
rect -5203 10179 -5169 10205
rect -4945 11123 -4911 11149
rect -4945 11115 -4911 11123
rect -4945 11055 -4911 11077
rect -4945 11043 -4911 11055
rect -4945 10987 -4911 11005
rect -4945 10971 -4911 10987
rect -4945 10919 -4911 10933
rect -4945 10899 -4911 10919
rect -4945 10851 -4911 10861
rect -4945 10827 -4911 10851
rect -4945 10783 -4911 10789
rect -4945 10755 -4911 10783
rect -4945 10715 -4911 10717
rect -4945 10683 -4911 10715
rect -4945 10613 -4911 10645
rect -4945 10611 -4911 10613
rect -4945 10545 -4911 10573
rect -4945 10539 -4911 10545
rect -4945 10477 -4911 10501
rect -4945 10467 -4911 10477
rect -4945 10409 -4911 10429
rect -4945 10395 -4911 10409
rect -4945 10341 -4911 10357
rect -4945 10323 -4911 10341
rect -4945 10273 -4911 10285
rect -4945 10251 -4911 10273
rect -4945 10205 -4911 10213
rect -4945 10179 -4911 10205
rect -4687 11123 -4653 11149
rect -4687 11115 -4653 11123
rect -4687 11055 -4653 11077
rect -4687 11043 -4653 11055
rect -4687 10987 -4653 11005
rect -4687 10971 -4653 10987
rect -4687 10919 -4653 10933
rect -4687 10899 -4653 10919
rect -4687 10851 -4653 10861
rect -4687 10827 -4653 10851
rect -4687 10783 -4653 10789
rect -4687 10755 -4653 10783
rect -4687 10715 -4653 10717
rect -4687 10683 -4653 10715
rect -4687 10613 -4653 10645
rect -4687 10611 -4653 10613
rect -4687 10545 -4653 10573
rect -4687 10539 -4653 10545
rect -4687 10477 -4653 10501
rect -4687 10467 -4653 10477
rect -4687 10409 -4653 10429
rect -4687 10395 -4653 10409
rect -4687 10341 -4653 10357
rect -4687 10323 -4653 10341
rect -4687 10273 -4653 10285
rect -4687 10251 -4653 10273
rect -4687 10205 -4653 10213
rect -4687 10179 -4653 10205
rect -4429 11123 -4395 11149
rect -4429 11115 -4395 11123
rect -4429 11055 -4395 11077
rect -4429 11043 -4395 11055
rect -4429 10987 -4395 11005
rect -4429 10971 -4395 10987
rect -4429 10919 -4395 10933
rect -4429 10899 -4395 10919
rect -4429 10851 -4395 10861
rect -4429 10827 -4395 10851
rect -4429 10783 -4395 10789
rect -4429 10755 -4395 10783
rect -4429 10715 -4395 10717
rect -4429 10683 -4395 10715
rect -4429 10613 -4395 10645
rect -4429 10611 -4395 10613
rect -4429 10545 -4395 10573
rect -4429 10539 -4395 10545
rect -4429 10477 -4395 10501
rect -4429 10467 -4395 10477
rect -4429 10409 -4395 10429
rect -4429 10395 -4395 10409
rect -4429 10341 -4395 10357
rect -4429 10323 -4395 10341
rect -4429 10273 -4395 10285
rect -4429 10251 -4395 10273
rect -4429 10205 -4395 10213
rect -4429 10179 -4395 10205
rect -4171 11123 -4137 11149
rect -4171 11115 -4137 11123
rect -4171 11055 -4137 11077
rect -4171 11043 -4137 11055
rect -4171 10987 -4137 11005
rect -4171 10971 -4137 10987
rect -4171 10919 -4137 10933
rect -4171 10899 -4137 10919
rect -4171 10851 -4137 10861
rect -4171 10827 -4137 10851
rect -4171 10783 -4137 10789
rect -4171 10755 -4137 10783
rect -4171 10715 -4137 10717
rect -4171 10683 -4137 10715
rect -4171 10613 -4137 10645
rect -4171 10611 -4137 10613
rect -4171 10545 -4137 10573
rect -4171 10539 -4137 10545
rect -4171 10477 -4137 10501
rect -4171 10467 -4137 10477
rect -4171 10409 -4137 10429
rect -4171 10395 -4137 10409
rect -4171 10341 -4137 10357
rect -4171 10323 -4137 10341
rect -4171 10273 -4137 10285
rect -4171 10251 -4137 10273
rect -4171 10205 -4137 10213
rect -4171 10179 -4137 10205
rect -3913 11123 -3879 11149
rect -3913 11115 -3879 11123
rect -3913 11055 -3879 11077
rect -3913 11043 -3879 11055
rect -3913 10987 -3879 11005
rect -3913 10971 -3879 10987
rect -3913 10919 -3879 10933
rect -3913 10899 -3879 10919
rect -3913 10851 -3879 10861
rect -3913 10827 -3879 10851
rect -3913 10783 -3879 10789
rect -3913 10755 -3879 10783
rect -3913 10715 -3879 10717
rect -3913 10683 -3879 10715
rect -3913 10613 -3879 10645
rect -3913 10611 -3879 10613
rect -3913 10545 -3879 10573
rect -3913 10539 -3879 10545
rect -3913 10477 -3879 10501
rect -3913 10467 -3879 10477
rect -3913 10409 -3879 10429
rect -3913 10395 -3879 10409
rect -3913 10341 -3879 10357
rect -3913 10323 -3879 10341
rect -3913 10273 -3879 10285
rect -3913 10251 -3879 10273
rect -3913 10205 -3879 10213
rect -3913 10179 -3879 10205
rect -3655 11123 -3621 11149
rect -3655 11115 -3621 11123
rect -3655 11055 -3621 11077
rect -3655 11043 -3621 11055
rect -3655 10987 -3621 11005
rect -3655 10971 -3621 10987
rect -3655 10919 -3621 10933
rect -3655 10899 -3621 10919
rect -3655 10851 -3621 10861
rect -3655 10827 -3621 10851
rect -3655 10783 -3621 10789
rect -3655 10755 -3621 10783
rect -3655 10715 -3621 10717
rect -3655 10683 -3621 10715
rect -3655 10613 -3621 10645
rect -3655 10611 -3621 10613
rect -3655 10545 -3621 10573
rect -3655 10539 -3621 10545
rect -3655 10477 -3621 10501
rect -3655 10467 -3621 10477
rect -3655 10409 -3621 10429
rect -3655 10395 -3621 10409
rect -3655 10341 -3621 10357
rect -3655 10323 -3621 10341
rect -3655 10273 -3621 10285
rect -3655 10251 -3621 10273
rect -3655 10205 -3621 10213
rect -3655 10179 -3621 10205
rect -8722 10092 -8720 10126
rect -8720 10092 -8688 10126
rect -8650 10092 -8618 10126
rect -8618 10092 -8616 10126
rect -8464 10092 -8462 10126
rect -8462 10092 -8430 10126
rect -8392 10092 -8360 10126
rect -8360 10092 -8358 10126
rect -8206 10092 -8204 10126
rect -8204 10092 -8172 10126
rect -8134 10092 -8102 10126
rect -8102 10092 -8100 10126
rect -7948 10092 -7946 10126
rect -7946 10092 -7914 10126
rect -7876 10092 -7844 10126
rect -7844 10092 -7842 10126
rect -7690 10092 -7688 10126
rect -7688 10092 -7656 10126
rect -7618 10092 -7586 10126
rect -7586 10092 -7584 10126
rect -7432 10092 -7430 10126
rect -7430 10092 -7398 10126
rect -7360 10092 -7328 10126
rect -7328 10092 -7326 10126
rect -7174 10092 -7172 10126
rect -7172 10092 -7140 10126
rect -7102 10092 -7070 10126
rect -7070 10092 -7068 10126
rect -6916 10092 -6914 10126
rect -6914 10092 -6882 10126
rect -6844 10092 -6812 10126
rect -6812 10092 -6810 10126
rect -6658 10092 -6656 10126
rect -6656 10092 -6624 10126
rect -6586 10092 -6554 10126
rect -6554 10092 -6552 10126
rect -6400 10092 -6398 10126
rect -6398 10092 -6366 10126
rect -6328 10092 -6296 10126
rect -6296 10092 -6294 10126
rect -6142 10092 -6140 10126
rect -6140 10092 -6108 10126
rect -6070 10092 -6038 10126
rect -6038 10092 -6036 10126
rect -5884 10092 -5882 10126
rect -5882 10092 -5850 10126
rect -5812 10092 -5780 10126
rect -5780 10092 -5778 10126
rect -5626 10092 -5624 10126
rect -5624 10092 -5592 10126
rect -5554 10092 -5522 10126
rect -5522 10092 -5520 10126
rect -5368 10092 -5366 10126
rect -5366 10092 -5334 10126
rect -5296 10092 -5264 10126
rect -5264 10092 -5262 10126
rect -5110 10092 -5108 10126
rect -5108 10092 -5076 10126
rect -5038 10092 -5006 10126
rect -5006 10092 -5004 10126
rect -4852 10092 -4850 10126
rect -4850 10092 -4818 10126
rect -4780 10092 -4748 10126
rect -4748 10092 -4746 10126
rect -4594 10092 -4592 10126
rect -4592 10092 -4560 10126
rect -4522 10092 -4490 10126
rect -4490 10092 -4488 10126
rect -4336 10092 -4334 10126
rect -4334 10092 -4302 10126
rect -4264 10092 -4232 10126
rect -4232 10092 -4230 10126
rect -4078 10092 -4076 10126
rect -4076 10092 -4044 10126
rect -4006 10092 -3974 10126
rect -3974 10092 -3972 10126
rect -3820 10092 -3818 10126
rect -3818 10092 -3786 10126
rect -3748 10092 -3716 10126
rect -3716 10092 -3714 10126
rect -7687 9837 -7685 9871
rect -7685 9837 -7653 9871
rect -7615 9837 -7583 9871
rect -7583 9837 -7581 9871
rect -7221 9837 -7219 9871
rect -7219 9837 -7187 9871
rect -7149 9837 -7117 9871
rect -7117 9837 -7115 9871
rect -6963 9837 -6961 9871
rect -6961 9837 -6929 9871
rect -6891 9837 -6859 9871
rect -6859 9837 -6857 9871
rect -6705 9837 -6703 9871
rect -6703 9837 -6671 9871
rect -6633 9837 -6601 9871
rect -6601 9837 -6599 9871
rect -6447 9837 -6445 9871
rect -6445 9837 -6413 9871
rect -6375 9837 -6343 9871
rect -6343 9837 -6341 9871
rect -6189 9837 -6187 9871
rect -6187 9837 -6155 9871
rect -6117 9837 -6085 9871
rect -6085 9837 -6083 9871
rect -5931 9837 -5929 9871
rect -5929 9837 -5897 9871
rect -5859 9837 -5827 9871
rect -5827 9837 -5825 9871
rect -5673 9837 -5671 9871
rect -5671 9837 -5639 9871
rect -5601 9837 -5569 9871
rect -5569 9837 -5567 9871
rect -5415 9837 -5413 9871
rect -5413 9837 -5381 9871
rect -5343 9837 -5311 9871
rect -5311 9837 -5309 9871
rect -5157 9837 -5155 9871
rect -5155 9837 -5123 9871
rect -5085 9837 -5053 9871
rect -5053 9837 -5051 9871
rect -4899 9837 -4897 9871
rect -4897 9837 -4865 9871
rect -4827 9837 -4795 9871
rect -4795 9837 -4793 9871
rect -7780 9758 -7746 9784
rect -7780 9750 -7746 9758
rect -7780 9690 -7746 9712
rect -7780 9678 -7746 9690
rect -7780 9622 -7746 9640
rect -7780 9606 -7746 9622
rect -7780 9554 -7746 9568
rect -7780 9534 -7746 9554
rect -7780 9486 -7746 9496
rect -7780 9462 -7746 9486
rect -7780 9418 -7746 9424
rect -7780 9390 -7746 9418
rect -7780 9350 -7746 9352
rect -7780 9318 -7746 9350
rect -7780 9248 -7746 9280
rect -7780 9246 -7746 9248
rect -7780 9180 -7746 9208
rect -7780 9174 -7746 9180
rect -7780 9112 -7746 9136
rect -7780 9102 -7746 9112
rect -7780 9044 -7746 9064
rect -7780 9030 -7746 9044
rect -7780 8976 -7746 8992
rect -7780 8958 -7746 8976
rect -7780 8908 -7746 8920
rect -7780 8886 -7746 8908
rect -7780 8840 -7746 8848
rect -7780 8814 -7746 8840
rect -7522 9758 -7488 9784
rect -7522 9750 -7488 9758
rect -7522 9690 -7488 9712
rect -7522 9678 -7488 9690
rect -7522 9622 -7488 9640
rect -7522 9606 -7488 9622
rect -7522 9554 -7488 9568
rect -7522 9534 -7488 9554
rect -7522 9486 -7488 9496
rect -7522 9462 -7488 9486
rect -7522 9418 -7488 9424
rect -7522 9390 -7488 9418
rect -7522 9350 -7488 9352
rect -7522 9318 -7488 9350
rect -7522 9248 -7488 9280
rect -7522 9246 -7488 9248
rect -7522 9180 -7488 9208
rect -7522 9174 -7488 9180
rect -7522 9112 -7488 9136
rect -7522 9102 -7488 9112
rect -7522 9044 -7488 9064
rect -7522 9030 -7488 9044
rect -7522 8976 -7488 8992
rect -7522 8958 -7488 8976
rect -7522 8908 -7488 8920
rect -7522 8886 -7488 8908
rect -7522 8840 -7488 8848
rect -7522 8814 -7488 8840
rect -7314 9758 -7280 9784
rect -7314 9750 -7280 9758
rect -7314 9690 -7280 9712
rect -7314 9678 -7280 9690
rect -7314 9622 -7280 9640
rect -7314 9606 -7280 9622
rect -7314 9554 -7280 9568
rect -7314 9534 -7280 9554
rect -7314 9486 -7280 9496
rect -7314 9462 -7280 9486
rect -7314 9418 -7280 9424
rect -7314 9390 -7280 9418
rect -7314 9350 -7280 9352
rect -7314 9318 -7280 9350
rect -7314 9248 -7280 9280
rect -7314 9246 -7280 9248
rect -7314 9180 -7280 9208
rect -7314 9174 -7280 9180
rect -7314 9112 -7280 9136
rect -7314 9102 -7280 9112
rect -7314 9044 -7280 9064
rect -7314 9030 -7280 9044
rect -7314 8976 -7280 8992
rect -7314 8958 -7280 8976
rect -7314 8908 -7280 8920
rect -7314 8886 -7280 8908
rect -7314 8840 -7280 8848
rect -7314 8814 -7280 8840
rect -7056 9758 -7022 9784
rect -7056 9750 -7022 9758
rect -7056 9690 -7022 9712
rect -7056 9678 -7022 9690
rect -7056 9622 -7022 9640
rect -7056 9606 -7022 9622
rect -7056 9554 -7022 9568
rect -7056 9534 -7022 9554
rect -7056 9486 -7022 9496
rect -7056 9462 -7022 9486
rect -7056 9418 -7022 9424
rect -7056 9390 -7022 9418
rect -7056 9350 -7022 9352
rect -7056 9318 -7022 9350
rect -7056 9248 -7022 9280
rect -7056 9246 -7022 9248
rect -7056 9180 -7022 9208
rect -7056 9174 -7022 9180
rect -7056 9112 -7022 9136
rect -7056 9102 -7022 9112
rect -7056 9044 -7022 9064
rect -7056 9030 -7022 9044
rect -7056 8976 -7022 8992
rect -7056 8958 -7022 8976
rect -7056 8908 -7022 8920
rect -7056 8886 -7022 8908
rect -7056 8840 -7022 8848
rect -7056 8814 -7022 8840
rect -6798 9758 -6764 9784
rect -6798 9750 -6764 9758
rect -6798 9690 -6764 9712
rect -6798 9678 -6764 9690
rect -6798 9622 -6764 9640
rect -6798 9606 -6764 9622
rect -6798 9554 -6764 9568
rect -6798 9534 -6764 9554
rect -6798 9486 -6764 9496
rect -6798 9462 -6764 9486
rect -6798 9418 -6764 9424
rect -6798 9390 -6764 9418
rect -6798 9350 -6764 9352
rect -6798 9318 -6764 9350
rect -6798 9248 -6764 9280
rect -6798 9246 -6764 9248
rect -6798 9180 -6764 9208
rect -6798 9174 -6764 9180
rect -6798 9112 -6764 9136
rect -6798 9102 -6764 9112
rect -6798 9044 -6764 9064
rect -6798 9030 -6764 9044
rect -6798 8976 -6764 8992
rect -6798 8958 -6764 8976
rect -6798 8908 -6764 8920
rect -6798 8886 -6764 8908
rect -6798 8840 -6764 8848
rect -6798 8814 -6764 8840
rect -6540 9758 -6506 9784
rect -6540 9750 -6506 9758
rect -6540 9690 -6506 9712
rect -6540 9678 -6506 9690
rect -6540 9622 -6506 9640
rect -6540 9606 -6506 9622
rect -6540 9554 -6506 9568
rect -6540 9534 -6506 9554
rect -6540 9486 -6506 9496
rect -6540 9462 -6506 9486
rect -6540 9418 -6506 9424
rect -6540 9390 -6506 9418
rect -6540 9350 -6506 9352
rect -6540 9318 -6506 9350
rect -6540 9248 -6506 9280
rect -6540 9246 -6506 9248
rect -6540 9180 -6506 9208
rect -6540 9174 -6506 9180
rect -6540 9112 -6506 9136
rect -6540 9102 -6506 9112
rect -6540 9044 -6506 9064
rect -6540 9030 -6506 9044
rect -6540 8976 -6506 8992
rect -6540 8958 -6506 8976
rect -6540 8908 -6506 8920
rect -6540 8886 -6506 8908
rect -6540 8840 -6506 8848
rect -6540 8814 -6506 8840
rect -6282 9758 -6248 9784
rect -6282 9750 -6248 9758
rect -6282 9690 -6248 9712
rect -6282 9678 -6248 9690
rect -6282 9622 -6248 9640
rect -6282 9606 -6248 9622
rect -6282 9554 -6248 9568
rect -6282 9534 -6248 9554
rect -6282 9486 -6248 9496
rect -6282 9462 -6248 9486
rect -6282 9418 -6248 9424
rect -6282 9390 -6248 9418
rect -6282 9350 -6248 9352
rect -6282 9318 -6248 9350
rect -6282 9248 -6248 9280
rect -6282 9246 -6248 9248
rect -6282 9180 -6248 9208
rect -6282 9174 -6248 9180
rect -6282 9112 -6248 9136
rect -6282 9102 -6248 9112
rect -6282 9044 -6248 9064
rect -6282 9030 -6248 9044
rect -6282 8976 -6248 8992
rect -6282 8958 -6248 8976
rect -6282 8908 -6248 8920
rect -6282 8886 -6248 8908
rect -6282 8840 -6248 8848
rect -6282 8814 -6248 8840
rect -6024 9758 -5990 9784
rect -6024 9750 -5990 9758
rect -6024 9690 -5990 9712
rect -6024 9678 -5990 9690
rect -6024 9622 -5990 9640
rect -6024 9606 -5990 9622
rect -6024 9554 -5990 9568
rect -6024 9534 -5990 9554
rect -6024 9486 -5990 9496
rect -6024 9462 -5990 9486
rect -6024 9418 -5990 9424
rect -6024 9390 -5990 9418
rect -6024 9350 -5990 9352
rect -6024 9318 -5990 9350
rect -6024 9248 -5990 9280
rect -6024 9246 -5990 9248
rect -6024 9180 -5990 9208
rect -6024 9174 -5990 9180
rect -6024 9112 -5990 9136
rect -6024 9102 -5990 9112
rect -6024 9044 -5990 9064
rect -6024 9030 -5990 9044
rect -6024 8976 -5990 8992
rect -6024 8958 -5990 8976
rect -6024 8908 -5990 8920
rect -6024 8886 -5990 8908
rect -6024 8840 -5990 8848
rect -6024 8814 -5990 8840
rect -5766 9758 -5732 9784
rect -5766 9750 -5732 9758
rect -5766 9690 -5732 9712
rect -5766 9678 -5732 9690
rect -5766 9622 -5732 9640
rect -5766 9606 -5732 9622
rect -5766 9554 -5732 9568
rect -5766 9534 -5732 9554
rect -5766 9486 -5732 9496
rect -5766 9462 -5732 9486
rect -5766 9418 -5732 9424
rect -5766 9390 -5732 9418
rect -5766 9350 -5732 9352
rect -5766 9318 -5732 9350
rect -5766 9248 -5732 9280
rect -5766 9246 -5732 9248
rect -5766 9180 -5732 9208
rect -5766 9174 -5732 9180
rect -5766 9112 -5732 9136
rect -5766 9102 -5732 9112
rect -5766 9044 -5732 9064
rect -5766 9030 -5732 9044
rect -5766 8976 -5732 8992
rect -5766 8958 -5732 8976
rect -5766 8908 -5732 8920
rect -5766 8886 -5732 8908
rect -5766 8840 -5732 8848
rect -5766 8814 -5732 8840
rect -5508 9758 -5474 9784
rect -5508 9750 -5474 9758
rect -5508 9690 -5474 9712
rect -5508 9678 -5474 9690
rect -5508 9622 -5474 9640
rect -5508 9606 -5474 9622
rect -5508 9554 -5474 9568
rect -5508 9534 -5474 9554
rect -5508 9486 -5474 9496
rect -5508 9462 -5474 9486
rect -5508 9418 -5474 9424
rect -5508 9390 -5474 9418
rect -5508 9350 -5474 9352
rect -5508 9318 -5474 9350
rect -5508 9248 -5474 9280
rect -5508 9246 -5474 9248
rect -5508 9180 -5474 9208
rect -5508 9174 -5474 9180
rect -5508 9112 -5474 9136
rect -5508 9102 -5474 9112
rect -5508 9044 -5474 9064
rect -5508 9030 -5474 9044
rect -5508 8976 -5474 8992
rect -5508 8958 -5474 8976
rect -5508 8908 -5474 8920
rect -5508 8886 -5474 8908
rect -5508 8840 -5474 8848
rect -5508 8814 -5474 8840
rect -5250 9758 -5216 9784
rect -5250 9750 -5216 9758
rect -5250 9690 -5216 9712
rect -5250 9678 -5216 9690
rect -5250 9622 -5216 9640
rect -5250 9606 -5216 9622
rect -5250 9554 -5216 9568
rect -5250 9534 -5216 9554
rect -5250 9486 -5216 9496
rect -5250 9462 -5216 9486
rect -5250 9418 -5216 9424
rect -5250 9390 -5216 9418
rect -5250 9350 -5216 9352
rect -5250 9318 -5216 9350
rect -5250 9248 -5216 9280
rect -5250 9246 -5216 9248
rect -5250 9180 -5216 9208
rect -5250 9174 -5216 9180
rect -5250 9112 -5216 9136
rect -5250 9102 -5216 9112
rect -5250 9044 -5216 9064
rect -5250 9030 -5216 9044
rect -5250 8976 -5216 8992
rect -5250 8958 -5216 8976
rect -5250 8908 -5216 8920
rect -5250 8886 -5216 8908
rect -5250 8840 -5216 8848
rect -5250 8814 -5216 8840
rect -4992 9758 -4958 9784
rect -4992 9750 -4958 9758
rect -4992 9690 -4958 9712
rect -4992 9678 -4958 9690
rect -4992 9622 -4958 9640
rect -4992 9606 -4958 9622
rect -4992 9554 -4958 9568
rect -4992 9534 -4958 9554
rect -4992 9486 -4958 9496
rect -4992 9462 -4958 9486
rect -4992 9418 -4958 9424
rect -4992 9390 -4958 9418
rect -4992 9350 -4958 9352
rect -4992 9318 -4958 9350
rect -4992 9248 -4958 9280
rect -4992 9246 -4958 9248
rect -4992 9180 -4958 9208
rect -4992 9174 -4958 9180
rect -4992 9112 -4958 9136
rect -4992 9102 -4958 9112
rect -4992 9044 -4958 9064
rect -4992 9030 -4958 9044
rect -4992 8976 -4958 8992
rect -4992 8958 -4958 8976
rect -4992 8908 -4958 8920
rect -4992 8886 -4958 8908
rect -4992 8840 -4958 8848
rect -4992 8814 -4958 8840
rect -4734 9758 -4700 9784
rect -4734 9750 -4700 9758
rect -4734 9690 -4700 9712
rect -4734 9678 -4700 9690
rect -4734 9622 -4700 9640
rect -4734 9606 -4700 9622
rect -4734 9554 -4700 9568
rect -4734 9534 -4700 9554
rect -4734 9486 -4700 9496
rect -4734 9462 -4700 9486
rect -4734 9418 -4700 9424
rect -4734 9390 -4700 9418
rect -4734 9350 -4700 9352
rect -4734 9318 -4700 9350
rect -4734 9248 -4700 9280
rect -4734 9246 -4700 9248
rect -4734 9180 -4700 9208
rect -4734 9174 -4700 9180
rect -4734 9112 -4700 9136
rect -4734 9102 -4700 9112
rect -4734 9044 -4700 9064
rect -4734 9030 -4700 9044
rect -4734 8976 -4700 8992
rect -4734 8958 -4700 8976
rect -4734 8908 -4700 8920
rect -4734 8886 -4700 8908
rect -4734 8840 -4700 8848
rect -4734 8814 -4700 8840
rect -7687 8727 -7685 8761
rect -7685 8727 -7653 8761
rect -7615 8727 -7583 8761
rect -7583 8727 -7581 8761
rect -7221 8727 -7219 8761
rect -7219 8727 -7187 8761
rect -7149 8727 -7117 8761
rect -7117 8727 -7115 8761
rect -6963 8727 -6961 8761
rect -6961 8727 -6929 8761
rect -6891 8727 -6859 8761
rect -6859 8727 -6857 8761
rect -6705 8727 -6703 8761
rect -6703 8727 -6671 8761
rect -6633 8727 -6601 8761
rect -6601 8727 -6599 8761
rect -6447 8727 -6445 8761
rect -6445 8727 -6413 8761
rect -6375 8727 -6343 8761
rect -6343 8727 -6341 8761
rect -6189 8727 -6187 8761
rect -6187 8727 -6155 8761
rect -6117 8727 -6085 8761
rect -6085 8727 -6083 8761
rect -5931 8727 -5929 8761
rect -5929 8727 -5897 8761
rect -5859 8727 -5827 8761
rect -5827 8727 -5825 8761
rect -5673 8727 -5671 8761
rect -5671 8727 -5639 8761
rect -5601 8727 -5569 8761
rect -5569 8727 -5567 8761
rect -5415 8727 -5413 8761
rect -5413 8727 -5381 8761
rect -5343 8727 -5311 8761
rect -5311 8727 -5309 8761
rect -5157 8727 -5155 8761
rect -5155 8727 -5123 8761
rect -5085 8727 -5053 8761
rect -5053 8727 -5051 8761
rect -4899 8727 -4897 8761
rect -4897 8727 -4865 8761
rect -4827 8727 -4795 8761
rect -4795 8727 -4793 8761
rect 13152 10944 13174 10950
rect 13174 10944 13186 10950
rect 13252 10944 13264 10950
rect 13264 10944 13286 10950
rect 13352 10944 13354 10950
rect 13354 10944 13386 10950
rect 13152 10916 13186 10944
rect 13252 10916 13286 10944
rect 13352 10916 13386 10944
rect 13452 10916 13486 10950
rect 13552 10916 13586 10950
rect 13652 10944 13680 10950
rect 13680 10944 13686 10950
rect 13652 10916 13686 10944
rect 13152 10816 13186 10850
rect 13252 10816 13286 10850
rect 13352 10816 13386 10850
rect 13452 10816 13486 10850
rect 13552 10816 13586 10850
rect 13652 10816 13686 10850
rect 13152 10716 13186 10750
rect 13252 10716 13286 10750
rect 13352 10716 13386 10750
rect 13452 10716 13486 10750
rect 13552 10716 13586 10750
rect 13652 10716 13686 10750
rect 13152 10618 13186 10650
rect 13252 10618 13286 10650
rect 13352 10618 13386 10650
rect 13152 10616 13174 10618
rect 13174 10616 13186 10618
rect 13252 10616 13264 10618
rect 13264 10616 13286 10618
rect 13352 10616 13354 10618
rect 13354 10616 13386 10618
rect 13452 10616 13486 10650
rect 13552 10616 13586 10650
rect 13652 10618 13686 10650
rect 13652 10616 13680 10618
rect 13680 10616 13686 10618
rect 13152 10528 13186 10550
rect 13252 10528 13286 10550
rect 13352 10528 13386 10550
rect 13152 10516 13174 10528
rect 13174 10516 13186 10528
rect 13252 10516 13264 10528
rect 13264 10516 13286 10528
rect 13352 10516 13354 10528
rect 13354 10516 13386 10528
rect 13452 10516 13486 10550
rect 13552 10516 13586 10550
rect 13652 10528 13686 10550
rect 13652 10516 13680 10528
rect 13680 10516 13686 10528
rect 13152 10438 13186 10450
rect 13252 10438 13286 10450
rect 13352 10438 13386 10450
rect 13152 10416 13174 10438
rect 13174 10416 13186 10438
rect 13252 10416 13264 10438
rect 13264 10416 13286 10438
rect 13352 10416 13354 10438
rect 13354 10416 13386 10438
rect 13452 10416 13486 10450
rect 13552 10416 13586 10450
rect 13652 10438 13686 10450
rect 13652 10416 13680 10438
rect 13680 10416 13686 10438
rect 15051 11294 15075 11328
rect 15075 11294 15085 11328
rect 15123 11294 15143 11328
rect 15143 11294 15157 11328
rect 15195 11294 15211 11328
rect 15211 11294 15229 11328
rect 15267 11294 15279 11328
rect 15279 11294 15301 11328
rect 15339 11294 15347 11328
rect 15347 11294 15373 11328
rect 15411 11294 15415 11328
rect 15415 11294 15445 11328
rect 15483 11294 15517 11328
rect 15555 11294 15585 11328
rect 15585 11294 15589 11328
rect 15627 11294 15653 11328
rect 15653 11294 15661 11328
rect 15699 11294 15721 11328
rect 15721 11294 15733 11328
rect 15771 11294 15789 11328
rect 15789 11294 15805 11328
rect 15843 11294 15857 11328
rect 15857 11294 15877 11328
rect 15915 11294 15925 11328
rect 15925 11294 15949 11328
rect 16109 11294 16133 11328
rect 16133 11294 16143 11328
rect 16181 11294 16201 11328
rect 16201 11294 16215 11328
rect 16253 11294 16269 11328
rect 16269 11294 16287 11328
rect 16325 11294 16337 11328
rect 16337 11294 16359 11328
rect 16397 11294 16405 11328
rect 16405 11294 16431 11328
rect 16469 11294 16473 11328
rect 16473 11294 16503 11328
rect 16541 11294 16575 11328
rect 16613 11294 16643 11328
rect 16643 11294 16647 11328
rect 16685 11294 16711 11328
rect 16711 11294 16719 11328
rect 16757 11294 16779 11328
rect 16779 11294 16791 11328
rect 16829 11294 16847 11328
rect 16847 11294 16863 11328
rect 16901 11294 16915 11328
rect 16915 11294 16935 11328
rect 16973 11294 16983 11328
rect 16983 11294 17007 11328
rect 13152 9454 13174 9460
rect 13174 9454 13186 9460
rect 13252 9454 13264 9460
rect 13264 9454 13286 9460
rect 13352 9454 13354 9460
rect 13354 9454 13386 9460
rect 13152 9426 13186 9454
rect 13252 9426 13286 9454
rect 13352 9426 13386 9454
rect 13452 9426 13486 9460
rect 13552 9426 13586 9460
rect 13652 9454 13680 9460
rect 13680 9454 13686 9460
rect 13652 9426 13686 9454
rect 13152 9326 13186 9360
rect 13252 9326 13286 9360
rect 13352 9326 13386 9360
rect 13452 9326 13486 9360
rect 13552 9326 13586 9360
rect 13652 9326 13686 9360
rect 13152 9226 13186 9260
rect 13252 9226 13286 9260
rect 13352 9226 13386 9260
rect 13452 9226 13486 9260
rect 13552 9226 13586 9260
rect 13652 9226 13686 9260
rect 13152 9128 13186 9160
rect 13252 9128 13286 9160
rect 13352 9128 13386 9160
rect 13152 9126 13174 9128
rect 13174 9126 13186 9128
rect 13252 9126 13264 9128
rect 13264 9126 13286 9128
rect 13352 9126 13354 9128
rect 13354 9126 13386 9128
rect 13452 9126 13486 9160
rect 13552 9126 13586 9160
rect 13652 9128 13686 9160
rect 13652 9126 13680 9128
rect 13680 9126 13686 9128
rect 13152 9038 13186 9060
rect 13252 9038 13286 9060
rect 13352 9038 13386 9060
rect 13152 9026 13174 9038
rect 13174 9026 13186 9038
rect 13252 9026 13264 9038
rect 13264 9026 13286 9038
rect 13352 9026 13354 9038
rect 13354 9026 13386 9038
rect 13452 9026 13486 9060
rect 13552 9026 13586 9060
rect 13652 9038 13686 9060
rect 13652 9026 13680 9038
rect 13680 9026 13686 9038
rect 13152 8948 13186 8960
rect 13252 8948 13286 8960
rect 13352 8948 13386 8960
rect 13152 8926 13174 8948
rect 13174 8926 13186 8948
rect 13252 8926 13264 8948
rect 13264 8926 13286 8948
rect 13352 8926 13354 8948
rect 13354 8926 13386 8948
rect 13452 8926 13486 8960
rect 13552 8926 13586 8960
rect 13652 8948 13686 8960
rect 13652 8926 13680 8948
rect 13680 8926 13686 8948
rect -7687 7576 -7685 7610
rect -7685 7576 -7653 7610
rect -7615 7576 -7583 7610
rect -7583 7576 -7581 7610
rect -7429 7576 -7427 7610
rect -7427 7576 -7395 7610
rect -7357 7576 -7325 7610
rect -7325 7576 -7323 7610
rect -7171 7576 -7169 7610
rect -7169 7576 -7137 7610
rect -7099 7576 -7067 7610
rect -7067 7576 -7065 7610
rect -6913 7576 -6911 7610
rect -6911 7576 -6879 7610
rect -6841 7576 -6809 7610
rect -6809 7576 -6807 7610
rect -6655 7576 -6653 7610
rect -6653 7576 -6621 7610
rect -6583 7576 -6551 7610
rect -6551 7576 -6549 7610
rect -6397 7576 -6395 7610
rect -6395 7576 -6363 7610
rect -6325 7576 -6293 7610
rect -6293 7576 -6291 7610
rect -6139 7576 -6137 7610
rect -6137 7576 -6105 7610
rect -6067 7576 -6035 7610
rect -6035 7576 -6033 7610
rect -5881 7576 -5879 7610
rect -5879 7576 -5847 7610
rect -5809 7576 -5777 7610
rect -5777 7576 -5775 7610
rect -5623 7576 -5621 7610
rect -5621 7576 -5589 7610
rect -5551 7576 -5519 7610
rect -5519 7576 -5517 7610
rect -5365 7576 -5363 7610
rect -5363 7576 -5331 7610
rect -5293 7576 -5261 7610
rect -5261 7576 -5259 7610
rect -5107 7576 -5105 7610
rect -5105 7576 -5073 7610
rect -5035 7576 -5003 7610
rect -5003 7576 -5001 7610
rect -4849 7576 -4847 7610
rect -4847 7576 -4815 7610
rect -4777 7576 -4745 7610
rect -4745 7576 -4743 7610
rect -4591 7576 -4589 7610
rect -4589 7576 -4557 7610
rect -4519 7576 -4487 7610
rect -4487 7576 -4485 7610
rect -4333 7576 -4331 7610
rect -4331 7576 -4299 7610
rect -4261 7576 -4229 7610
rect -4229 7576 -4227 7610
rect -4075 7576 -4073 7610
rect -4073 7576 -4041 7610
rect -4003 7576 -3971 7610
rect -3971 7576 -3969 7610
rect -3817 7576 -3815 7610
rect -3815 7576 -3783 7610
rect -3745 7576 -3713 7610
rect -3713 7576 -3711 7610
rect -7969 5880 -7968 5886
rect -7968 5880 -7935 5886
rect -7969 5852 -7935 5880
rect -7969 5812 -7968 5814
rect -7968 5812 -7935 5814
rect -7969 5780 -7935 5812
rect -7969 5710 -7935 5742
rect -7969 5708 -7968 5710
rect -7968 5708 -7935 5710
rect -7780 7473 -7746 7491
rect -7780 7457 -7746 7473
rect -7780 7405 -7746 7419
rect -7780 7385 -7746 7405
rect -7780 7337 -7746 7347
rect -7780 7313 -7746 7337
rect -7780 7269 -7746 7275
rect -7780 7241 -7746 7269
rect -7780 7201 -7746 7203
rect -7780 7169 -7746 7201
rect -7780 7099 -7746 7131
rect -7780 7097 -7746 7099
rect -7780 7031 -7746 7059
rect -7780 7025 -7746 7031
rect -7780 6963 -7746 6987
rect -7780 6953 -7746 6963
rect -7780 6895 -7746 6915
rect -7780 6881 -7746 6895
rect -7780 6827 -7746 6843
rect -7780 6809 -7746 6827
rect -7780 6759 -7746 6771
rect -7780 6737 -7746 6759
rect -7780 6691 -7746 6699
rect -7780 6665 -7746 6691
rect -7780 6623 -7746 6627
rect -7780 6593 -7746 6623
rect -7780 6521 -7746 6555
rect -7780 6453 -7746 6483
rect -7780 6449 -7746 6453
rect -7780 6385 -7746 6411
rect -7780 6377 -7746 6385
rect -7780 6317 -7746 6339
rect -7780 6305 -7746 6317
rect -7780 6249 -7746 6267
rect -7780 6233 -7746 6249
rect -7780 6181 -7746 6195
rect -7780 6161 -7746 6181
rect -7780 6113 -7746 6123
rect -7780 6089 -7746 6113
rect -7780 6045 -7746 6051
rect -7780 6017 -7746 6045
rect -7780 5977 -7746 5979
rect -7780 5945 -7746 5977
rect -7780 5875 -7746 5907
rect -7780 5873 -7746 5875
rect -7780 5807 -7746 5835
rect -7780 5801 -7746 5807
rect -7780 5739 -7746 5763
rect -7780 5729 -7746 5739
rect -7780 5671 -7746 5691
rect -7780 5657 -7746 5671
rect -7780 5603 -7746 5619
rect -7780 5585 -7746 5603
rect -7522 7473 -7488 7491
rect -7522 7457 -7488 7473
rect -7522 7405 -7488 7419
rect -7522 7385 -7488 7405
rect -7522 7337 -7488 7347
rect -7522 7313 -7488 7337
rect -7522 7269 -7488 7275
rect -7522 7241 -7488 7269
rect -7522 7201 -7488 7203
rect -7522 7169 -7488 7201
rect -7522 7099 -7488 7131
rect -7522 7097 -7488 7099
rect -7522 7031 -7488 7059
rect -7522 7025 -7488 7031
rect -7522 6963 -7488 6987
rect -7522 6953 -7488 6963
rect -7522 6895 -7488 6915
rect -7522 6881 -7488 6895
rect -7522 6827 -7488 6843
rect -7522 6809 -7488 6827
rect -7522 6759 -7488 6771
rect -7522 6737 -7488 6759
rect -7522 6691 -7488 6699
rect -7522 6665 -7488 6691
rect -7522 6623 -7488 6627
rect -7522 6593 -7488 6623
rect -7522 6521 -7488 6555
rect -7522 6453 -7488 6483
rect -7522 6449 -7488 6453
rect -7522 6385 -7488 6411
rect -7522 6377 -7488 6385
rect -7522 6317 -7488 6339
rect -7522 6305 -7488 6317
rect -7522 6249 -7488 6267
rect -7522 6233 -7488 6249
rect -7522 6181 -7488 6195
rect -7522 6161 -7488 6181
rect -7522 6113 -7488 6123
rect -7522 6089 -7488 6113
rect -7522 6045 -7488 6051
rect -7522 6017 -7488 6045
rect -7522 5977 -7488 5979
rect -7522 5945 -7488 5977
rect -7522 5875 -7488 5907
rect -7522 5873 -7488 5875
rect -7522 5807 -7488 5835
rect -7522 5801 -7488 5807
rect -7522 5739 -7488 5763
rect -7522 5729 -7488 5739
rect -7522 5671 -7488 5691
rect -7522 5657 -7488 5671
rect -7522 5603 -7488 5619
rect -7522 5585 -7488 5603
rect -7264 7473 -7230 7491
rect -7264 7457 -7230 7473
rect -7264 7405 -7230 7419
rect -7264 7385 -7230 7405
rect -7264 7337 -7230 7347
rect -7264 7313 -7230 7337
rect -7264 7269 -7230 7275
rect -7264 7241 -7230 7269
rect -7264 7201 -7230 7203
rect -7264 7169 -7230 7201
rect -7264 7099 -7230 7131
rect -7264 7097 -7230 7099
rect -7264 7031 -7230 7059
rect -7264 7025 -7230 7031
rect -7264 6963 -7230 6987
rect -7264 6953 -7230 6963
rect -7264 6895 -7230 6915
rect -7264 6881 -7230 6895
rect -7264 6827 -7230 6843
rect -7264 6809 -7230 6827
rect -7264 6759 -7230 6771
rect -7264 6737 -7230 6759
rect -7264 6691 -7230 6699
rect -7264 6665 -7230 6691
rect -7264 6623 -7230 6627
rect -7264 6593 -7230 6623
rect -7264 6521 -7230 6555
rect -7264 6453 -7230 6483
rect -7264 6449 -7230 6453
rect -7264 6385 -7230 6411
rect -7264 6377 -7230 6385
rect -7264 6317 -7230 6339
rect -7264 6305 -7230 6317
rect -7264 6249 -7230 6267
rect -7264 6233 -7230 6249
rect -7264 6181 -7230 6195
rect -7264 6161 -7230 6181
rect -7264 6113 -7230 6123
rect -7264 6089 -7230 6113
rect -7264 6045 -7230 6051
rect -7264 6017 -7230 6045
rect -7264 5977 -7230 5979
rect -7264 5945 -7230 5977
rect -7264 5875 -7230 5907
rect -7264 5873 -7230 5875
rect -7264 5807 -7230 5835
rect -7264 5801 -7230 5807
rect -7264 5739 -7230 5763
rect -7264 5729 -7230 5739
rect -7264 5671 -7230 5691
rect -7264 5657 -7230 5671
rect -7264 5603 -7230 5619
rect -7264 5585 -7230 5603
rect -7006 7473 -6972 7491
rect -7006 7457 -6972 7473
rect -7006 7405 -6972 7419
rect -7006 7385 -6972 7405
rect -7006 7337 -6972 7347
rect -7006 7313 -6972 7337
rect -7006 7269 -6972 7275
rect -7006 7241 -6972 7269
rect -7006 7201 -6972 7203
rect -7006 7169 -6972 7201
rect -7006 7099 -6972 7131
rect -7006 7097 -6972 7099
rect -7006 7031 -6972 7059
rect -7006 7025 -6972 7031
rect -7006 6963 -6972 6987
rect -7006 6953 -6972 6963
rect -7006 6895 -6972 6915
rect -7006 6881 -6972 6895
rect -7006 6827 -6972 6843
rect -7006 6809 -6972 6827
rect -7006 6759 -6972 6771
rect -7006 6737 -6972 6759
rect -7006 6691 -6972 6699
rect -7006 6665 -6972 6691
rect -7006 6623 -6972 6627
rect -7006 6593 -6972 6623
rect -7006 6521 -6972 6555
rect -7006 6453 -6972 6483
rect -7006 6449 -6972 6453
rect -7006 6385 -6972 6411
rect -7006 6377 -6972 6385
rect -7006 6317 -6972 6339
rect -7006 6305 -6972 6317
rect -7006 6249 -6972 6267
rect -7006 6233 -6972 6249
rect -7006 6181 -6972 6195
rect -7006 6161 -6972 6181
rect -7006 6113 -6972 6123
rect -7006 6089 -6972 6113
rect -7006 6045 -6972 6051
rect -7006 6017 -6972 6045
rect -7006 5977 -6972 5979
rect -7006 5945 -6972 5977
rect -7006 5875 -6972 5907
rect -7006 5873 -6972 5875
rect -7006 5807 -6972 5835
rect -7006 5801 -6972 5807
rect -7006 5739 -6972 5763
rect -7006 5729 -6972 5739
rect -7006 5671 -6972 5691
rect -7006 5657 -6972 5671
rect -7006 5603 -6972 5619
rect -7006 5585 -6972 5603
rect -6748 7473 -6714 7491
rect -6748 7457 -6714 7473
rect -6748 7405 -6714 7419
rect -6748 7385 -6714 7405
rect -6748 7337 -6714 7347
rect -6748 7313 -6714 7337
rect -6748 7269 -6714 7275
rect -6748 7241 -6714 7269
rect -6748 7201 -6714 7203
rect -6748 7169 -6714 7201
rect -6748 7099 -6714 7131
rect -6748 7097 -6714 7099
rect -6748 7031 -6714 7059
rect -6748 7025 -6714 7031
rect -6748 6963 -6714 6987
rect -6748 6953 -6714 6963
rect -6748 6895 -6714 6915
rect -6748 6881 -6714 6895
rect -6748 6827 -6714 6843
rect -6748 6809 -6714 6827
rect -6748 6759 -6714 6771
rect -6748 6737 -6714 6759
rect -6748 6691 -6714 6699
rect -6748 6665 -6714 6691
rect -6748 6623 -6714 6627
rect -6748 6593 -6714 6623
rect -6748 6521 -6714 6555
rect -6748 6453 -6714 6483
rect -6748 6449 -6714 6453
rect -6748 6385 -6714 6411
rect -6748 6377 -6714 6385
rect -6748 6317 -6714 6339
rect -6748 6305 -6714 6317
rect -6748 6249 -6714 6267
rect -6748 6233 -6714 6249
rect -6748 6181 -6714 6195
rect -6748 6161 -6714 6181
rect -6748 6113 -6714 6123
rect -6748 6089 -6714 6113
rect -6748 6045 -6714 6051
rect -6748 6017 -6714 6045
rect -6748 5977 -6714 5979
rect -6748 5945 -6714 5977
rect -6748 5875 -6714 5907
rect -6748 5873 -6714 5875
rect -6748 5807 -6714 5835
rect -6748 5801 -6714 5807
rect -6748 5739 -6714 5763
rect -6748 5729 -6714 5739
rect -6748 5671 -6714 5691
rect -6748 5657 -6714 5671
rect -6748 5603 -6714 5619
rect -6748 5585 -6714 5603
rect -6490 7473 -6456 7491
rect -6490 7457 -6456 7473
rect -6490 7405 -6456 7419
rect -6490 7385 -6456 7405
rect -6490 7337 -6456 7347
rect -6490 7313 -6456 7337
rect -6490 7269 -6456 7275
rect -6490 7241 -6456 7269
rect -6490 7201 -6456 7203
rect -6490 7169 -6456 7201
rect -6490 7099 -6456 7131
rect -6490 7097 -6456 7099
rect -6490 7031 -6456 7059
rect -6490 7025 -6456 7031
rect -6490 6963 -6456 6987
rect -6490 6953 -6456 6963
rect -6490 6895 -6456 6915
rect -6490 6881 -6456 6895
rect -6490 6827 -6456 6843
rect -6490 6809 -6456 6827
rect -6490 6759 -6456 6771
rect -6490 6737 -6456 6759
rect -6490 6691 -6456 6699
rect -6490 6665 -6456 6691
rect -6490 6623 -6456 6627
rect -6490 6593 -6456 6623
rect -6490 6521 -6456 6555
rect -6490 6453 -6456 6483
rect -6490 6449 -6456 6453
rect -6490 6385 -6456 6411
rect -6490 6377 -6456 6385
rect -6490 6317 -6456 6339
rect -6490 6305 -6456 6317
rect -6490 6249 -6456 6267
rect -6490 6233 -6456 6249
rect -6490 6181 -6456 6195
rect -6490 6161 -6456 6181
rect -6490 6113 -6456 6123
rect -6490 6089 -6456 6113
rect -6490 6045 -6456 6051
rect -6490 6017 -6456 6045
rect -6490 5977 -6456 5979
rect -6490 5945 -6456 5977
rect -6490 5875 -6456 5907
rect -6490 5873 -6456 5875
rect -6490 5807 -6456 5835
rect -6490 5801 -6456 5807
rect -6490 5739 -6456 5763
rect -6490 5729 -6456 5739
rect -6490 5671 -6456 5691
rect -6490 5657 -6456 5671
rect -6490 5603 -6456 5619
rect -6490 5585 -6456 5603
rect -6232 7473 -6198 7491
rect -6232 7457 -6198 7473
rect -6232 7405 -6198 7419
rect -6232 7385 -6198 7405
rect -6232 7337 -6198 7347
rect -6232 7313 -6198 7337
rect -6232 7269 -6198 7275
rect -6232 7241 -6198 7269
rect -6232 7201 -6198 7203
rect -6232 7169 -6198 7201
rect -6232 7099 -6198 7131
rect -6232 7097 -6198 7099
rect -6232 7031 -6198 7059
rect -6232 7025 -6198 7031
rect -6232 6963 -6198 6987
rect -6232 6953 -6198 6963
rect -6232 6895 -6198 6915
rect -6232 6881 -6198 6895
rect -6232 6827 -6198 6843
rect -6232 6809 -6198 6827
rect -6232 6759 -6198 6771
rect -6232 6737 -6198 6759
rect -6232 6691 -6198 6699
rect -6232 6665 -6198 6691
rect -6232 6623 -6198 6627
rect -6232 6593 -6198 6623
rect -6232 6521 -6198 6555
rect -6232 6453 -6198 6483
rect -6232 6449 -6198 6453
rect -6232 6385 -6198 6411
rect -6232 6377 -6198 6385
rect -6232 6317 -6198 6339
rect -6232 6305 -6198 6317
rect -6232 6249 -6198 6267
rect -6232 6233 -6198 6249
rect -6232 6181 -6198 6195
rect -6232 6161 -6198 6181
rect -6232 6113 -6198 6123
rect -6232 6089 -6198 6113
rect -6232 6045 -6198 6051
rect -6232 6017 -6198 6045
rect -6232 5977 -6198 5979
rect -6232 5945 -6198 5977
rect -6232 5875 -6198 5907
rect -6232 5873 -6198 5875
rect -6232 5807 -6198 5835
rect -6232 5801 -6198 5807
rect -6232 5739 -6198 5763
rect -6232 5729 -6198 5739
rect -6232 5671 -6198 5691
rect -6232 5657 -6198 5671
rect -6232 5603 -6198 5619
rect -6232 5585 -6198 5603
rect -5974 7473 -5940 7491
rect -5974 7457 -5940 7473
rect -5974 7405 -5940 7419
rect -5974 7385 -5940 7405
rect -5974 7337 -5940 7347
rect -5974 7313 -5940 7337
rect -5974 7269 -5940 7275
rect -5974 7241 -5940 7269
rect -5974 7201 -5940 7203
rect -5974 7169 -5940 7201
rect -5974 7099 -5940 7131
rect -5974 7097 -5940 7099
rect -5974 7031 -5940 7059
rect -5974 7025 -5940 7031
rect -5974 6963 -5940 6987
rect -5974 6953 -5940 6963
rect -5974 6895 -5940 6915
rect -5974 6881 -5940 6895
rect -5974 6827 -5940 6843
rect -5974 6809 -5940 6827
rect -5974 6759 -5940 6771
rect -5974 6737 -5940 6759
rect -5974 6691 -5940 6699
rect -5974 6665 -5940 6691
rect -5974 6623 -5940 6627
rect -5974 6593 -5940 6623
rect -5974 6521 -5940 6555
rect -5974 6453 -5940 6483
rect -5974 6449 -5940 6453
rect -5974 6385 -5940 6411
rect -5974 6377 -5940 6385
rect -5974 6317 -5940 6339
rect -5974 6305 -5940 6317
rect -5974 6249 -5940 6267
rect -5974 6233 -5940 6249
rect -5974 6181 -5940 6195
rect -5974 6161 -5940 6181
rect -5974 6113 -5940 6123
rect -5974 6089 -5940 6113
rect -5974 6045 -5940 6051
rect -5974 6017 -5940 6045
rect -5974 5977 -5940 5979
rect -5974 5945 -5940 5977
rect -5974 5875 -5940 5907
rect -5974 5873 -5940 5875
rect -5974 5807 -5940 5835
rect -5974 5801 -5940 5807
rect -5974 5739 -5940 5763
rect -5974 5729 -5940 5739
rect -5974 5671 -5940 5691
rect -5974 5657 -5940 5671
rect -5974 5603 -5940 5619
rect -5974 5585 -5940 5603
rect -5716 7473 -5682 7491
rect -5716 7457 -5682 7473
rect -5716 7405 -5682 7419
rect -5716 7385 -5682 7405
rect -5716 7337 -5682 7347
rect -5716 7313 -5682 7337
rect -5716 7269 -5682 7275
rect -5716 7241 -5682 7269
rect -5716 7201 -5682 7203
rect -5716 7169 -5682 7201
rect -5716 7099 -5682 7131
rect -5716 7097 -5682 7099
rect -5716 7031 -5682 7059
rect -5716 7025 -5682 7031
rect -5716 6963 -5682 6987
rect -5716 6953 -5682 6963
rect -5716 6895 -5682 6915
rect -5716 6881 -5682 6895
rect -5716 6827 -5682 6843
rect -5716 6809 -5682 6827
rect -5716 6759 -5682 6771
rect -5716 6737 -5682 6759
rect -5716 6691 -5682 6699
rect -5716 6665 -5682 6691
rect -5716 6623 -5682 6627
rect -5716 6593 -5682 6623
rect -5716 6521 -5682 6555
rect -5716 6453 -5682 6483
rect -5716 6449 -5682 6453
rect -5716 6385 -5682 6411
rect -5716 6377 -5682 6385
rect -5716 6317 -5682 6339
rect -5716 6305 -5682 6317
rect -5716 6249 -5682 6267
rect -5716 6233 -5682 6249
rect -5716 6181 -5682 6195
rect -5716 6161 -5682 6181
rect -5716 6113 -5682 6123
rect -5716 6089 -5682 6113
rect -5716 6045 -5682 6051
rect -5716 6017 -5682 6045
rect -5716 5977 -5682 5979
rect -5716 5945 -5682 5977
rect -5716 5875 -5682 5907
rect -5716 5873 -5682 5875
rect -5716 5807 -5682 5835
rect -5716 5801 -5682 5807
rect -5716 5739 -5682 5763
rect -5716 5729 -5682 5739
rect -5716 5671 -5682 5691
rect -5716 5657 -5682 5671
rect -5716 5603 -5682 5619
rect -5716 5585 -5682 5603
rect -5458 7473 -5424 7491
rect -5458 7457 -5424 7473
rect -5458 7405 -5424 7419
rect -5458 7385 -5424 7405
rect -5458 7337 -5424 7347
rect -5458 7313 -5424 7337
rect -5458 7269 -5424 7275
rect -5458 7241 -5424 7269
rect -5458 7201 -5424 7203
rect -5458 7169 -5424 7201
rect -5458 7099 -5424 7131
rect -5458 7097 -5424 7099
rect -5458 7031 -5424 7059
rect -5458 7025 -5424 7031
rect -5458 6963 -5424 6987
rect -5458 6953 -5424 6963
rect -5458 6895 -5424 6915
rect -5458 6881 -5424 6895
rect -5458 6827 -5424 6843
rect -5458 6809 -5424 6827
rect -5458 6759 -5424 6771
rect -5458 6737 -5424 6759
rect -5458 6691 -5424 6699
rect -5458 6665 -5424 6691
rect -5458 6623 -5424 6627
rect -5458 6593 -5424 6623
rect -5458 6521 -5424 6555
rect -5458 6453 -5424 6483
rect -5458 6449 -5424 6453
rect -5458 6385 -5424 6411
rect -5458 6377 -5424 6385
rect -5458 6317 -5424 6339
rect -5458 6305 -5424 6317
rect -5458 6249 -5424 6267
rect -5458 6233 -5424 6249
rect -5458 6181 -5424 6195
rect -5458 6161 -5424 6181
rect -5458 6113 -5424 6123
rect -5458 6089 -5424 6113
rect -5458 6045 -5424 6051
rect -5458 6017 -5424 6045
rect -5458 5977 -5424 5979
rect -5458 5945 -5424 5977
rect -5458 5875 -5424 5907
rect -5458 5873 -5424 5875
rect -5458 5807 -5424 5835
rect -5458 5801 -5424 5807
rect -5458 5739 -5424 5763
rect -5458 5729 -5424 5739
rect -5458 5671 -5424 5691
rect -5458 5657 -5424 5671
rect -5458 5603 -5424 5619
rect -5458 5585 -5424 5603
rect -5200 7473 -5166 7491
rect -5200 7457 -5166 7473
rect -5200 7405 -5166 7419
rect -5200 7385 -5166 7405
rect -5200 7337 -5166 7347
rect -5200 7313 -5166 7337
rect -5200 7269 -5166 7275
rect -5200 7241 -5166 7269
rect -5200 7201 -5166 7203
rect -5200 7169 -5166 7201
rect -5200 7099 -5166 7131
rect -5200 7097 -5166 7099
rect -5200 7031 -5166 7059
rect -5200 7025 -5166 7031
rect -5200 6963 -5166 6987
rect -5200 6953 -5166 6963
rect -5200 6895 -5166 6915
rect -5200 6881 -5166 6895
rect -5200 6827 -5166 6843
rect -5200 6809 -5166 6827
rect -5200 6759 -5166 6771
rect -5200 6737 -5166 6759
rect -5200 6691 -5166 6699
rect -5200 6665 -5166 6691
rect -5200 6623 -5166 6627
rect -5200 6593 -5166 6623
rect -5200 6521 -5166 6555
rect -5200 6453 -5166 6483
rect -5200 6449 -5166 6453
rect -5200 6385 -5166 6411
rect -5200 6377 -5166 6385
rect -5200 6317 -5166 6339
rect -5200 6305 -5166 6317
rect -5200 6249 -5166 6267
rect -5200 6233 -5166 6249
rect -5200 6181 -5166 6195
rect -5200 6161 -5166 6181
rect -5200 6113 -5166 6123
rect -5200 6089 -5166 6113
rect -5200 6045 -5166 6051
rect -5200 6017 -5166 6045
rect -5200 5977 -5166 5979
rect -5200 5945 -5166 5977
rect -5200 5875 -5166 5907
rect -5200 5873 -5166 5875
rect -5200 5807 -5166 5835
rect -5200 5801 -5166 5807
rect -5200 5739 -5166 5763
rect -5200 5729 -5166 5739
rect -5200 5671 -5166 5691
rect -5200 5657 -5166 5671
rect -5200 5603 -5166 5619
rect -5200 5585 -5166 5603
rect -4942 7473 -4908 7491
rect -4942 7457 -4908 7473
rect -4942 7405 -4908 7419
rect -4942 7385 -4908 7405
rect -4942 7337 -4908 7347
rect -4942 7313 -4908 7337
rect -4942 7269 -4908 7275
rect -4942 7241 -4908 7269
rect -4942 7201 -4908 7203
rect -4942 7169 -4908 7201
rect -4942 7099 -4908 7131
rect -4942 7097 -4908 7099
rect -4942 7031 -4908 7059
rect -4942 7025 -4908 7031
rect -4942 6963 -4908 6987
rect -4942 6953 -4908 6963
rect -4942 6895 -4908 6915
rect -4942 6881 -4908 6895
rect -4942 6827 -4908 6843
rect -4942 6809 -4908 6827
rect -4942 6759 -4908 6771
rect -4942 6737 -4908 6759
rect -4942 6691 -4908 6699
rect -4942 6665 -4908 6691
rect -4942 6623 -4908 6627
rect -4942 6593 -4908 6623
rect -4942 6521 -4908 6555
rect -4942 6453 -4908 6483
rect -4942 6449 -4908 6453
rect -4942 6385 -4908 6411
rect -4942 6377 -4908 6385
rect -4942 6317 -4908 6339
rect -4942 6305 -4908 6317
rect -4942 6249 -4908 6267
rect -4942 6233 -4908 6249
rect -4942 6181 -4908 6195
rect -4942 6161 -4908 6181
rect -4942 6113 -4908 6123
rect -4942 6089 -4908 6113
rect -4942 6045 -4908 6051
rect -4942 6017 -4908 6045
rect -4942 5977 -4908 5979
rect -4942 5945 -4908 5977
rect -4942 5875 -4908 5907
rect -4942 5873 -4908 5875
rect -4942 5807 -4908 5835
rect -4942 5801 -4908 5807
rect -4942 5739 -4908 5763
rect -4942 5729 -4908 5739
rect -4942 5671 -4908 5691
rect -4942 5657 -4908 5671
rect -4942 5603 -4908 5619
rect -4942 5585 -4908 5603
rect -4684 7473 -4650 7491
rect -4684 7457 -4650 7473
rect -4684 7405 -4650 7419
rect -4684 7385 -4650 7405
rect -4684 7337 -4650 7347
rect -4684 7313 -4650 7337
rect -4684 7269 -4650 7275
rect -4684 7241 -4650 7269
rect -4684 7201 -4650 7203
rect -4684 7169 -4650 7201
rect -4684 7099 -4650 7131
rect -4684 7097 -4650 7099
rect -4684 7031 -4650 7059
rect -4684 7025 -4650 7031
rect -4684 6963 -4650 6987
rect -4684 6953 -4650 6963
rect -4684 6895 -4650 6915
rect -4684 6881 -4650 6895
rect -4684 6827 -4650 6843
rect -4684 6809 -4650 6827
rect -4684 6759 -4650 6771
rect -4684 6737 -4650 6759
rect -4684 6691 -4650 6699
rect -4684 6665 -4650 6691
rect -4684 6623 -4650 6627
rect -4684 6593 -4650 6623
rect -4684 6521 -4650 6555
rect -4684 6453 -4650 6483
rect -4684 6449 -4650 6453
rect -4684 6385 -4650 6411
rect -4684 6377 -4650 6385
rect -4684 6317 -4650 6339
rect -4684 6305 -4650 6317
rect -4684 6249 -4650 6267
rect -4684 6233 -4650 6249
rect -4684 6181 -4650 6195
rect -4684 6161 -4650 6181
rect -4684 6113 -4650 6123
rect -4684 6089 -4650 6113
rect -4684 6045 -4650 6051
rect -4684 6017 -4650 6045
rect -4684 5977 -4650 5979
rect -4684 5945 -4650 5977
rect -4684 5875 -4650 5907
rect -4684 5873 -4650 5875
rect -4684 5807 -4650 5835
rect -4684 5801 -4650 5807
rect -4684 5739 -4650 5763
rect -4684 5729 -4650 5739
rect -4684 5671 -4650 5691
rect -4684 5657 -4650 5671
rect -4684 5603 -4650 5619
rect -4684 5585 -4650 5603
rect -4426 7473 -4392 7491
rect -4426 7457 -4392 7473
rect -4426 7405 -4392 7419
rect -4426 7385 -4392 7405
rect -4426 7337 -4392 7347
rect -4426 7313 -4392 7337
rect -4426 7269 -4392 7275
rect -4426 7241 -4392 7269
rect -4426 7201 -4392 7203
rect -4426 7169 -4392 7201
rect -4426 7099 -4392 7131
rect -4426 7097 -4392 7099
rect -4426 7031 -4392 7059
rect -4426 7025 -4392 7031
rect -4426 6963 -4392 6987
rect -4426 6953 -4392 6963
rect -4426 6895 -4392 6915
rect -4426 6881 -4392 6895
rect -4426 6827 -4392 6843
rect -4426 6809 -4392 6827
rect -4426 6759 -4392 6771
rect -4426 6737 -4392 6759
rect -4426 6691 -4392 6699
rect -4426 6665 -4392 6691
rect -4426 6623 -4392 6627
rect -4426 6593 -4392 6623
rect -4426 6521 -4392 6555
rect -4426 6453 -4392 6483
rect -4426 6449 -4392 6453
rect -4426 6385 -4392 6411
rect -4426 6377 -4392 6385
rect -4426 6317 -4392 6339
rect -4426 6305 -4392 6317
rect -4426 6249 -4392 6267
rect -4426 6233 -4392 6249
rect -4426 6181 -4392 6195
rect -4426 6161 -4392 6181
rect -4426 6113 -4392 6123
rect -4426 6089 -4392 6113
rect -4426 6045 -4392 6051
rect -4426 6017 -4392 6045
rect -4426 5977 -4392 5979
rect -4426 5945 -4392 5977
rect -4426 5875 -4392 5907
rect -4426 5873 -4392 5875
rect -4426 5807 -4392 5835
rect -4426 5801 -4392 5807
rect -4426 5739 -4392 5763
rect -4426 5729 -4392 5739
rect -4426 5671 -4392 5691
rect -4426 5657 -4392 5671
rect -4426 5603 -4392 5619
rect -4426 5585 -4392 5603
rect -4168 7473 -4134 7491
rect -4168 7457 -4134 7473
rect -4168 7405 -4134 7419
rect -4168 7385 -4134 7405
rect -4168 7337 -4134 7347
rect -4168 7313 -4134 7337
rect -4168 7269 -4134 7275
rect -4168 7241 -4134 7269
rect -4168 7201 -4134 7203
rect -4168 7169 -4134 7201
rect -4168 7099 -4134 7131
rect -4168 7097 -4134 7099
rect -4168 7031 -4134 7059
rect -4168 7025 -4134 7031
rect -4168 6963 -4134 6987
rect -4168 6953 -4134 6963
rect -4168 6895 -4134 6915
rect -4168 6881 -4134 6895
rect -4168 6827 -4134 6843
rect -4168 6809 -4134 6827
rect -4168 6759 -4134 6771
rect -4168 6737 -4134 6759
rect -4168 6691 -4134 6699
rect -4168 6665 -4134 6691
rect -4168 6623 -4134 6627
rect -4168 6593 -4134 6623
rect -4168 6521 -4134 6555
rect -4168 6453 -4134 6483
rect -4168 6449 -4134 6453
rect -4168 6385 -4134 6411
rect -4168 6377 -4134 6385
rect -4168 6317 -4134 6339
rect -4168 6305 -4134 6317
rect -4168 6249 -4134 6267
rect -4168 6233 -4134 6249
rect -4168 6181 -4134 6195
rect -4168 6161 -4134 6181
rect -4168 6113 -4134 6123
rect -4168 6089 -4134 6113
rect -4168 6045 -4134 6051
rect -4168 6017 -4134 6045
rect -4168 5977 -4134 5979
rect -4168 5945 -4134 5977
rect -4168 5875 -4134 5907
rect -4168 5873 -4134 5875
rect -4168 5807 -4134 5835
rect -4168 5801 -4134 5807
rect -4168 5739 -4134 5763
rect -4168 5729 -4134 5739
rect -4168 5671 -4134 5691
rect -4168 5657 -4134 5671
rect -4168 5603 -4134 5619
rect -4168 5585 -4134 5603
rect -3910 7473 -3876 7491
rect -3910 7457 -3876 7473
rect -3910 7405 -3876 7419
rect -3910 7385 -3876 7405
rect -3910 7337 -3876 7347
rect -3910 7313 -3876 7337
rect -3910 7269 -3876 7275
rect -3910 7241 -3876 7269
rect -3910 7201 -3876 7203
rect -3910 7169 -3876 7201
rect -3910 7099 -3876 7131
rect -3910 7097 -3876 7099
rect -3910 7031 -3876 7059
rect -3910 7025 -3876 7031
rect -3910 6963 -3876 6987
rect -3910 6953 -3876 6963
rect -3910 6895 -3876 6915
rect -3910 6881 -3876 6895
rect -3910 6827 -3876 6843
rect -3910 6809 -3876 6827
rect -3910 6759 -3876 6771
rect -3910 6737 -3876 6759
rect -3910 6691 -3876 6699
rect -3910 6665 -3876 6691
rect -3910 6623 -3876 6627
rect -3910 6593 -3876 6623
rect -3910 6521 -3876 6555
rect -3910 6453 -3876 6483
rect -3910 6449 -3876 6453
rect -3910 6385 -3876 6411
rect -3910 6377 -3876 6385
rect -3910 6317 -3876 6339
rect -3910 6305 -3876 6317
rect -3910 6249 -3876 6267
rect -3910 6233 -3876 6249
rect -3910 6181 -3876 6195
rect -3910 6161 -3876 6181
rect -3910 6113 -3876 6123
rect -3910 6089 -3876 6113
rect -3910 6045 -3876 6051
rect -3910 6017 -3876 6045
rect -3910 5977 -3876 5979
rect -3910 5945 -3876 5977
rect -3910 5875 -3876 5907
rect -3910 5873 -3876 5875
rect -3910 5807 -3876 5835
rect -3910 5801 -3876 5807
rect -3910 5739 -3876 5763
rect -3910 5729 -3876 5739
rect -3910 5671 -3876 5691
rect -3910 5657 -3876 5671
rect -3910 5603 -3876 5619
rect -3910 5585 -3876 5603
rect -3652 7473 -3618 7491
rect -3652 7457 -3618 7473
rect -3652 7405 -3618 7419
rect -3652 7385 -3618 7405
rect -3652 7337 -3618 7347
rect -3652 7313 -3618 7337
rect -3652 7269 -3618 7275
rect -3652 7241 -3618 7269
rect -3652 7201 -3618 7203
rect -3652 7169 -3618 7201
rect -3652 7099 -3618 7131
rect -3652 7097 -3618 7099
rect -3652 7031 -3618 7059
rect -3652 7025 -3618 7031
rect -3652 6963 -3618 6987
rect -3652 6953 -3618 6963
rect -3652 6895 -3618 6915
rect -3652 6881 -3618 6895
rect -3652 6827 -3618 6843
rect -3652 6809 -3618 6827
rect -3652 6759 -3618 6771
rect -3652 6737 -3618 6759
rect -3652 6691 -3618 6699
rect -3652 6665 -3618 6691
rect -3652 6623 -3618 6627
rect -3652 6593 -3618 6623
rect -3652 6521 -3618 6555
rect -3652 6453 -3618 6483
rect -3652 6449 -3618 6453
rect -3652 6385 -3618 6411
rect -3652 6377 -3618 6385
rect -3652 6317 -3618 6339
rect -3652 6305 -3618 6317
rect -3652 6249 -3618 6267
rect -3652 6233 -3618 6249
rect -3652 6181 -3618 6195
rect -3652 6161 -3618 6181
rect -3652 6113 -3618 6123
rect -3652 6089 -3618 6113
rect -3652 6045 -3618 6051
rect -3652 6017 -3618 6045
rect -3652 5977 -3618 5979
rect -3652 5945 -3618 5977
rect -3652 5875 -3618 5907
rect -3652 5873 -3618 5875
rect -3652 5807 -3618 5835
rect -3652 5801 -3618 5807
rect -3652 5739 -3618 5763
rect -3652 5729 -3618 5739
rect -3652 5671 -3618 5691
rect -3652 5657 -3618 5671
rect -3652 5603 -3618 5619
rect -3652 5585 -3618 5603
rect -3456 5858 -3422 5885
rect -3456 5851 -3422 5858
rect -3456 5790 -3422 5813
rect -3456 5779 -3422 5790
rect -3456 5722 -3422 5741
rect -3456 5707 -3422 5722
rect -7687 5466 -7685 5500
rect -7685 5466 -7653 5500
rect -7615 5466 -7583 5500
rect -7583 5466 -7581 5500
rect -7429 5466 -7427 5500
rect -7427 5466 -7395 5500
rect -7357 5466 -7325 5500
rect -7325 5466 -7323 5500
rect -7171 5466 -7169 5500
rect -7169 5466 -7137 5500
rect -7099 5466 -7067 5500
rect -7067 5466 -7065 5500
rect -6913 5466 -6911 5500
rect -6911 5466 -6879 5500
rect -6841 5466 -6809 5500
rect -6809 5466 -6807 5500
rect -6655 5466 -6653 5500
rect -6653 5466 -6621 5500
rect -6583 5466 -6551 5500
rect -6551 5466 -6549 5500
rect -6397 5466 -6395 5500
rect -6395 5466 -6363 5500
rect -6325 5466 -6293 5500
rect -6293 5466 -6291 5500
rect -6139 5466 -6137 5500
rect -6137 5466 -6105 5500
rect -6067 5466 -6035 5500
rect -6035 5466 -6033 5500
rect -5881 5466 -5879 5500
rect -5879 5466 -5847 5500
rect -5809 5466 -5777 5500
rect -5777 5466 -5775 5500
rect -5623 5466 -5621 5500
rect -5621 5466 -5589 5500
rect -5551 5466 -5519 5500
rect -5519 5466 -5517 5500
rect -5365 5466 -5363 5500
rect -5363 5466 -5331 5500
rect -5293 5466 -5261 5500
rect -5261 5466 -5259 5500
rect -5107 5466 -5105 5500
rect -5105 5466 -5073 5500
rect -5035 5466 -5003 5500
rect -5003 5466 -5001 5500
rect -4849 5466 -4847 5500
rect -4847 5466 -4815 5500
rect -4777 5466 -4745 5500
rect -4745 5466 -4743 5500
rect -4591 5466 -4589 5500
rect -4589 5466 -4557 5500
rect -4519 5466 -4487 5500
rect -4487 5466 -4485 5500
rect -4333 5466 -4331 5500
rect -4331 5466 -4299 5500
rect -4261 5466 -4229 5500
rect -4229 5466 -4227 5500
rect -4075 5466 -4073 5500
rect -4073 5466 -4041 5500
rect -4003 5466 -3971 5500
rect -3971 5466 -3969 5500
rect -3817 5466 -3815 5500
rect -3815 5466 -3783 5500
rect -3745 5466 -3713 5500
rect -3713 5466 -3711 5500
rect 13142 8044 13164 8050
rect 13164 8044 13176 8050
rect 13242 8044 13254 8050
rect 13254 8044 13276 8050
rect 13342 8044 13344 8050
rect 13344 8044 13376 8050
rect 13142 8016 13176 8044
rect 13242 8016 13276 8044
rect 13342 8016 13376 8044
rect 13442 8016 13476 8050
rect 13542 8016 13576 8050
rect 13642 8044 13670 8050
rect 13670 8044 13676 8050
rect 13642 8016 13676 8044
rect 13142 7916 13176 7950
rect 13242 7916 13276 7950
rect 13342 7916 13376 7950
rect 13442 7916 13476 7950
rect 13542 7916 13576 7950
rect 13642 7916 13676 7950
rect 13142 7816 13176 7850
rect 13242 7816 13276 7850
rect 13342 7816 13376 7850
rect 13442 7816 13476 7850
rect 13542 7816 13576 7850
rect 13642 7816 13676 7850
rect 13142 7718 13176 7750
rect 13242 7718 13276 7750
rect 13342 7718 13376 7750
rect 13142 7716 13164 7718
rect 13164 7716 13176 7718
rect 13242 7716 13254 7718
rect 13254 7716 13276 7718
rect 13342 7716 13344 7718
rect 13344 7716 13376 7718
rect 13442 7716 13476 7750
rect 13542 7716 13576 7750
rect 13642 7718 13676 7750
rect 13642 7716 13670 7718
rect 13670 7716 13676 7718
rect 13142 7628 13176 7650
rect 13242 7628 13276 7650
rect 13342 7628 13376 7650
rect 13142 7616 13164 7628
rect 13164 7616 13176 7628
rect 13242 7616 13254 7628
rect 13254 7616 13276 7628
rect 13342 7616 13344 7628
rect 13344 7616 13376 7628
rect 13442 7616 13476 7650
rect 13542 7616 13576 7650
rect 13642 7628 13676 7650
rect 13642 7616 13670 7628
rect 13670 7616 13676 7628
rect 13142 7538 13176 7550
rect 13242 7538 13276 7550
rect 13342 7538 13376 7550
rect 13142 7516 13164 7538
rect 13164 7516 13176 7538
rect 13242 7516 13254 7538
rect 13254 7516 13276 7538
rect 13342 7516 13344 7538
rect 13344 7516 13376 7538
rect 13442 7516 13476 7550
rect 13542 7516 13576 7550
rect 13642 7538 13676 7550
rect 13642 7516 13670 7538
rect 13670 7516 13676 7538
rect 14954 11192 14988 11204
rect 14954 11170 14988 11192
rect 14954 11124 14988 11132
rect 14954 11098 14988 11124
rect 14954 11056 14988 11060
rect 14954 11026 14988 11056
rect 14954 10954 14988 10988
rect 14954 10886 14988 10916
rect 14954 10882 14988 10886
rect 14954 10818 14988 10844
rect 14954 10810 14988 10818
rect 14954 10750 14988 10772
rect 14954 10738 14988 10750
rect 14954 10682 14988 10700
rect 14954 10666 14988 10682
rect 14954 10614 14988 10628
rect 14954 10594 14988 10614
rect 14954 10546 14988 10556
rect 14954 10522 14988 10546
rect 14954 10478 14988 10484
rect 14954 10450 14988 10478
rect 14954 10410 14988 10412
rect 14954 10378 14988 10410
rect 14954 10308 14988 10340
rect 14954 10306 14988 10308
rect 14954 10240 14988 10268
rect 14954 10234 14988 10240
rect 14954 10172 14988 10196
rect 14954 10162 14988 10172
rect 14954 10104 14988 10124
rect 14954 10090 14988 10104
rect 14954 10036 14988 10052
rect 14954 10018 14988 10036
rect 14954 9968 14988 9980
rect 14954 9946 14988 9968
rect 14954 9900 14988 9908
rect 14954 9874 14988 9900
rect 14954 9832 14988 9836
rect 14954 9802 14988 9832
rect 14954 9730 14988 9764
rect 14954 9662 14988 9692
rect 14954 9658 14988 9662
rect 14954 9594 14988 9620
rect 14954 9586 14988 9594
rect 14954 9526 14988 9548
rect 14954 9514 14988 9526
rect 14954 9458 14988 9476
rect 14954 9442 14988 9458
rect 14954 9390 14988 9404
rect 14954 9370 14988 9390
rect 14954 9322 14988 9332
rect 14954 9298 14988 9322
rect 14954 9254 14988 9260
rect 14954 9226 14988 9254
rect 14954 9186 14988 9188
rect 14954 9154 14988 9186
rect 14954 9084 14988 9116
rect 14954 9082 14988 9084
rect 14954 9016 14988 9044
rect 14954 9010 14988 9016
rect 14954 8948 14988 8972
rect 14954 8938 14988 8948
rect 14954 8880 14988 8900
rect 14954 8866 14988 8880
rect 14954 8812 14988 8828
rect 14954 8794 14988 8812
rect 14954 8744 14988 8756
rect 14954 8722 14988 8744
rect 14954 8676 14988 8684
rect 14954 8650 14988 8676
rect 14954 8608 14988 8612
rect 14954 8578 14988 8608
rect 14954 8506 14988 8540
rect 14954 8438 14988 8468
rect 14954 8434 14988 8438
rect 14954 8370 14988 8396
rect 14954 8362 14988 8370
rect 14954 8302 14988 8324
rect 14954 8290 14988 8302
rect 16012 11192 16046 11204
rect 16012 11170 16046 11192
rect 16012 11124 16046 11132
rect 16012 11098 16046 11124
rect 16012 11056 16046 11060
rect 16012 11026 16046 11056
rect 16012 10954 16046 10988
rect 16012 10886 16046 10916
rect 16012 10882 16046 10886
rect 16012 10818 16046 10844
rect 16012 10810 16046 10818
rect 16012 10750 16046 10772
rect 16012 10738 16046 10750
rect 16012 10682 16046 10700
rect 16012 10666 16046 10682
rect 16012 10614 16046 10628
rect 16012 10594 16046 10614
rect 16012 10546 16046 10556
rect 16012 10522 16046 10546
rect 16012 10478 16046 10484
rect 16012 10450 16046 10478
rect 16012 10410 16046 10412
rect 16012 10378 16046 10410
rect 16012 10308 16046 10340
rect 16012 10306 16046 10308
rect 16012 10240 16046 10268
rect 16012 10234 16046 10240
rect 16012 10172 16046 10196
rect 16012 10162 16046 10172
rect 16012 10104 16046 10124
rect 16012 10090 16046 10104
rect 16012 10036 16046 10052
rect 16012 10018 16046 10036
rect 16012 9968 16046 9980
rect 16012 9946 16046 9968
rect 16012 9900 16046 9908
rect 16012 9874 16046 9900
rect 16012 9832 16046 9836
rect 16012 9802 16046 9832
rect 16012 9730 16046 9764
rect 16012 9662 16046 9692
rect 16012 9658 16046 9662
rect 16012 9594 16046 9620
rect 16012 9586 16046 9594
rect 16012 9526 16046 9548
rect 16012 9514 16046 9526
rect 16012 9458 16046 9476
rect 16012 9442 16046 9458
rect 16012 9390 16046 9404
rect 16012 9370 16046 9390
rect 16012 9322 16046 9332
rect 16012 9298 16046 9322
rect 16012 9254 16046 9260
rect 16012 9226 16046 9254
rect 16012 9186 16046 9188
rect 16012 9154 16046 9186
rect 16012 9084 16046 9116
rect 16012 9082 16046 9084
rect 16012 9016 16046 9044
rect 16012 9010 16046 9016
rect 16012 8948 16046 8972
rect 16012 8938 16046 8948
rect 16012 8880 16046 8900
rect 16012 8866 16046 8880
rect 16012 8812 16046 8828
rect 16012 8794 16046 8812
rect 16012 8744 16046 8756
rect 16012 8722 16046 8744
rect 16012 8676 16046 8684
rect 16012 8650 16046 8676
rect 16012 8608 16046 8612
rect 16012 8578 16046 8608
rect 16012 8506 16046 8540
rect 16012 8438 16046 8468
rect 16012 8434 16046 8438
rect 16012 8370 16046 8396
rect 16012 8362 16046 8370
rect 16012 8302 16046 8324
rect 16012 8290 16046 8302
rect 17070 11192 17104 11204
rect 17070 11170 17104 11192
rect 17070 11124 17104 11132
rect 17070 11098 17104 11124
rect 17070 11056 17104 11060
rect 17070 11026 17104 11056
rect 17070 10954 17104 10988
rect 17070 10886 17104 10916
rect 17070 10882 17104 10886
rect 17070 10818 17104 10844
rect 17070 10810 17104 10818
rect 17070 10750 17104 10772
rect 17070 10738 17104 10750
rect 17070 10682 17104 10700
rect 17070 10666 17104 10682
rect 17070 10614 17104 10628
rect 17070 10594 17104 10614
rect 17070 10546 17104 10556
rect 17070 10522 17104 10546
rect 17070 10478 17104 10484
rect 17070 10450 17104 10478
rect 17070 10410 17104 10412
rect 17070 10378 17104 10410
rect 17070 10308 17104 10340
rect 17070 10306 17104 10308
rect 17070 10240 17104 10268
rect 17070 10234 17104 10240
rect 17070 10172 17104 10196
rect 17070 10162 17104 10172
rect 17070 10104 17104 10124
rect 17070 10090 17104 10104
rect 17070 10036 17104 10052
rect 17070 10018 17104 10036
rect 17070 9968 17104 9980
rect 17070 9946 17104 9968
rect 17070 9900 17104 9908
rect 17070 9874 17104 9900
rect 17070 9832 17104 9836
rect 17070 9802 17104 9832
rect 17070 9730 17104 9764
rect 17070 9662 17104 9692
rect 17070 9658 17104 9662
rect 17070 9594 17104 9620
rect 17070 9586 17104 9594
rect 17070 9526 17104 9548
rect 17070 9514 17104 9526
rect 17070 9458 17104 9476
rect 17070 9442 17104 9458
rect 17070 9390 17104 9404
rect 17070 9370 17104 9390
rect 17070 9322 17104 9332
rect 17070 9298 17104 9322
rect 17070 9254 17104 9260
rect 17070 9226 17104 9254
rect 17070 9186 17104 9188
rect 17070 9154 17104 9186
rect 17070 9084 17104 9116
rect 17070 9082 17104 9084
rect 17070 9016 17104 9044
rect 17070 9010 17104 9016
rect 17070 8948 17104 8972
rect 17070 8938 17104 8948
rect 17070 8880 17104 8900
rect 17070 8866 17104 8880
rect 17070 8812 17104 8828
rect 17070 8794 17104 8812
rect 17070 8744 17104 8756
rect 17070 8722 17104 8744
rect 17070 8676 17104 8684
rect 17070 8650 17104 8676
rect 17070 8608 17104 8612
rect 17070 8578 17104 8608
rect 17070 8506 17104 8540
rect 17070 8438 17104 8468
rect 17070 8434 17104 8438
rect 17070 8370 17104 8396
rect 17070 8362 17104 8370
rect 17070 8302 17104 8324
rect 17070 8290 17104 8302
rect 15051 8166 15075 8200
rect 15075 8166 15085 8200
rect 15123 8166 15143 8200
rect 15143 8166 15157 8200
rect 15195 8166 15211 8200
rect 15211 8166 15229 8200
rect 15267 8166 15279 8200
rect 15279 8166 15301 8200
rect 15339 8166 15347 8200
rect 15347 8166 15373 8200
rect 15411 8166 15415 8200
rect 15415 8166 15445 8200
rect 15483 8166 15517 8200
rect 15555 8166 15585 8200
rect 15585 8166 15589 8200
rect 15627 8166 15653 8200
rect 15653 8166 15661 8200
rect 15699 8166 15721 8200
rect 15721 8166 15733 8200
rect 15771 8166 15789 8200
rect 15789 8166 15805 8200
rect 15843 8166 15857 8200
rect 15857 8166 15877 8200
rect 15915 8166 15925 8200
rect 15925 8166 15949 8200
rect 16109 8166 16133 8200
rect 16133 8166 16143 8200
rect 16181 8166 16201 8200
rect 16201 8166 16215 8200
rect 16253 8166 16269 8200
rect 16269 8166 16287 8200
rect 16325 8166 16337 8200
rect 16337 8166 16359 8200
rect 16397 8166 16405 8200
rect 16405 8166 16431 8200
rect 16469 8166 16473 8200
rect 16473 8166 16503 8200
rect 16541 8166 16575 8200
rect 16613 8166 16643 8200
rect 16643 8166 16647 8200
rect 16685 8166 16711 8200
rect 16711 8166 16719 8200
rect 16757 8166 16779 8200
rect 16779 8166 16791 8200
rect 16829 8166 16847 8200
rect 16847 8166 16863 8200
rect 16901 8166 16915 8200
rect 16915 8166 16935 8200
rect 16973 8166 16983 8200
rect 16983 8166 17007 8200
rect 17575 11268 17599 11302
rect 17599 11268 17609 11302
rect 17647 11268 17667 11302
rect 17667 11268 17681 11302
rect 17719 11268 17735 11302
rect 17735 11268 17753 11302
rect 17791 11268 17803 11302
rect 17803 11268 17825 11302
rect 17863 11268 17871 11302
rect 17871 11268 17897 11302
rect 17935 11268 17939 11302
rect 17939 11268 17969 11302
rect 18007 11268 18041 11302
rect 18079 11268 18109 11302
rect 18109 11268 18113 11302
rect 18151 11268 18177 11302
rect 18177 11268 18185 11302
rect 18223 11268 18245 11302
rect 18245 11268 18257 11302
rect 18295 11268 18313 11302
rect 18313 11268 18329 11302
rect 18367 11268 18381 11302
rect 18381 11268 18401 11302
rect 18439 11268 18449 11302
rect 18449 11268 18473 11302
rect 18633 11268 18657 11302
rect 18657 11268 18667 11302
rect 18705 11268 18725 11302
rect 18725 11268 18739 11302
rect 18777 11268 18793 11302
rect 18793 11268 18811 11302
rect 18849 11268 18861 11302
rect 18861 11268 18883 11302
rect 18921 11268 18929 11302
rect 18929 11268 18955 11302
rect 18993 11268 18997 11302
rect 18997 11268 19027 11302
rect 19065 11268 19099 11302
rect 19137 11268 19167 11302
rect 19167 11268 19171 11302
rect 19209 11268 19235 11302
rect 19235 11268 19243 11302
rect 19281 11268 19303 11302
rect 19303 11268 19315 11302
rect 19353 11268 19371 11302
rect 19371 11268 19387 11302
rect 19425 11268 19439 11302
rect 19439 11268 19459 11302
rect 19497 11268 19507 11302
rect 19507 11268 19531 11302
rect 17478 11166 17512 11178
rect 17478 11144 17512 11166
rect 17478 11098 17512 11106
rect 17478 11072 17512 11098
rect 17478 11030 17512 11034
rect 17478 11000 17512 11030
rect 17478 10928 17512 10962
rect 17478 10860 17512 10890
rect 17478 10856 17512 10860
rect 17478 10792 17512 10818
rect 17478 10784 17512 10792
rect 17478 10724 17512 10746
rect 17478 10712 17512 10724
rect 17478 10656 17512 10674
rect 17478 10640 17512 10656
rect 17478 10588 17512 10602
rect 17478 10568 17512 10588
rect 17478 10520 17512 10530
rect 17478 10496 17512 10520
rect 17478 10452 17512 10458
rect 17478 10424 17512 10452
rect 17478 10384 17512 10386
rect 17478 10352 17512 10384
rect 17478 10282 17512 10314
rect 17478 10280 17512 10282
rect 17478 10214 17512 10242
rect 17478 10208 17512 10214
rect 17478 10146 17512 10170
rect 17478 10136 17512 10146
rect 17478 10078 17512 10098
rect 17478 10064 17512 10078
rect 17478 10010 17512 10026
rect 17478 9992 17512 10010
rect 17478 9942 17512 9954
rect 17478 9920 17512 9942
rect 17478 9874 17512 9882
rect 17478 9848 17512 9874
rect 17478 9806 17512 9810
rect 17478 9776 17512 9806
rect 17478 9704 17512 9738
rect 17478 9636 17512 9666
rect 17478 9632 17512 9636
rect 17478 9568 17512 9594
rect 17478 9560 17512 9568
rect 17478 9500 17512 9522
rect 17478 9488 17512 9500
rect 17478 9432 17512 9450
rect 17478 9416 17512 9432
rect 17478 9364 17512 9378
rect 17478 9344 17512 9364
rect 17478 9296 17512 9306
rect 17478 9272 17512 9296
rect 17478 9228 17512 9234
rect 17478 9200 17512 9228
rect 17478 9160 17512 9162
rect 17478 9128 17512 9160
rect 17478 9058 17512 9090
rect 17478 9056 17512 9058
rect 17478 8990 17512 9018
rect 17478 8984 17512 8990
rect 17478 8922 17512 8946
rect 17478 8912 17512 8922
rect 17478 8854 17512 8874
rect 17478 8840 17512 8854
rect 17478 8786 17512 8802
rect 17478 8768 17512 8786
rect 17478 8718 17512 8730
rect 17478 8696 17512 8718
rect 17478 8650 17512 8658
rect 17478 8624 17512 8650
rect 17478 8582 17512 8586
rect 17478 8552 17512 8582
rect 17478 8480 17512 8514
rect 17478 8412 17512 8442
rect 17478 8408 17512 8412
rect 17478 8344 17512 8370
rect 17478 8336 17512 8344
rect 17478 8276 17512 8298
rect 17478 8264 17512 8276
rect 18536 11166 18570 11178
rect 18536 11144 18570 11166
rect 18536 11098 18570 11106
rect 18536 11072 18570 11098
rect 18536 11030 18570 11034
rect 18536 11000 18570 11030
rect 18536 10928 18570 10962
rect 18536 10860 18570 10890
rect 18536 10856 18570 10860
rect 18536 10792 18570 10818
rect 18536 10784 18570 10792
rect 18536 10724 18570 10746
rect 18536 10712 18570 10724
rect 18536 10656 18570 10674
rect 18536 10640 18570 10656
rect 18536 10588 18570 10602
rect 18536 10568 18570 10588
rect 18536 10520 18570 10530
rect 18536 10496 18570 10520
rect 18536 10452 18570 10458
rect 18536 10424 18570 10452
rect 18536 10384 18570 10386
rect 18536 10352 18570 10384
rect 18536 10282 18570 10314
rect 18536 10280 18570 10282
rect 18536 10214 18570 10242
rect 18536 10208 18570 10214
rect 18536 10146 18570 10170
rect 18536 10136 18570 10146
rect 18536 10078 18570 10098
rect 18536 10064 18570 10078
rect 18536 10010 18570 10026
rect 18536 9992 18570 10010
rect 18536 9942 18570 9954
rect 18536 9920 18570 9942
rect 18536 9874 18570 9882
rect 18536 9848 18570 9874
rect 18536 9806 18570 9810
rect 18536 9776 18570 9806
rect 18536 9704 18570 9738
rect 18536 9636 18570 9666
rect 18536 9632 18570 9636
rect 18536 9568 18570 9594
rect 18536 9560 18570 9568
rect 18536 9500 18570 9522
rect 18536 9488 18570 9500
rect 18536 9432 18570 9450
rect 18536 9416 18570 9432
rect 18536 9364 18570 9378
rect 18536 9344 18570 9364
rect 18536 9296 18570 9306
rect 18536 9272 18570 9296
rect 18536 9228 18570 9234
rect 18536 9200 18570 9228
rect 18536 9160 18570 9162
rect 18536 9128 18570 9160
rect 18536 9058 18570 9090
rect 18536 9056 18570 9058
rect 18536 8990 18570 9018
rect 18536 8984 18570 8990
rect 18536 8922 18570 8946
rect 18536 8912 18570 8922
rect 18536 8854 18570 8874
rect 18536 8840 18570 8854
rect 18536 8786 18570 8802
rect 18536 8768 18570 8786
rect 18536 8718 18570 8730
rect 18536 8696 18570 8718
rect 18536 8650 18570 8658
rect 18536 8624 18570 8650
rect 18536 8582 18570 8586
rect 18536 8552 18570 8582
rect 18536 8480 18570 8514
rect 18536 8412 18570 8442
rect 18536 8408 18570 8412
rect 18536 8344 18570 8370
rect 18536 8336 18570 8344
rect 18536 8276 18570 8298
rect 18536 8264 18570 8276
rect 19594 11166 19628 11178
rect 19594 11144 19628 11166
rect 19594 11098 19628 11106
rect 19594 11072 19628 11098
rect 19594 11030 19628 11034
rect 19594 11000 19628 11030
rect 19594 10928 19628 10962
rect 19594 10860 19628 10890
rect 19594 10856 19628 10860
rect 19594 10792 19628 10818
rect 19594 10784 19628 10792
rect 19594 10724 19628 10746
rect 19594 10712 19628 10724
rect 19594 10656 19628 10674
rect 19594 10640 19628 10656
rect 19594 10588 19628 10602
rect 19594 10568 19628 10588
rect 19594 10520 19628 10530
rect 19594 10496 19628 10520
rect 19594 10452 19628 10458
rect 19594 10424 19628 10452
rect 19594 10384 19628 10386
rect 19594 10352 19628 10384
rect 19594 10282 19628 10314
rect 19594 10280 19628 10282
rect 19594 10214 19628 10242
rect 19594 10208 19628 10214
rect 19594 10146 19628 10170
rect 19594 10136 19628 10146
rect 19594 10078 19628 10098
rect 19594 10064 19628 10078
rect 19594 10010 19628 10026
rect 19594 9992 19628 10010
rect 19594 9942 19628 9954
rect 19594 9920 19628 9942
rect 19594 9874 19628 9882
rect 19594 9848 19628 9874
rect 19594 9806 19628 9810
rect 19594 9776 19628 9806
rect 19594 9704 19628 9738
rect 19594 9636 19628 9666
rect 19594 9632 19628 9636
rect 19594 9568 19628 9594
rect 19594 9560 19628 9568
rect 19594 9500 19628 9522
rect 19594 9488 19628 9500
rect 19594 9432 19628 9450
rect 19594 9416 19628 9432
rect 19594 9364 19628 9378
rect 19594 9344 19628 9364
rect 19594 9296 19628 9306
rect 19594 9272 19628 9296
rect 19594 9228 19628 9234
rect 19594 9200 19628 9228
rect 19594 9160 19628 9162
rect 19594 9128 19628 9160
rect 19594 9058 19628 9090
rect 19594 9056 19628 9058
rect 19594 8990 19628 9018
rect 19594 8984 19628 8990
rect 19594 8922 19628 8946
rect 19594 8912 19628 8922
rect 19594 8854 19628 8874
rect 19594 8840 19628 8854
rect 19594 8786 19628 8802
rect 19594 8768 19628 8786
rect 19594 8718 19628 8730
rect 19594 8696 19628 8718
rect 19594 8650 19628 8658
rect 19594 8624 19628 8650
rect 19594 8582 19628 8586
rect 19594 8552 19628 8582
rect 19594 8480 19628 8514
rect 19594 8412 19628 8442
rect 19594 8408 19628 8412
rect 19594 8344 19628 8370
rect 19594 8336 19628 8344
rect 19594 8276 19628 8298
rect 19594 8264 19628 8276
rect 17575 8140 17599 8174
rect 17599 8140 17609 8174
rect 17647 8140 17667 8174
rect 17667 8140 17681 8174
rect 17719 8140 17735 8174
rect 17735 8140 17753 8174
rect 17791 8140 17803 8174
rect 17803 8140 17825 8174
rect 17863 8140 17871 8174
rect 17871 8140 17897 8174
rect 17935 8140 17939 8174
rect 17939 8140 17969 8174
rect 18007 8140 18041 8174
rect 18079 8140 18109 8174
rect 18109 8140 18113 8174
rect 18151 8140 18177 8174
rect 18177 8140 18185 8174
rect 18223 8140 18245 8174
rect 18245 8140 18257 8174
rect 18295 8140 18313 8174
rect 18313 8140 18329 8174
rect 18367 8140 18381 8174
rect 18381 8140 18401 8174
rect 18439 8140 18449 8174
rect 18449 8140 18473 8174
rect 18633 8140 18657 8174
rect 18657 8140 18667 8174
rect 18705 8140 18725 8174
rect 18725 8140 18739 8174
rect 18777 8140 18793 8174
rect 18793 8140 18811 8174
rect 18849 8140 18861 8174
rect 18861 8140 18883 8174
rect 18921 8140 18929 8174
rect 18929 8140 18955 8174
rect 18993 8140 18997 8174
rect 18997 8140 19027 8174
rect 19065 8140 19099 8174
rect 19137 8140 19167 8174
rect 19167 8140 19171 8174
rect 19209 8140 19235 8174
rect 19235 8140 19243 8174
rect 19281 8140 19303 8174
rect 19303 8140 19315 8174
rect 19353 8140 19371 8174
rect 19371 8140 19387 8174
rect 19425 8140 19439 8174
rect 19439 8140 19459 8174
rect 19497 8140 19507 8174
rect 19507 8140 19531 8174
rect 17531 7586 17555 7620
rect 17555 7586 17565 7620
rect 17603 7586 17623 7620
rect 17623 7586 17637 7620
rect 17675 7586 17691 7620
rect 17691 7586 17709 7620
rect 17747 7586 17759 7620
rect 17759 7586 17781 7620
rect 17819 7586 17827 7620
rect 17827 7586 17853 7620
rect 17891 7586 17895 7620
rect 17895 7586 17925 7620
rect 17963 7586 17997 7620
rect 18035 7586 18065 7620
rect 18065 7586 18069 7620
rect 18107 7586 18133 7620
rect 18133 7586 18141 7620
rect 18179 7586 18201 7620
rect 18201 7586 18213 7620
rect 18251 7586 18269 7620
rect 18269 7586 18285 7620
rect 18323 7586 18337 7620
rect 18337 7586 18357 7620
rect 18395 7586 18405 7620
rect 18405 7586 18429 7620
rect 13142 6694 13164 6700
rect 13164 6694 13176 6700
rect 13242 6694 13254 6700
rect 13254 6694 13276 6700
rect 13342 6694 13344 6700
rect 13344 6694 13376 6700
rect 13142 6666 13176 6694
rect 13242 6666 13276 6694
rect 13342 6666 13376 6694
rect 13442 6666 13476 6700
rect 13542 6666 13576 6700
rect 13642 6694 13670 6700
rect 13670 6694 13676 6700
rect 13642 6666 13676 6694
rect 13142 6566 13176 6600
rect 13242 6566 13276 6600
rect 13342 6566 13376 6600
rect 13442 6566 13476 6600
rect 13542 6566 13576 6600
rect 13642 6566 13676 6600
rect 13142 6466 13176 6500
rect 13242 6466 13276 6500
rect 13342 6466 13376 6500
rect 13442 6466 13476 6500
rect 13542 6466 13576 6500
rect 13642 6466 13676 6500
rect 13142 6368 13176 6400
rect 13242 6368 13276 6400
rect 13342 6368 13376 6400
rect 13142 6366 13164 6368
rect 13164 6366 13176 6368
rect 13242 6366 13254 6368
rect 13254 6366 13276 6368
rect 13342 6366 13344 6368
rect 13344 6366 13376 6368
rect 13442 6366 13476 6400
rect 13542 6366 13576 6400
rect 13642 6368 13676 6400
rect 13642 6366 13670 6368
rect 13670 6366 13676 6368
rect 13142 6278 13176 6300
rect 13242 6278 13276 6300
rect 13342 6278 13376 6300
rect 13142 6266 13164 6278
rect 13164 6266 13176 6278
rect 13242 6266 13254 6278
rect 13254 6266 13276 6278
rect 13342 6266 13344 6278
rect 13344 6266 13376 6278
rect 13442 6266 13476 6300
rect 13542 6266 13576 6300
rect 13642 6278 13676 6300
rect 13642 6266 13670 6278
rect 13670 6266 13676 6278
rect 13142 6188 13176 6200
rect 13242 6188 13276 6200
rect 13342 6188 13376 6200
rect 13142 6166 13164 6188
rect 13164 6166 13176 6188
rect 13242 6166 13254 6188
rect 13254 6166 13276 6188
rect 13342 6166 13344 6188
rect 13344 6166 13376 6188
rect 13442 6166 13476 6200
rect 13542 6166 13576 6200
rect 13642 6188 13676 6200
rect 13642 6166 13670 6188
rect 13670 6166 13676 6188
rect 14792 6724 14814 6730
rect 14814 6724 14826 6730
rect 14892 6724 14904 6730
rect 14904 6724 14926 6730
rect 14992 6724 14994 6730
rect 14994 6724 15026 6730
rect 14792 6696 14826 6724
rect 14892 6696 14926 6724
rect 14992 6696 15026 6724
rect 15092 6696 15126 6730
rect 15192 6696 15226 6730
rect 15292 6724 15320 6730
rect 15320 6724 15326 6730
rect 15292 6696 15326 6724
rect 14792 6596 14826 6630
rect 14892 6596 14926 6630
rect 14992 6596 15026 6630
rect 15092 6596 15126 6630
rect 15192 6596 15226 6630
rect 15292 6596 15326 6630
rect 14792 6496 14826 6530
rect 14892 6496 14926 6530
rect 14992 6496 15026 6530
rect 15092 6496 15126 6530
rect 15192 6496 15226 6530
rect 15292 6496 15326 6530
rect 14792 6398 14826 6430
rect 14892 6398 14926 6430
rect 14992 6398 15026 6430
rect 14792 6396 14814 6398
rect 14814 6396 14826 6398
rect 14892 6396 14904 6398
rect 14904 6396 14926 6398
rect 14992 6396 14994 6398
rect 14994 6396 15026 6398
rect 15092 6396 15126 6430
rect 15192 6396 15226 6430
rect 15292 6398 15326 6430
rect 15292 6396 15320 6398
rect 15320 6396 15326 6398
rect 14792 6308 14826 6330
rect 14892 6308 14926 6330
rect 14992 6308 15026 6330
rect 14792 6296 14814 6308
rect 14814 6296 14826 6308
rect 14892 6296 14904 6308
rect 14904 6296 14926 6308
rect 14992 6296 14994 6308
rect 14994 6296 15026 6308
rect 15092 6296 15126 6330
rect 15192 6296 15226 6330
rect 15292 6308 15326 6330
rect 15292 6296 15320 6308
rect 15320 6296 15326 6308
rect 14792 6218 14826 6230
rect 14892 6218 14926 6230
rect 14992 6218 15026 6230
rect 14792 6196 14814 6218
rect 14814 6196 14826 6218
rect 14892 6196 14904 6218
rect 14904 6196 14926 6218
rect 14992 6196 14994 6218
rect 14994 6196 15026 6218
rect 15092 6196 15126 6230
rect 15192 6196 15226 6230
rect 15292 6218 15326 6230
rect 15292 6196 15320 6218
rect 15320 6196 15326 6218
rect 16228 7056 16262 7090
rect 16228 6984 16262 7018
rect 16228 6912 16262 6946
rect 16228 6840 16262 6874
rect 16228 6768 16262 6802
rect 16228 6696 16262 6730
rect 16546 7056 16580 7090
rect 16546 6984 16580 7018
rect 16546 6912 16580 6946
rect 16546 6840 16580 6874
rect 16546 6768 16580 6802
rect 16546 6696 16580 6730
rect 16864 7056 16898 7090
rect 16864 6984 16898 7018
rect 16864 6912 16898 6946
rect 16864 6840 16898 6874
rect 16864 6768 16898 6802
rect 16864 6696 16898 6730
rect 13142 5344 13164 5350
rect 13164 5344 13176 5350
rect 13242 5344 13254 5350
rect 13254 5344 13276 5350
rect 13342 5344 13344 5350
rect 13344 5344 13376 5350
rect 13142 5316 13176 5344
rect 13242 5316 13276 5344
rect 13342 5316 13376 5344
rect 13442 5316 13476 5350
rect 13542 5316 13576 5350
rect 13642 5344 13670 5350
rect 13670 5344 13676 5350
rect 13642 5316 13676 5344
rect 13142 5216 13176 5250
rect 13242 5216 13276 5250
rect 13342 5216 13376 5250
rect 13442 5216 13476 5250
rect 13542 5216 13576 5250
rect 13642 5216 13676 5250
rect 13142 5116 13176 5150
rect 13242 5116 13276 5150
rect 13342 5116 13376 5150
rect 13442 5116 13476 5150
rect 13542 5116 13576 5150
rect 13642 5116 13676 5150
rect 13142 5018 13176 5050
rect 13242 5018 13276 5050
rect 13342 5018 13376 5050
rect 13142 5016 13164 5018
rect 13164 5016 13176 5018
rect 13242 5016 13254 5018
rect 13254 5016 13276 5018
rect 13342 5016 13344 5018
rect 13344 5016 13376 5018
rect 13442 5016 13476 5050
rect 13542 5016 13576 5050
rect 13642 5018 13676 5050
rect 13642 5016 13670 5018
rect 13670 5016 13676 5018
rect 13142 4928 13176 4950
rect 13242 4928 13276 4950
rect 13342 4928 13376 4950
rect 13142 4916 13164 4928
rect 13164 4916 13176 4928
rect 13242 4916 13254 4928
rect 13254 4916 13276 4928
rect 13342 4916 13344 4928
rect 13344 4916 13376 4928
rect 13442 4916 13476 4950
rect 13542 4916 13576 4950
rect 13642 4928 13676 4950
rect 13642 4916 13670 4928
rect 13670 4916 13676 4928
rect 13142 4838 13176 4850
rect 13242 4838 13276 4850
rect 13342 4838 13376 4850
rect 13142 4816 13164 4838
rect 13164 4816 13176 4838
rect 13242 4816 13254 4838
rect 13254 4816 13276 4838
rect 13342 4816 13344 4838
rect 13344 4816 13376 4838
rect 13442 4816 13476 4850
rect 13542 4816 13576 4850
rect 13642 4838 13676 4850
rect 13642 4816 13670 4838
rect 13670 4816 13676 4838
rect 14792 5364 14814 5370
rect 14814 5364 14826 5370
rect 14892 5364 14904 5370
rect 14904 5364 14926 5370
rect 14992 5364 14994 5370
rect 14994 5364 15026 5370
rect 14792 5336 14826 5364
rect 14892 5336 14926 5364
rect 14992 5336 15026 5364
rect 15092 5336 15126 5370
rect 15192 5336 15226 5370
rect 15292 5364 15320 5370
rect 15320 5364 15326 5370
rect 15292 5336 15326 5364
rect 14792 5236 14826 5270
rect 14892 5236 14926 5270
rect 14992 5236 15026 5270
rect 15092 5236 15126 5270
rect 15192 5236 15226 5270
rect 15292 5236 15326 5270
rect 14792 5136 14826 5170
rect 14892 5136 14926 5170
rect 14992 5136 15026 5170
rect 15092 5136 15126 5170
rect 15192 5136 15226 5170
rect 15292 5136 15326 5170
rect 14792 5038 14826 5070
rect 14892 5038 14926 5070
rect 14992 5038 15026 5070
rect 14792 5036 14814 5038
rect 14814 5036 14826 5038
rect 14892 5036 14904 5038
rect 14904 5036 14926 5038
rect 14992 5036 14994 5038
rect 14994 5036 15026 5038
rect 15092 5036 15126 5070
rect 15192 5036 15226 5070
rect 15292 5038 15326 5070
rect 15292 5036 15320 5038
rect 15320 5036 15326 5038
rect 14792 4948 14826 4970
rect 14892 4948 14926 4970
rect 14992 4948 15026 4970
rect 14792 4936 14814 4948
rect 14814 4936 14826 4948
rect 14892 4936 14904 4948
rect 14904 4936 14926 4948
rect 14992 4936 14994 4948
rect 14994 4936 15026 4948
rect 15092 4936 15126 4970
rect 15192 4936 15226 4970
rect 15292 4948 15326 4970
rect 15292 4936 15320 4948
rect 15320 4936 15326 4948
rect 14792 4858 14826 4870
rect 14892 4858 14926 4870
rect 14992 4858 15026 4870
rect 14792 4836 14814 4858
rect 14814 4836 14826 4858
rect 14892 4836 14904 4858
rect 14904 4836 14926 4858
rect 14992 4836 14994 4858
rect 14994 4836 15026 4858
rect 15092 4836 15126 4870
rect 15192 4836 15226 4870
rect 15292 4858 15326 4870
rect 15292 4836 15320 4858
rect 15320 4836 15326 4858
rect 16228 5025 16262 5059
rect 16228 4953 16262 4987
rect 16228 4881 16262 4915
rect 16228 4809 16262 4843
rect 16228 4737 16262 4771
rect 16228 4665 16262 4699
rect 16546 5025 16580 5059
rect 16546 4953 16580 4987
rect 16546 4881 16580 4915
rect 16546 4809 16580 4843
rect 16546 4737 16580 4771
rect 16546 4665 16580 4699
rect 16864 5025 16898 5059
rect 16864 4953 16898 4987
rect 16864 4881 16898 4915
rect 16864 4809 16898 4843
rect 16864 4737 16898 4771
rect 16864 4665 16898 4699
rect 17434 7493 17468 7505
rect 17434 7471 17468 7493
rect 17434 7425 17468 7433
rect 17434 7399 17468 7425
rect 17434 7357 17468 7361
rect 17434 7327 17468 7357
rect 17434 7255 17468 7289
rect 17434 7187 17468 7217
rect 17434 7183 17468 7187
rect 17434 7119 17468 7145
rect 17434 7111 17468 7119
rect 17434 7051 17468 7073
rect 17434 7039 17468 7051
rect 17434 6983 17468 7001
rect 17434 6967 17468 6983
rect 17434 6915 17468 6929
rect 17434 6895 17468 6915
rect 17434 6847 17468 6857
rect 17434 6823 17468 6847
rect 17434 6779 17468 6785
rect 17434 6751 17468 6779
rect 17434 6711 17468 6713
rect 17434 6679 17468 6711
rect 17434 6609 17468 6641
rect 17434 6607 17468 6609
rect 17434 6541 17468 6569
rect 17434 6535 17468 6541
rect 17434 6473 17468 6497
rect 17434 6463 17468 6473
rect 17434 6405 17468 6425
rect 17434 6391 17468 6405
rect 17434 6337 17468 6353
rect 17434 6319 17468 6337
rect 17434 6269 17468 6281
rect 17434 6247 17468 6269
rect 17434 6201 17468 6209
rect 17434 6175 17468 6201
rect 17434 6133 17468 6137
rect 17434 6103 17468 6133
rect 17434 6031 17468 6065
rect 17434 5963 17468 5993
rect 17434 5959 17468 5963
rect 17434 5895 17468 5921
rect 17434 5887 17468 5895
rect 17434 5827 17468 5849
rect 17434 5815 17468 5827
rect 17434 5759 17468 5777
rect 17434 5743 17468 5759
rect 17434 5691 17468 5705
rect 17434 5671 17468 5691
rect 17434 5623 17468 5633
rect 17434 5599 17468 5623
rect 17434 5555 17468 5561
rect 17434 5527 17468 5555
rect 17434 5487 17468 5489
rect 17434 5455 17468 5487
rect 17434 5385 17468 5417
rect 17434 5383 17468 5385
rect 17434 5317 17468 5345
rect 17434 5311 17468 5317
rect 17434 5249 17468 5273
rect 17434 5239 17468 5249
rect 17434 5181 17468 5201
rect 17434 5167 17468 5181
rect 17434 5113 17468 5129
rect 17434 5095 17468 5113
rect 17434 5045 17468 5057
rect 17434 5023 17468 5045
rect 17434 4977 17468 4985
rect 17434 4951 17468 4977
rect 17434 4909 17468 4913
rect 17434 4879 17468 4909
rect 17434 4807 17468 4841
rect 17434 4739 17468 4769
rect 17434 4735 17468 4739
rect 17434 4671 17468 4697
rect 17434 4663 17468 4671
rect 17434 4603 17468 4625
rect 17434 4591 17468 4603
rect 18492 7493 18526 7505
rect 18492 7471 18526 7493
rect 18492 7425 18526 7433
rect 18492 7399 18526 7425
rect 18492 7357 18526 7361
rect 18492 7327 18526 7357
rect 18492 7255 18526 7289
rect 18492 7187 18526 7217
rect 18492 7183 18526 7187
rect 18492 7119 18526 7145
rect 18492 7111 18526 7119
rect 18492 7051 18526 7073
rect 18492 7039 18526 7051
rect 18492 6983 18526 7001
rect 18492 6967 18526 6983
rect 18492 6915 18526 6929
rect 18492 6895 18526 6915
rect 18492 6847 18526 6857
rect 18492 6823 18526 6847
rect 18492 6779 18526 6785
rect 18492 6751 18526 6779
rect 18492 6711 18526 6713
rect 18492 6679 18526 6711
rect 18492 6609 18526 6641
rect 18492 6607 18526 6609
rect 18492 6541 18526 6569
rect 18492 6535 18526 6541
rect 18492 6473 18526 6497
rect 18492 6463 18526 6473
rect 18492 6405 18526 6425
rect 18492 6391 18526 6405
rect 18492 6337 18526 6353
rect 18492 6319 18526 6337
rect 18492 6269 18526 6281
rect 18492 6247 18526 6269
rect 18492 6201 18526 6209
rect 18492 6175 18526 6201
rect 18492 6133 18526 6137
rect 18492 6103 18526 6133
rect 18492 6031 18526 6065
rect 18492 5963 18526 5993
rect 18492 5959 18526 5963
rect 18492 5895 18526 5921
rect 18492 5887 18526 5895
rect 18492 5827 18526 5849
rect 18492 5815 18526 5827
rect 18492 5759 18526 5777
rect 18492 5743 18526 5759
rect 18492 5691 18526 5705
rect 18492 5671 18526 5691
rect 18492 5623 18526 5633
rect 18492 5599 18526 5623
rect 18492 5555 18526 5561
rect 18492 5527 18526 5555
rect 18492 5487 18526 5489
rect 18492 5455 18526 5487
rect 18492 5385 18526 5417
rect 18492 5383 18526 5385
rect 18492 5317 18526 5345
rect 18492 5311 18526 5317
rect 18492 5249 18526 5273
rect 18492 5239 18526 5249
rect 18492 5181 18526 5201
rect 18492 5167 18526 5181
rect 18492 5113 18526 5129
rect 18492 5095 18526 5113
rect 18492 5045 18526 5057
rect 18492 5023 18526 5045
rect 18492 4977 18526 4985
rect 18492 4951 18526 4977
rect 18492 4909 18526 4913
rect 18492 4879 18526 4909
rect 18492 4807 18526 4841
rect 18492 4739 18526 4769
rect 18492 4735 18526 4739
rect 18492 4671 18526 4697
rect 18492 4663 18526 4671
rect 18492 4603 18526 4625
rect 18492 4591 18526 4603
rect 17531 4476 17555 4510
rect 17555 4476 17565 4510
rect 17603 4476 17623 4510
rect 17623 4476 17637 4510
rect 17675 4476 17691 4510
rect 17691 4476 17709 4510
rect 17747 4476 17759 4510
rect 17759 4476 17781 4510
rect 17819 4476 17827 4510
rect 17827 4476 17853 4510
rect 17891 4476 17895 4510
rect 17895 4476 17925 4510
rect 17963 4476 17997 4510
rect 18035 4476 18065 4510
rect 18065 4476 18069 4510
rect 18107 4476 18133 4510
rect 18133 4476 18141 4510
rect 18179 4476 18201 4510
rect 18201 4476 18213 4510
rect 18251 4476 18269 4510
rect 18269 4476 18285 4510
rect 18323 4476 18337 4510
rect 18337 4476 18357 4510
rect 18395 4476 18405 4510
rect 18405 4476 18429 4510
rect 18981 7586 19005 7620
rect 19005 7586 19015 7620
rect 19053 7586 19073 7620
rect 19073 7586 19087 7620
rect 19125 7586 19141 7620
rect 19141 7586 19159 7620
rect 19197 7586 19209 7620
rect 19209 7586 19231 7620
rect 19269 7586 19277 7620
rect 19277 7586 19303 7620
rect 19341 7586 19345 7620
rect 19345 7586 19375 7620
rect 19413 7586 19447 7620
rect 19485 7586 19515 7620
rect 19515 7586 19519 7620
rect 19557 7586 19583 7620
rect 19583 7586 19591 7620
rect 19629 7586 19651 7620
rect 19651 7586 19663 7620
rect 19701 7586 19719 7620
rect 19719 7586 19735 7620
rect 19773 7586 19787 7620
rect 19787 7586 19807 7620
rect 19845 7586 19855 7620
rect 19855 7586 19879 7620
rect 18884 7493 18918 7505
rect 18884 7471 18918 7493
rect 18884 7425 18918 7433
rect 18884 7399 18918 7425
rect 18884 7357 18918 7361
rect 18884 7327 18918 7357
rect 18884 7255 18918 7289
rect 18884 7187 18918 7217
rect 18884 7183 18918 7187
rect 18884 7119 18918 7145
rect 18884 7111 18918 7119
rect 18884 7051 18918 7073
rect 18884 7039 18918 7051
rect 18884 6983 18918 7001
rect 18884 6967 18918 6983
rect 18884 6915 18918 6929
rect 18884 6895 18918 6915
rect 18884 6847 18918 6857
rect 18884 6823 18918 6847
rect 18884 6779 18918 6785
rect 18884 6751 18918 6779
rect 18884 6711 18918 6713
rect 18884 6679 18918 6711
rect 18884 6609 18918 6641
rect 18884 6607 18918 6609
rect 18884 6541 18918 6569
rect 18884 6535 18918 6541
rect 18884 6473 18918 6497
rect 18884 6463 18918 6473
rect 18884 6405 18918 6425
rect 18884 6391 18918 6405
rect 18884 6337 18918 6353
rect 18884 6319 18918 6337
rect 18884 6269 18918 6281
rect 18884 6247 18918 6269
rect 18884 6201 18918 6209
rect 18884 6175 18918 6201
rect 18884 6133 18918 6137
rect 18884 6103 18918 6133
rect 18884 6031 18918 6065
rect 18884 5963 18918 5993
rect 18884 5959 18918 5963
rect 18884 5895 18918 5921
rect 18884 5887 18918 5895
rect 18884 5827 18918 5849
rect 18884 5815 18918 5827
rect 18884 5759 18918 5777
rect 18884 5743 18918 5759
rect 18884 5691 18918 5705
rect 18884 5671 18918 5691
rect 18884 5623 18918 5633
rect 18884 5599 18918 5623
rect 18884 5555 18918 5561
rect 18884 5527 18918 5555
rect 18884 5487 18918 5489
rect 18884 5455 18918 5487
rect 18884 5385 18918 5417
rect 18884 5383 18918 5385
rect 18884 5317 18918 5345
rect 18884 5311 18918 5317
rect 18884 5249 18918 5273
rect 18884 5239 18918 5249
rect 18884 5181 18918 5201
rect 18884 5167 18918 5181
rect 18884 5113 18918 5129
rect 18884 5095 18918 5113
rect 18884 5045 18918 5057
rect 18884 5023 18918 5045
rect 18884 4977 18918 4985
rect 18884 4951 18918 4977
rect 18884 4909 18918 4913
rect 18884 4879 18918 4909
rect 18884 4807 18918 4841
rect 18884 4739 18918 4769
rect 18884 4735 18918 4739
rect 18884 4671 18918 4697
rect 18884 4663 18918 4671
rect 18884 4603 18918 4625
rect 18884 4591 18918 4603
rect 19942 7493 19976 7505
rect 19942 7471 19976 7493
rect 19942 7425 19976 7433
rect 19942 7399 19976 7425
rect 19942 7357 19976 7361
rect 19942 7327 19976 7357
rect 19942 7255 19976 7289
rect 19942 7187 19976 7217
rect 19942 7183 19976 7187
rect 19942 7119 19976 7145
rect 19942 7111 19976 7119
rect 19942 7051 19976 7073
rect 19942 7039 19976 7051
rect 19942 6983 19976 7001
rect 19942 6967 19976 6983
rect 19942 6915 19976 6929
rect 19942 6895 19976 6915
rect 19942 6847 19976 6857
rect 19942 6823 19976 6847
rect 19942 6779 19976 6785
rect 19942 6751 19976 6779
rect 19942 6711 19976 6713
rect 19942 6679 19976 6711
rect 19942 6609 19976 6641
rect 19942 6607 19976 6609
rect 19942 6541 19976 6569
rect 19942 6535 19976 6541
rect 19942 6473 19976 6497
rect 19942 6463 19976 6473
rect 19942 6405 19976 6425
rect 19942 6391 19976 6405
rect 19942 6337 19976 6353
rect 19942 6319 19976 6337
rect 19942 6269 19976 6281
rect 19942 6247 19976 6269
rect 19942 6201 19976 6209
rect 19942 6175 19976 6201
rect 19942 6133 19976 6137
rect 19942 6103 19976 6133
rect 19942 6031 19976 6065
rect 19942 5963 19976 5993
rect 19942 5959 19976 5963
rect 19942 5895 19976 5921
rect 19942 5887 19976 5895
rect 19942 5827 19976 5849
rect 19942 5815 19976 5827
rect 19942 5759 19976 5777
rect 19942 5743 19976 5759
rect 19942 5691 19976 5705
rect 19942 5671 19976 5691
rect 19942 5623 19976 5633
rect 19942 5599 19976 5623
rect 19942 5555 19976 5561
rect 19942 5527 19976 5555
rect 19942 5487 19976 5489
rect 19942 5455 19976 5487
rect 19942 5385 19976 5417
rect 19942 5383 19976 5385
rect 19942 5317 19976 5345
rect 19942 5311 19976 5317
rect 19942 5249 19976 5273
rect 19942 5239 19976 5249
rect 19942 5181 19976 5201
rect 19942 5167 19976 5181
rect 19942 5113 19976 5129
rect 19942 5095 19976 5113
rect 19942 5045 19976 5057
rect 19942 5023 19976 5045
rect 19942 4977 19976 4985
rect 19942 4951 19976 4977
rect 19942 4909 19976 4913
rect 19942 4879 19976 4909
rect 19942 4807 19976 4841
rect 19942 4739 19976 4769
rect 19942 4735 19976 4739
rect 19942 4671 19976 4697
rect 19942 4663 19976 4671
rect 19942 4603 19976 4625
rect 19942 4591 19976 4603
rect 23480 15462 23502 15468
rect 23502 15462 23514 15468
rect 23580 15462 23592 15468
rect 23592 15462 23614 15468
rect 23680 15462 23682 15468
rect 23682 15462 23714 15468
rect 23480 15434 23514 15462
rect 23580 15434 23614 15462
rect 23680 15434 23714 15462
rect 23780 15434 23814 15468
rect 23880 15434 23914 15468
rect 23980 15462 24008 15468
rect 24008 15462 24014 15468
rect 23980 15434 24014 15462
rect 23480 15334 23514 15368
rect 23580 15334 23614 15368
rect 23680 15334 23714 15368
rect 23780 15334 23814 15368
rect 23880 15334 23914 15368
rect 23980 15334 24014 15368
rect 24609 15614 24643 15648
rect 24681 15614 24715 15648
rect 24753 15614 24787 15648
rect 24825 15614 24859 15648
rect 24897 15614 24931 15648
rect 24969 15614 25003 15648
rect 27140 15614 27174 15648
rect 27212 15614 27246 15648
rect 27284 15614 27318 15648
rect 27356 15614 27390 15648
rect 27428 15614 27462 15648
rect 27500 15614 27534 15648
rect 23480 15234 23514 15268
rect 23580 15234 23614 15268
rect 23680 15234 23714 15268
rect 23780 15234 23814 15268
rect 23880 15234 23914 15268
rect 23980 15234 24014 15268
rect 23480 15136 23514 15168
rect 23580 15136 23614 15168
rect 23680 15136 23714 15168
rect 23480 15134 23502 15136
rect 23502 15134 23514 15136
rect 23580 15134 23592 15136
rect 23592 15134 23614 15136
rect 23680 15134 23682 15136
rect 23682 15134 23714 15136
rect 23780 15134 23814 15168
rect 23880 15134 23914 15168
rect 23980 15136 24014 15168
rect 38517 15807 38767 15913
rect 39533 15806 39855 15912
rect 40586 15887 40620 15921
rect 40586 15815 40620 15849
rect 24609 15296 24643 15330
rect 24681 15296 24715 15330
rect 24753 15296 24787 15330
rect 24825 15296 24859 15330
rect 24897 15296 24931 15330
rect 24969 15296 25003 15330
rect 27140 15296 27174 15330
rect 27212 15296 27246 15330
rect 27284 15296 27318 15330
rect 27356 15296 27390 15330
rect 27428 15296 27462 15330
rect 27500 15296 27534 15330
rect 28982 15208 29016 15242
rect 23980 15134 24008 15136
rect 24008 15134 24014 15136
rect 23480 15046 23514 15068
rect 23580 15046 23614 15068
rect 23680 15046 23714 15068
rect 23480 15034 23502 15046
rect 23502 15034 23514 15046
rect 23580 15034 23592 15046
rect 23592 15034 23614 15046
rect 23680 15034 23682 15046
rect 23682 15034 23714 15046
rect 23780 15034 23814 15068
rect 23880 15034 23914 15068
rect 23980 15046 24014 15068
rect 23980 15034 24008 15046
rect 24008 15034 24014 15046
rect 23480 14956 23514 14968
rect 23580 14956 23614 14968
rect 23680 14956 23714 14968
rect 23480 14934 23502 14956
rect 23502 14934 23514 14956
rect 23580 14934 23592 14956
rect 23592 14934 23614 14956
rect 23680 14934 23682 14956
rect 23682 14934 23714 14956
rect 23780 14934 23814 14968
rect 23880 14934 23914 14968
rect 23980 14956 24014 14968
rect 23980 14934 24008 14956
rect 24008 14934 24014 14956
rect 28982 15136 29016 15170
rect 28982 15064 29016 15098
rect 28982 14992 29016 15026
rect 28982 14920 29016 14954
rect 28982 14848 29016 14882
rect 29300 15208 29334 15242
rect 29300 15136 29334 15170
rect 29300 15064 29334 15098
rect 29300 14992 29334 15026
rect 29300 14920 29334 14954
rect 29300 14848 29334 14882
rect 29618 15208 29652 15242
rect 29618 15136 29652 15170
rect 29618 15064 29652 15098
rect 29618 14992 29652 15026
rect 29618 14920 29652 14954
rect 29618 14848 29652 14882
rect 28982 14137 29016 14171
rect 28982 14065 29016 14099
rect 28982 13993 29016 14027
rect 28982 13921 29016 13955
rect 28982 13849 29016 13883
rect 28982 13777 29016 13811
rect 29300 14137 29334 14171
rect 29300 14065 29334 14099
rect 29300 13993 29334 14027
rect 29300 13921 29334 13955
rect 29300 13849 29334 13883
rect 29300 13777 29334 13811
rect 29618 14137 29652 14171
rect 29618 14065 29652 14099
rect 29618 13993 29652 14027
rect 29618 13921 29652 13955
rect 29618 13849 29652 13883
rect 29618 13777 29652 13811
rect 38133 15520 38167 15538
rect 38133 15504 38167 15520
rect 38133 15452 38167 15466
rect 38133 15432 38167 15452
rect 38133 15384 38167 15394
rect 38133 15360 38167 15384
rect 38133 15316 38167 15322
rect 38133 15288 38167 15316
rect 38133 15248 38167 15250
rect 38133 15216 38167 15248
rect 38133 15146 38167 15178
rect 38133 15144 38167 15146
rect 38133 15078 38167 15106
rect 38133 15072 38167 15078
rect 38133 15010 38167 15034
rect 38133 15000 38167 15010
rect 38133 14942 38167 14962
rect 38133 14928 38167 14942
rect 38133 14874 38167 14890
rect 38133 14856 38167 14874
rect 38133 14806 38167 14818
rect 38133 14784 38167 14806
rect 38133 14738 38167 14746
rect 38133 14712 38167 14738
rect 38133 14670 38167 14674
rect 38133 14640 38167 14670
rect 38133 14568 38167 14602
rect 38133 14500 38167 14530
rect 38133 14496 38167 14500
rect 38133 14432 38167 14458
rect 38133 14424 38167 14432
rect 38133 14364 38167 14386
rect 38133 14352 38167 14364
rect 38133 14296 38167 14314
rect 38133 14280 38167 14296
rect 38133 14228 38167 14242
rect 38133 14208 38167 14228
rect 38133 14160 38167 14170
rect 38133 14136 38167 14160
rect 38133 14092 38167 14098
rect 38133 14064 38167 14092
rect 38133 14024 38167 14026
rect 38133 13992 38167 14024
rect 38133 13922 38167 13954
rect 38133 13920 38167 13922
rect 38133 13854 38167 13882
rect 38133 13848 38167 13854
rect 38133 13786 38167 13810
rect 38133 13776 38167 13786
rect 38133 13718 38167 13738
rect 38133 13704 38167 13718
rect 38133 13650 38167 13666
rect 38133 13632 38167 13650
rect 38391 15520 38425 15538
rect 38391 15504 38425 15520
rect 38391 15452 38425 15466
rect 38391 15432 38425 15452
rect 38391 15384 38425 15394
rect 38391 15360 38425 15384
rect 38391 15316 38425 15322
rect 38391 15288 38425 15316
rect 38391 15248 38425 15250
rect 38391 15216 38425 15248
rect 38391 15146 38425 15178
rect 38391 15144 38425 15146
rect 38391 15078 38425 15106
rect 38391 15072 38425 15078
rect 38391 15010 38425 15034
rect 38391 15000 38425 15010
rect 38391 14942 38425 14962
rect 38391 14928 38425 14942
rect 38391 14874 38425 14890
rect 38391 14856 38425 14874
rect 38391 14806 38425 14818
rect 38391 14784 38425 14806
rect 38391 14738 38425 14746
rect 38391 14712 38425 14738
rect 38391 14670 38425 14674
rect 38391 14640 38425 14670
rect 38391 14568 38425 14602
rect 38391 14500 38425 14530
rect 38391 14496 38425 14500
rect 38391 14432 38425 14458
rect 38391 14424 38425 14432
rect 38391 14364 38425 14386
rect 38391 14352 38425 14364
rect 38391 14296 38425 14314
rect 38391 14280 38425 14296
rect 38391 14228 38425 14242
rect 38391 14208 38425 14228
rect 38391 14160 38425 14170
rect 38391 14136 38425 14160
rect 38391 14092 38425 14098
rect 38391 14064 38425 14092
rect 38391 14024 38425 14026
rect 38391 13992 38425 14024
rect 38391 13922 38425 13954
rect 38391 13920 38425 13922
rect 38391 13854 38425 13882
rect 38391 13848 38425 13854
rect 38391 13786 38425 13810
rect 38391 13776 38425 13786
rect 38391 13718 38425 13738
rect 38391 13704 38425 13718
rect 38391 13650 38425 13666
rect 38391 13632 38425 13650
rect 38649 15520 38683 15538
rect 38649 15504 38683 15520
rect 38649 15452 38683 15466
rect 38649 15432 38683 15452
rect 38649 15384 38683 15394
rect 38649 15360 38683 15384
rect 38649 15316 38683 15322
rect 38649 15288 38683 15316
rect 38649 15248 38683 15250
rect 38649 15216 38683 15248
rect 38649 15146 38683 15178
rect 38649 15144 38683 15146
rect 38649 15078 38683 15106
rect 38649 15072 38683 15078
rect 38649 15010 38683 15034
rect 38649 15000 38683 15010
rect 38649 14942 38683 14962
rect 38649 14928 38683 14942
rect 38649 14874 38683 14890
rect 38649 14856 38683 14874
rect 38649 14806 38683 14818
rect 38649 14784 38683 14806
rect 38649 14738 38683 14746
rect 38649 14712 38683 14738
rect 38649 14670 38683 14674
rect 38649 14640 38683 14670
rect 38649 14568 38683 14602
rect 38649 14500 38683 14530
rect 38649 14496 38683 14500
rect 38649 14432 38683 14458
rect 38649 14424 38683 14432
rect 38649 14364 38683 14386
rect 38649 14352 38683 14364
rect 38649 14296 38683 14314
rect 38649 14280 38683 14296
rect 38649 14228 38683 14242
rect 38649 14208 38683 14228
rect 38649 14160 38683 14170
rect 38649 14136 38683 14160
rect 38649 14092 38683 14098
rect 38649 14064 38683 14092
rect 38649 14024 38683 14026
rect 38649 13992 38683 14024
rect 38649 13922 38683 13954
rect 38649 13920 38683 13922
rect 38649 13854 38683 13882
rect 38649 13848 38683 13854
rect 38649 13786 38683 13810
rect 38649 13776 38683 13786
rect 38649 13718 38683 13738
rect 38649 13704 38683 13718
rect 38649 13650 38683 13666
rect 38649 13632 38683 13650
rect 38907 15520 38941 15538
rect 38907 15504 38941 15520
rect 38907 15452 38941 15466
rect 38907 15432 38941 15452
rect 38907 15384 38941 15394
rect 38907 15360 38941 15384
rect 38907 15316 38941 15322
rect 38907 15288 38941 15316
rect 38907 15248 38941 15250
rect 38907 15216 38941 15248
rect 38907 15146 38941 15178
rect 38907 15144 38941 15146
rect 38907 15078 38941 15106
rect 38907 15072 38941 15078
rect 38907 15010 38941 15034
rect 38907 15000 38941 15010
rect 38907 14942 38941 14962
rect 38907 14928 38941 14942
rect 38907 14874 38941 14890
rect 38907 14856 38941 14874
rect 38907 14806 38941 14818
rect 38907 14784 38941 14806
rect 38907 14738 38941 14746
rect 38907 14712 38941 14738
rect 38907 14670 38941 14674
rect 38907 14640 38941 14670
rect 38907 14568 38941 14602
rect 38907 14500 38941 14530
rect 38907 14496 38941 14500
rect 38907 14432 38941 14458
rect 38907 14424 38941 14432
rect 38907 14364 38941 14386
rect 38907 14352 38941 14364
rect 38907 14296 38941 14314
rect 38907 14280 38941 14296
rect 38907 14228 38941 14242
rect 38907 14208 38941 14228
rect 38907 14160 38941 14170
rect 38907 14136 38941 14160
rect 38907 14092 38941 14098
rect 38907 14064 38941 14092
rect 38907 14024 38941 14026
rect 38907 13992 38941 14024
rect 38907 13922 38941 13954
rect 38907 13920 38941 13922
rect 38907 13854 38941 13882
rect 38907 13848 38941 13854
rect 38907 13786 38941 13810
rect 38907 13776 38941 13786
rect 38907 13718 38941 13738
rect 38907 13704 38941 13718
rect 38907 13650 38941 13666
rect 38907 13632 38941 13650
rect 39165 15520 39199 15538
rect 39165 15504 39199 15520
rect 39165 15452 39199 15466
rect 39165 15432 39199 15452
rect 39165 15384 39199 15394
rect 39165 15360 39199 15384
rect 39165 15316 39199 15322
rect 39165 15288 39199 15316
rect 39165 15248 39199 15250
rect 39165 15216 39199 15248
rect 39165 15146 39199 15178
rect 39165 15144 39199 15146
rect 39165 15078 39199 15106
rect 39165 15072 39199 15078
rect 39165 15010 39199 15034
rect 39165 15000 39199 15010
rect 39165 14942 39199 14962
rect 39165 14928 39199 14942
rect 39165 14874 39199 14890
rect 39165 14856 39199 14874
rect 39165 14806 39199 14818
rect 39165 14784 39199 14806
rect 39165 14738 39199 14746
rect 39165 14712 39199 14738
rect 39165 14670 39199 14674
rect 39165 14640 39199 14670
rect 39165 14568 39199 14602
rect 39165 14500 39199 14530
rect 39165 14496 39199 14500
rect 39165 14432 39199 14458
rect 39165 14424 39199 14432
rect 39165 14364 39199 14386
rect 39165 14352 39199 14364
rect 39165 14296 39199 14314
rect 39165 14280 39199 14296
rect 39165 14228 39199 14242
rect 39165 14208 39199 14228
rect 39165 14160 39199 14170
rect 39165 14136 39199 14160
rect 39165 14092 39199 14098
rect 39165 14064 39199 14092
rect 39165 14024 39199 14026
rect 39165 13992 39199 14024
rect 39165 13922 39199 13954
rect 39165 13920 39199 13922
rect 39165 13854 39199 13882
rect 39165 13848 39199 13854
rect 39165 13786 39199 13810
rect 39165 13776 39199 13786
rect 39165 13718 39199 13738
rect 39165 13704 39199 13718
rect 39165 13650 39199 13666
rect 39165 13632 39199 13650
rect 39423 15520 39457 15538
rect 39423 15504 39457 15520
rect 39423 15452 39457 15466
rect 39423 15432 39457 15452
rect 39423 15384 39457 15394
rect 39423 15360 39457 15384
rect 39423 15316 39457 15322
rect 39423 15288 39457 15316
rect 39423 15248 39457 15250
rect 39423 15216 39457 15248
rect 39423 15146 39457 15178
rect 39423 15144 39457 15146
rect 39423 15078 39457 15106
rect 39423 15072 39457 15078
rect 39423 15010 39457 15034
rect 39423 15000 39457 15010
rect 39423 14942 39457 14962
rect 39423 14928 39457 14942
rect 39423 14874 39457 14890
rect 39423 14856 39457 14874
rect 39423 14806 39457 14818
rect 39423 14784 39457 14806
rect 39423 14738 39457 14746
rect 39423 14712 39457 14738
rect 39423 14670 39457 14674
rect 39423 14640 39457 14670
rect 39423 14568 39457 14602
rect 39423 14500 39457 14530
rect 39423 14496 39457 14500
rect 39423 14432 39457 14458
rect 39423 14424 39457 14432
rect 39423 14364 39457 14386
rect 39423 14352 39457 14364
rect 39423 14296 39457 14314
rect 39423 14280 39457 14296
rect 39423 14228 39457 14242
rect 39423 14208 39457 14228
rect 39423 14160 39457 14170
rect 39423 14136 39457 14160
rect 39423 14092 39457 14098
rect 39423 14064 39457 14092
rect 39423 14024 39457 14026
rect 39423 13992 39457 14024
rect 39423 13922 39457 13954
rect 39423 13920 39457 13922
rect 39423 13854 39457 13882
rect 39423 13848 39457 13854
rect 39423 13786 39457 13810
rect 39423 13776 39457 13786
rect 39423 13718 39457 13738
rect 39423 13704 39457 13718
rect 39423 13650 39457 13666
rect 39423 13632 39457 13650
rect 23224 13322 23250 13356
rect 23250 13322 23258 13356
rect 23296 13322 23318 13356
rect 23318 13322 23330 13356
rect 23368 13322 23386 13356
rect 23386 13322 23402 13356
rect 23440 13322 23454 13356
rect 23454 13322 23474 13356
rect 23512 13322 23522 13356
rect 23522 13322 23546 13356
rect 23584 13322 23590 13356
rect 23590 13322 23618 13356
rect 23656 13322 23658 13356
rect 23658 13322 23690 13356
rect 23728 13322 23760 13356
rect 23760 13322 23762 13356
rect 23800 13322 23828 13356
rect 23828 13322 23834 13356
rect 23872 13322 23896 13356
rect 23896 13322 23906 13356
rect 23944 13322 23964 13356
rect 23964 13322 23978 13356
rect 24016 13322 24032 13356
rect 24032 13322 24050 13356
rect 24088 13322 24100 13356
rect 24100 13322 24122 13356
rect 24160 13322 24168 13356
rect 24168 13322 24194 13356
rect 23128 13235 23162 13259
rect 23128 13225 23162 13235
rect 23128 13167 23162 13187
rect 23128 13153 23162 13167
rect 23128 13099 23162 13115
rect 23128 13081 23162 13099
rect 23128 13031 23162 13043
rect 23128 13009 23162 13031
rect 23128 12963 23162 12971
rect 23128 12937 23162 12963
rect 23128 12895 23162 12899
rect 23128 12865 23162 12895
rect 23128 12793 23162 12827
rect 23128 12725 23162 12755
rect 23128 12721 23162 12725
rect 23128 12657 23162 12683
rect 23128 12649 23162 12657
rect 23128 12589 23162 12611
rect 23128 12577 23162 12589
rect 23128 12521 23162 12539
rect 23128 12505 23162 12521
rect 23128 12453 23162 12467
rect 23128 12433 23162 12453
rect 23128 12385 23162 12395
rect 23128 12361 23162 12385
rect 24256 13235 24290 13259
rect 24256 13225 24290 13235
rect 24256 13167 24290 13187
rect 24256 13153 24290 13167
rect 24256 13099 24290 13115
rect 24256 13081 24290 13099
rect 24256 13031 24290 13043
rect 24256 13009 24290 13031
rect 24256 12963 24290 12971
rect 24256 12937 24290 12963
rect 24256 12895 24290 12899
rect 24256 12865 24290 12895
rect 24256 12793 24290 12827
rect 24256 12725 24290 12755
rect 24256 12721 24290 12725
rect 24256 12657 24290 12683
rect 24256 12649 24290 12657
rect 24256 12589 24290 12611
rect 24256 12577 24290 12589
rect 24256 12521 24290 12539
rect 24256 12505 24290 12521
rect 24256 12453 24290 12467
rect 24256 12433 24290 12453
rect 24256 12385 24290 12395
rect 24256 12361 24290 12385
rect 23224 12264 23250 12298
rect 23250 12264 23258 12298
rect 23296 12264 23318 12298
rect 23318 12264 23330 12298
rect 23368 12264 23386 12298
rect 23386 12264 23402 12298
rect 23440 12264 23454 12298
rect 23454 12264 23474 12298
rect 23512 12264 23522 12298
rect 23522 12264 23546 12298
rect 23584 12264 23590 12298
rect 23590 12264 23618 12298
rect 23656 12264 23658 12298
rect 23658 12264 23690 12298
rect 23728 12264 23760 12298
rect 23760 12264 23762 12298
rect 23800 12264 23828 12298
rect 23828 12264 23834 12298
rect 23872 12264 23896 12298
rect 23896 12264 23906 12298
rect 23944 12264 23964 12298
rect 23964 12264 23978 12298
rect 24016 12264 24032 12298
rect 24032 12264 24050 12298
rect 24088 12264 24100 12298
rect 24100 12264 24122 12298
rect 24160 12264 24168 12298
rect 24168 12264 24194 12298
rect 24784 13316 24810 13350
rect 24810 13316 24818 13350
rect 24856 13316 24878 13350
rect 24878 13316 24890 13350
rect 24928 13316 24946 13350
rect 24946 13316 24962 13350
rect 25000 13316 25014 13350
rect 25014 13316 25034 13350
rect 25072 13316 25082 13350
rect 25082 13316 25106 13350
rect 25144 13316 25150 13350
rect 25150 13316 25178 13350
rect 25216 13316 25218 13350
rect 25218 13316 25250 13350
rect 25288 13316 25320 13350
rect 25320 13316 25322 13350
rect 25360 13316 25388 13350
rect 25388 13316 25394 13350
rect 25432 13316 25456 13350
rect 25456 13316 25466 13350
rect 25504 13316 25524 13350
rect 25524 13316 25538 13350
rect 25576 13316 25592 13350
rect 25592 13316 25610 13350
rect 25648 13316 25660 13350
rect 25660 13316 25682 13350
rect 25720 13316 25728 13350
rect 25728 13316 25754 13350
rect 24688 13229 24722 13253
rect 24688 13219 24722 13229
rect 24688 13161 24722 13181
rect 24688 13147 24722 13161
rect 24688 13093 24722 13109
rect 24688 13075 24722 13093
rect 24688 13025 24722 13037
rect 24688 13003 24722 13025
rect 24688 12957 24722 12965
rect 24688 12931 24722 12957
rect 24688 12889 24722 12893
rect 24688 12859 24722 12889
rect 24688 12787 24722 12821
rect 24688 12719 24722 12749
rect 24688 12715 24722 12719
rect 24688 12651 24722 12677
rect 24688 12643 24722 12651
rect 24688 12583 24722 12605
rect 24688 12571 24722 12583
rect 24688 12515 24722 12533
rect 24688 12499 24722 12515
rect 24688 12447 24722 12461
rect 24688 12427 24722 12447
rect 24688 12379 24722 12389
rect 24688 12355 24722 12379
rect 25816 13229 25850 13253
rect 25816 13219 25850 13229
rect 25816 13161 25850 13181
rect 25816 13147 25850 13161
rect 25816 13093 25850 13109
rect 25816 13075 25850 13093
rect 25816 13025 25850 13037
rect 25816 13003 25850 13025
rect 25816 12957 25850 12965
rect 25816 12931 25850 12957
rect 25816 12889 25850 12893
rect 25816 12859 25850 12889
rect 25816 12787 25850 12821
rect 25816 12719 25850 12749
rect 25816 12715 25850 12719
rect 25816 12651 25850 12677
rect 25816 12643 25850 12651
rect 25816 12583 25850 12605
rect 25816 12571 25850 12583
rect 25816 12515 25850 12533
rect 25816 12499 25850 12515
rect 25816 12447 25850 12461
rect 25816 12427 25850 12447
rect 25816 12379 25850 12389
rect 25816 12355 25850 12379
rect 26546 13290 26580 13324
rect 26546 13218 26580 13252
rect 26546 13146 26580 13180
rect 26546 13074 26580 13108
rect 26546 13002 26580 13036
rect 26546 12930 26580 12964
rect 26864 13290 26898 13324
rect 26864 13218 26898 13252
rect 26864 13146 26898 13180
rect 26864 13074 26898 13108
rect 26864 13002 26898 13036
rect 26864 12930 26898 12964
rect 27182 13290 27216 13324
rect 27182 13218 27216 13252
rect 27718 13274 27752 13308
rect 27182 13146 27216 13180
rect 27718 13202 27752 13236
rect 27718 13130 27752 13164
rect 27182 13074 27216 13108
rect 27718 13058 27752 13092
rect 27182 13002 27216 13036
rect 27718 12986 27752 13020
rect 27182 12930 27216 12964
rect 27718 12914 27752 12948
rect 24784 12258 24810 12292
rect 24810 12258 24818 12292
rect 24856 12258 24878 12292
rect 24878 12258 24890 12292
rect 24928 12258 24946 12292
rect 24946 12258 24962 12292
rect 25000 12258 25014 12292
rect 25014 12258 25034 12292
rect 25072 12258 25082 12292
rect 25082 12258 25106 12292
rect 25144 12258 25150 12292
rect 25150 12258 25178 12292
rect 25216 12258 25218 12292
rect 25218 12258 25250 12292
rect 25288 12258 25320 12292
rect 25320 12258 25322 12292
rect 25360 12258 25388 12292
rect 25388 12258 25394 12292
rect 25432 12258 25456 12292
rect 25456 12258 25466 12292
rect 25504 12258 25524 12292
rect 25524 12258 25538 12292
rect 25576 12258 25592 12292
rect 25592 12258 25610 12292
rect 25648 12258 25660 12292
rect 25660 12258 25682 12292
rect 25720 12258 25728 12292
rect 25728 12258 25754 12292
rect 23145 11782 23171 11816
rect 23171 11782 23179 11816
rect 23217 11782 23239 11816
rect 23239 11782 23251 11816
rect 23289 11782 23307 11816
rect 23307 11782 23323 11816
rect 23361 11782 23375 11816
rect 23375 11782 23395 11816
rect 23433 11782 23443 11816
rect 23443 11782 23467 11816
rect 23505 11782 23511 11816
rect 23511 11782 23539 11816
rect 23577 11782 23579 11816
rect 23579 11782 23611 11816
rect 23649 11782 23681 11816
rect 23681 11782 23683 11816
rect 23721 11782 23749 11816
rect 23749 11782 23755 11816
rect 23793 11782 23817 11816
rect 23817 11782 23827 11816
rect 23865 11782 23885 11816
rect 23885 11782 23899 11816
rect 23937 11782 23953 11816
rect 23953 11782 23971 11816
rect 24009 11782 24021 11816
rect 24021 11782 24043 11816
rect 24081 11782 24089 11816
rect 24089 11782 24115 11816
rect 23058 11695 23092 11719
rect 23058 11685 23092 11695
rect 23058 11627 23092 11647
rect 23058 11613 23092 11627
rect 23058 11559 23092 11575
rect 23058 11541 23092 11559
rect 23058 11491 23092 11503
rect 23058 11469 23092 11491
rect 23058 11423 23092 11431
rect 23058 11397 23092 11423
rect 23058 11355 23092 11359
rect 23058 11325 23092 11355
rect 23058 11253 23092 11287
rect 23058 11185 23092 11215
rect 23058 11181 23092 11185
rect 23058 11117 23092 11143
rect 23058 11109 23092 11117
rect 23058 11049 23092 11071
rect 23058 11037 23092 11049
rect 23058 10981 23092 10999
rect 23058 10965 23092 10981
rect 23058 10913 23092 10927
rect 23058 10893 23092 10913
rect 23058 10845 23092 10855
rect 23058 10821 23092 10845
rect 24168 11695 24202 11719
rect 24168 11685 24202 11695
rect 24168 11627 24202 11647
rect 24168 11613 24202 11627
rect 24168 11559 24202 11575
rect 24168 11541 24202 11559
rect 24168 11491 24202 11503
rect 24168 11469 24202 11491
rect 24168 11423 24202 11431
rect 24168 11397 24202 11423
rect 24168 11355 24202 11359
rect 24168 11325 24202 11355
rect 24168 11253 24202 11287
rect 24168 11185 24202 11215
rect 24168 11181 24202 11185
rect 24168 11117 24202 11143
rect 24168 11109 24202 11117
rect 24168 11049 24202 11071
rect 24168 11037 24202 11049
rect 24168 10981 24202 10999
rect 24168 10965 24202 10981
rect 24168 10913 24202 10927
rect 24168 10893 24202 10913
rect 24168 10845 24202 10855
rect 24168 10821 24202 10845
rect 23145 10724 23171 10758
rect 23171 10724 23179 10758
rect 23217 10724 23239 10758
rect 23239 10724 23251 10758
rect 23289 10724 23307 10758
rect 23307 10724 23323 10758
rect 23361 10724 23375 10758
rect 23375 10724 23395 10758
rect 23433 10724 23443 10758
rect 23443 10724 23467 10758
rect 23505 10724 23511 10758
rect 23511 10724 23539 10758
rect 23577 10724 23579 10758
rect 23579 10724 23611 10758
rect 23649 10724 23681 10758
rect 23681 10724 23683 10758
rect 23721 10724 23749 10758
rect 23749 10724 23755 10758
rect 23793 10724 23817 10758
rect 23817 10724 23827 10758
rect 23865 10724 23885 10758
rect 23885 10724 23899 10758
rect 23937 10724 23953 10758
rect 23953 10724 23971 10758
rect 24009 10724 24021 10758
rect 24021 10724 24043 10758
rect 24081 10724 24089 10758
rect 24089 10724 24115 10758
rect 24688 12171 24722 12195
rect 24688 12161 24722 12171
rect 24688 12103 24722 12123
rect 24688 12089 24722 12103
rect 24688 12035 24722 12051
rect 24688 12017 24722 12035
rect 24688 11967 24722 11979
rect 24688 11945 24722 11967
rect 24688 11899 24722 11907
rect 24688 11873 24722 11899
rect 24688 11831 24722 11835
rect 24688 11801 24722 11831
rect 24688 11729 24722 11763
rect 24688 11661 24722 11691
rect 24688 11657 24722 11661
rect 24688 11593 24722 11619
rect 24688 11585 24722 11593
rect 24688 11525 24722 11547
rect 24688 11513 24722 11525
rect 24688 11457 24722 11475
rect 24688 11441 24722 11457
rect 24688 11389 24722 11403
rect 24688 11369 24722 11389
rect 24688 11321 24722 11331
rect 24688 11297 24722 11321
rect 25816 12171 25850 12195
rect 25816 12161 25850 12171
rect 25816 12103 25850 12123
rect 25816 12089 25850 12103
rect 25816 12035 25850 12051
rect 25816 12017 25850 12035
rect 25816 11967 25850 11979
rect 25816 11945 25850 11967
rect 25816 11899 25850 11907
rect 25816 11873 25850 11899
rect 25816 11831 25850 11835
rect 25816 11801 25850 11831
rect 25816 11729 25850 11763
rect 25816 11661 25850 11691
rect 25816 11657 25850 11661
rect 25816 11593 25850 11619
rect 25816 11585 25850 11593
rect 25816 11525 25850 11547
rect 25816 11513 25850 11525
rect 25816 11457 25850 11475
rect 25816 11441 25850 11457
rect 25816 11389 25850 11403
rect 25816 11369 25850 11389
rect 25816 11321 25850 11331
rect 25816 11297 25850 11321
rect 24784 11200 24810 11234
rect 24810 11200 24818 11234
rect 24856 11200 24878 11234
rect 24878 11200 24890 11234
rect 24928 11200 24946 11234
rect 24946 11200 24962 11234
rect 25000 11200 25014 11234
rect 25014 11200 25034 11234
rect 25072 11200 25082 11234
rect 25082 11200 25106 11234
rect 25144 11200 25150 11234
rect 25150 11200 25178 11234
rect 25216 11200 25218 11234
rect 25218 11200 25250 11234
rect 25288 11200 25320 11234
rect 25320 11200 25322 11234
rect 25360 11200 25388 11234
rect 25388 11200 25394 11234
rect 25432 11200 25456 11234
rect 25456 11200 25466 11234
rect 25504 11200 25524 11234
rect 25524 11200 25538 11234
rect 25576 11200 25592 11234
rect 25592 11200 25610 11234
rect 25648 11200 25660 11234
rect 25660 11200 25682 11234
rect 25720 11200 25728 11234
rect 25728 11200 25754 11234
rect 24688 11113 24722 11137
rect 24688 11103 24722 11113
rect 24688 11045 24722 11065
rect 24688 11031 24722 11045
rect 24688 10977 24722 10993
rect 24688 10959 24722 10977
rect 24688 10909 24722 10921
rect 24688 10887 24722 10909
rect 24688 10841 24722 10849
rect 24688 10815 24722 10841
rect 24688 10773 24722 10777
rect 24688 10743 24722 10773
rect 24688 10671 24722 10705
rect 24688 10603 24722 10633
rect 24688 10599 24722 10603
rect 24688 10535 24722 10561
rect 24688 10527 24722 10535
rect 24688 10467 24722 10489
rect 24688 10455 24722 10467
rect 24688 10399 24722 10417
rect 24688 10383 24722 10399
rect 24688 10331 24722 10345
rect 24688 10311 24722 10331
rect 24688 10263 24722 10273
rect 24688 10239 24722 10263
rect 25816 11113 25850 11137
rect 25816 11103 25850 11113
rect 25816 11045 25850 11065
rect 25816 11031 25850 11045
rect 25816 10977 25850 10993
rect 25816 10959 25850 10977
rect 25816 10909 25850 10921
rect 25816 10887 25850 10909
rect 25816 10841 25850 10849
rect 25816 10815 25850 10841
rect 25816 10773 25850 10777
rect 25816 10743 25850 10773
rect 25816 10671 25850 10705
rect 25816 10603 25850 10633
rect 25816 10599 25850 10603
rect 25816 10535 25850 10561
rect 25816 10527 25850 10535
rect 25816 10467 25850 10489
rect 25816 10455 25850 10467
rect 25816 10399 25850 10417
rect 25816 10383 25850 10399
rect 25816 10331 25850 10345
rect 25816 10311 25850 10331
rect 25816 10263 25850 10273
rect 25816 10239 25850 10263
rect 24784 10142 24810 10176
rect 24810 10142 24818 10176
rect 24856 10142 24878 10176
rect 24878 10142 24890 10176
rect 24928 10142 24946 10176
rect 24946 10142 24962 10176
rect 25000 10142 25014 10176
rect 25014 10142 25034 10176
rect 25072 10142 25082 10176
rect 25082 10142 25106 10176
rect 25144 10142 25150 10176
rect 25150 10142 25178 10176
rect 25216 10142 25218 10176
rect 25218 10142 25250 10176
rect 25288 10142 25320 10176
rect 25320 10142 25322 10176
rect 25360 10142 25388 10176
rect 25388 10142 25394 10176
rect 25432 10142 25456 10176
rect 25456 10142 25466 10176
rect 25504 10142 25524 10176
rect 25524 10142 25538 10176
rect 25576 10142 25592 10176
rect 25592 10142 25610 10176
rect 25648 10142 25660 10176
rect 25660 10142 25682 10176
rect 25720 10142 25728 10176
rect 25728 10142 25754 10176
rect 24688 10055 24722 10079
rect 24688 10045 24722 10055
rect 24688 9987 24722 10007
rect 24688 9973 24722 9987
rect 24688 9919 24722 9935
rect 24688 9901 24722 9919
rect 24688 9851 24722 9863
rect 24688 9829 24722 9851
rect 24688 9783 24722 9791
rect 24688 9757 24722 9783
rect 24688 9715 24722 9719
rect 24688 9685 24722 9715
rect 24688 9613 24722 9647
rect 24688 9545 24722 9575
rect 24688 9541 24722 9545
rect 24688 9477 24722 9503
rect 24688 9469 24722 9477
rect 24688 9409 24722 9431
rect 24688 9397 24722 9409
rect 24688 9341 24722 9359
rect 24688 9325 24722 9341
rect 24688 9273 24722 9287
rect 24688 9253 24722 9273
rect 24688 9205 24722 9215
rect 24688 9181 24722 9205
rect 25816 10055 25850 10079
rect 25816 10045 25850 10055
rect 25816 9987 25850 10007
rect 25816 9973 25850 9987
rect 25816 9919 25850 9935
rect 25816 9901 25850 9919
rect 25816 9851 25850 9863
rect 25816 9829 25850 9851
rect 25816 9783 25850 9791
rect 25816 9757 25850 9783
rect 25816 9715 25850 9719
rect 25816 9685 25850 9715
rect 25816 9613 25850 9647
rect 25816 9545 25850 9575
rect 25816 9541 25850 9545
rect 25816 9477 25850 9503
rect 25816 9469 25850 9477
rect 25816 9409 25850 9431
rect 25816 9397 25850 9409
rect 25816 9341 25850 9359
rect 25816 9325 25850 9341
rect 25816 9273 25850 9287
rect 25816 9253 25850 9273
rect 25816 9205 25850 9215
rect 25816 9181 25850 9205
rect 24784 9084 24810 9118
rect 24810 9084 24818 9118
rect 24856 9084 24878 9118
rect 24878 9084 24890 9118
rect 24928 9084 24946 9118
rect 24946 9084 24962 9118
rect 25000 9084 25014 9118
rect 25014 9084 25034 9118
rect 25072 9084 25082 9118
rect 25082 9084 25106 9118
rect 25144 9084 25150 9118
rect 25150 9084 25178 9118
rect 25216 9084 25218 9118
rect 25218 9084 25250 9118
rect 25288 9084 25320 9118
rect 25320 9084 25322 9118
rect 25360 9084 25388 9118
rect 25388 9084 25394 9118
rect 25432 9084 25456 9118
rect 25456 9084 25466 9118
rect 25504 9084 25524 9118
rect 25524 9084 25538 9118
rect 25576 9084 25592 9118
rect 25592 9084 25610 9118
rect 25648 9084 25660 9118
rect 25660 9084 25682 9118
rect 25720 9084 25728 9118
rect 25728 9084 25754 9118
rect 21898 7093 22436 7631
rect 23625 7846 23651 7880
rect 23651 7846 23659 7880
rect 23697 7846 23719 7880
rect 23719 7846 23731 7880
rect 23769 7846 23787 7880
rect 23787 7846 23803 7880
rect 23841 7846 23855 7880
rect 23855 7846 23875 7880
rect 23913 7846 23923 7880
rect 23923 7846 23947 7880
rect 23985 7846 23991 7880
rect 23991 7846 24019 7880
rect 24057 7846 24059 7880
rect 24059 7846 24091 7880
rect 24129 7846 24161 7880
rect 24161 7846 24163 7880
rect 24201 7846 24229 7880
rect 24229 7846 24235 7880
rect 24273 7846 24297 7880
rect 24297 7846 24307 7880
rect 24345 7846 24365 7880
rect 24365 7846 24379 7880
rect 24417 7846 24433 7880
rect 24433 7846 24451 7880
rect 24489 7846 24501 7880
rect 24501 7846 24523 7880
rect 24561 7846 24569 7880
rect 24569 7846 24595 7880
rect 20530 5099 20564 5133
rect 20530 5027 20564 5061
rect 20530 4955 20564 4989
rect 20530 4883 20564 4917
rect 20530 4811 20564 4845
rect 20530 4739 20564 4773
rect 20848 5099 20882 5133
rect 20848 5027 20882 5061
rect 20848 4955 20882 4989
rect 20848 4883 20882 4917
rect 20848 4811 20882 4845
rect 20848 4739 20882 4773
rect 21166 5099 21200 5133
rect 21166 5027 21200 5061
rect 21166 4955 21200 4989
rect 21166 4883 21200 4917
rect 21166 4811 21200 4845
rect 21166 4739 21200 4773
rect 21484 5099 21518 5133
rect 23538 7759 23572 7783
rect 23538 7749 23572 7759
rect 23538 7691 23572 7711
rect 23538 7677 23572 7691
rect 23538 7623 23572 7639
rect 23538 7605 23572 7623
rect 23538 7555 23572 7567
rect 23538 7533 23572 7555
rect 23538 7487 23572 7495
rect 23538 7461 23572 7487
rect 23538 7419 23572 7423
rect 23538 7389 23572 7419
rect 23538 7317 23572 7351
rect 23538 7249 23572 7279
rect 23538 7245 23572 7249
rect 23538 7181 23572 7207
rect 23538 7173 23572 7181
rect 23538 7113 23572 7135
rect 23538 7101 23572 7113
rect 23538 7045 23572 7063
rect 23538 7029 23572 7045
rect 23538 6977 23572 6991
rect 23538 6957 23572 6977
rect 23538 6909 23572 6919
rect 23538 6885 23572 6909
rect 24648 7759 24682 7783
rect 24648 7749 24682 7759
rect 24648 7691 24682 7711
rect 24648 7677 24682 7691
rect 24648 7623 24682 7639
rect 24648 7605 24682 7623
rect 24648 7555 24682 7567
rect 24648 7533 24682 7555
rect 24648 7487 24682 7495
rect 24648 7461 24682 7487
rect 24648 7419 24682 7423
rect 24648 7389 24682 7419
rect 24648 7317 24682 7351
rect 24648 7249 24682 7279
rect 24648 7245 24682 7249
rect 24648 7181 24682 7207
rect 24648 7173 24682 7181
rect 24648 7113 24682 7135
rect 24648 7101 24682 7113
rect 24648 7045 24682 7063
rect 24648 7029 24682 7045
rect 24648 6977 24682 6991
rect 24648 6957 24682 6977
rect 24648 6909 24682 6919
rect 24648 6885 24682 6909
rect 23625 6788 23651 6822
rect 23651 6788 23659 6822
rect 23697 6788 23719 6822
rect 23719 6788 23731 6822
rect 23769 6788 23787 6822
rect 23787 6788 23803 6822
rect 23841 6788 23855 6822
rect 23855 6788 23875 6822
rect 23913 6788 23923 6822
rect 23923 6788 23947 6822
rect 23985 6788 23991 6822
rect 23991 6788 24019 6822
rect 24057 6788 24059 6822
rect 24059 6788 24091 6822
rect 24129 6788 24161 6822
rect 24161 6788 24163 6822
rect 24201 6788 24229 6822
rect 24229 6788 24235 6822
rect 24273 6788 24297 6822
rect 24297 6788 24307 6822
rect 24345 6788 24365 6822
rect 24365 6788 24379 6822
rect 24417 6788 24433 6822
rect 24433 6788 24451 6822
rect 24489 6788 24501 6822
rect 24501 6788 24523 6822
rect 24561 6788 24569 6822
rect 24569 6788 24595 6822
rect 23538 6701 23572 6725
rect 23538 6691 23572 6701
rect 23538 6633 23572 6653
rect 23538 6619 23572 6633
rect 23538 6565 23572 6581
rect 23538 6547 23572 6565
rect 23538 6497 23572 6509
rect 23538 6475 23572 6497
rect 23538 6429 23572 6437
rect 23538 6403 23572 6429
rect 23538 6361 23572 6365
rect 23538 6331 23572 6361
rect 23538 6259 23572 6293
rect 23538 6191 23572 6221
rect 23538 6187 23572 6191
rect 23538 6123 23572 6149
rect 23538 6115 23572 6123
rect 23538 6055 23572 6077
rect 23538 6043 23572 6055
rect 23538 5987 23572 6005
rect 23538 5971 23572 5987
rect 23538 5919 23572 5933
rect 23538 5899 23572 5919
rect 23538 5851 23572 5861
rect 23538 5827 23572 5851
rect 24648 6701 24682 6725
rect 24648 6691 24682 6701
rect 24648 6633 24682 6653
rect 24648 6619 24682 6633
rect 24648 6565 24682 6581
rect 24648 6547 24682 6565
rect 24648 6497 24682 6509
rect 24648 6475 24682 6497
rect 24648 6429 24682 6437
rect 24648 6403 24682 6429
rect 24648 6361 24682 6365
rect 24648 6331 24682 6361
rect 24648 6259 24682 6293
rect 24648 6191 24682 6221
rect 24648 6187 24682 6191
rect 24648 6123 24682 6149
rect 24648 6115 24682 6123
rect 24648 6055 24682 6077
rect 24648 6043 24682 6055
rect 24648 5987 24682 6005
rect 24648 5971 24682 5987
rect 24648 5919 24682 5933
rect 24648 5899 24682 5919
rect 24648 5851 24682 5861
rect 24648 5827 24682 5851
rect 23625 5730 23651 5764
rect 23651 5730 23659 5764
rect 23697 5730 23719 5764
rect 23719 5730 23731 5764
rect 23769 5730 23787 5764
rect 23787 5730 23803 5764
rect 23841 5730 23855 5764
rect 23855 5730 23875 5764
rect 23913 5730 23923 5764
rect 23923 5730 23947 5764
rect 23985 5730 23991 5764
rect 23991 5730 24019 5764
rect 24057 5730 24059 5764
rect 24059 5730 24091 5764
rect 24129 5730 24161 5764
rect 24161 5730 24163 5764
rect 24201 5730 24229 5764
rect 24229 5730 24235 5764
rect 24273 5730 24297 5764
rect 24297 5730 24307 5764
rect 24345 5730 24365 5764
rect 24365 5730 24379 5764
rect 24417 5730 24433 5764
rect 24433 5730 24451 5764
rect 24489 5730 24501 5764
rect 24501 5730 24523 5764
rect 24561 5730 24569 5764
rect 24569 5730 24595 5764
rect 21484 5027 21518 5061
rect 21484 4955 21518 4989
rect 21484 4883 21518 4917
rect 21484 4811 21518 4845
rect 21484 4739 21518 4773
rect 23538 5643 23572 5667
rect 23538 5633 23572 5643
rect 23538 5575 23572 5595
rect 23538 5561 23572 5575
rect 23538 5507 23572 5523
rect 23538 5489 23572 5507
rect 23538 5439 23572 5451
rect 23538 5417 23572 5439
rect 23538 5371 23572 5379
rect 23538 5345 23572 5371
rect 23538 5303 23572 5307
rect 23538 5273 23572 5303
rect 23538 5201 23572 5235
rect 23538 5133 23572 5163
rect 23538 5129 23572 5133
rect 23538 5065 23572 5091
rect 23538 5057 23572 5065
rect 23538 4997 23572 5019
rect 23538 4985 23572 4997
rect 23538 4929 23572 4947
rect 23538 4913 23572 4929
rect 23538 4861 23572 4875
rect 23538 4841 23572 4861
rect 23538 4793 23572 4803
rect 23538 4769 23572 4793
rect 24648 5643 24682 5667
rect 24648 5633 24682 5643
rect 24648 5575 24682 5595
rect 24648 5561 24682 5575
rect 24648 5507 24682 5523
rect 24648 5489 24682 5507
rect 24648 5439 24682 5451
rect 24648 5417 24682 5439
rect 24648 5371 24682 5379
rect 24648 5345 24682 5371
rect 24648 5303 24682 5307
rect 24648 5273 24682 5303
rect 24648 5201 24682 5235
rect 24648 5133 24682 5163
rect 24648 5129 24682 5133
rect 24648 5065 24682 5091
rect 24648 5057 24682 5065
rect 24648 4997 24682 5019
rect 24648 4985 24682 4997
rect 24648 4929 24682 4947
rect 24648 4913 24682 4929
rect 24648 4861 24682 4875
rect 24648 4841 24682 4861
rect 24648 4793 24682 4803
rect 24648 4769 24682 4793
rect 23625 4672 23651 4706
rect 23651 4672 23659 4706
rect 23697 4672 23719 4706
rect 23719 4672 23731 4706
rect 23769 4672 23787 4706
rect 23787 4672 23803 4706
rect 23841 4672 23855 4706
rect 23855 4672 23875 4706
rect 23913 4672 23923 4706
rect 23923 4672 23947 4706
rect 23985 4672 23991 4706
rect 23991 4672 24019 4706
rect 24057 4672 24059 4706
rect 24059 4672 24091 4706
rect 24129 4672 24161 4706
rect 24161 4672 24163 4706
rect 24201 4672 24229 4706
rect 24229 4672 24235 4706
rect 24273 4672 24297 4706
rect 24297 4672 24307 4706
rect 24345 4672 24365 4706
rect 24365 4672 24379 4706
rect 24417 4672 24433 4706
rect 24433 4672 24451 4706
rect 24489 4672 24501 4706
rect 24501 4672 24523 4706
rect 24561 4672 24569 4706
rect 24569 4672 24595 4706
rect 18981 4476 19005 4510
rect 19005 4476 19015 4510
rect 19053 4476 19073 4510
rect 19073 4476 19087 4510
rect 19125 4476 19141 4510
rect 19141 4476 19159 4510
rect 19197 4476 19209 4510
rect 19209 4476 19231 4510
rect 19269 4476 19277 4510
rect 19277 4476 19303 4510
rect 19341 4476 19345 4510
rect 19345 4476 19375 4510
rect 19413 4476 19447 4510
rect 19485 4476 19515 4510
rect 19515 4476 19519 4510
rect 19557 4476 19583 4510
rect 19583 4476 19591 4510
rect 19629 4476 19651 4510
rect 19651 4476 19663 4510
rect 19701 4476 19719 4510
rect 19719 4476 19735 4510
rect 19773 4476 19787 4510
rect 19787 4476 19807 4510
rect 19845 4476 19855 4510
rect 19855 4476 19879 4510
rect 12824 3815 22650 4209
rect 23538 4585 23572 4609
rect 23538 4575 23572 4585
rect 23538 4517 23572 4537
rect 23538 4503 23572 4517
rect 23538 4449 23572 4465
rect 23538 4431 23572 4449
rect 23538 4381 23572 4393
rect 23538 4359 23572 4381
rect 23538 4313 23572 4321
rect 23538 4287 23572 4313
rect 23538 4245 23572 4249
rect 23538 4215 23572 4245
rect 23538 4143 23572 4177
rect 23538 4075 23572 4105
rect 23538 4071 23572 4075
rect 23538 4007 23572 4033
rect 23538 3999 23572 4007
rect 23538 3939 23572 3961
rect 23538 3927 23572 3939
rect 23538 3871 23572 3889
rect 23538 3855 23572 3871
rect 23538 3803 23572 3817
rect 23538 3783 23572 3803
rect 23538 3735 23572 3745
rect 23538 3711 23572 3735
rect 24648 4585 24682 4609
rect 24648 4575 24682 4585
rect 24648 4517 24682 4537
rect 24648 4503 24682 4517
rect 24648 4449 24682 4465
rect 24648 4431 24682 4449
rect 24648 4381 24682 4393
rect 24648 4359 24682 4381
rect 24648 4313 24682 4321
rect 24648 4287 24682 4313
rect 24648 4245 24682 4249
rect 24648 4215 24682 4245
rect 24648 4143 24682 4177
rect 24648 4075 24682 4105
rect 24648 4071 24682 4075
rect 24648 4007 24682 4033
rect 24648 3999 24682 4007
rect 24648 3939 24682 3961
rect 24648 3927 24682 3939
rect 24648 3871 24682 3889
rect 24648 3855 24682 3871
rect 24648 3803 24682 3817
rect 24648 3783 24682 3803
rect 24648 3735 24682 3745
rect 24648 3711 24682 3735
rect 23625 3614 23651 3648
rect 23651 3614 23659 3648
rect 23697 3614 23719 3648
rect 23719 3614 23731 3648
rect 23769 3614 23787 3648
rect 23787 3614 23803 3648
rect 23841 3614 23855 3648
rect 23855 3614 23875 3648
rect 23913 3614 23923 3648
rect 23923 3614 23947 3648
rect 23985 3614 23991 3648
rect 23991 3614 24019 3648
rect 24057 3614 24059 3648
rect 24059 3614 24091 3648
rect 24129 3614 24161 3648
rect 24161 3614 24163 3648
rect 24201 3614 24229 3648
rect 24229 3614 24235 3648
rect 24273 3614 24297 3648
rect 24297 3614 24307 3648
rect 24345 3614 24365 3648
rect 24365 3614 24379 3648
rect 24417 3614 24433 3648
rect 24433 3614 24451 3648
rect 24489 3614 24501 3648
rect 24501 3614 24523 3648
rect 24561 3614 24569 3648
rect 24569 3614 24595 3648
rect 25125 7846 25151 7880
rect 25151 7846 25159 7880
rect 25197 7846 25219 7880
rect 25219 7846 25231 7880
rect 25269 7846 25287 7880
rect 25287 7846 25303 7880
rect 25341 7846 25355 7880
rect 25355 7846 25375 7880
rect 25413 7846 25423 7880
rect 25423 7846 25447 7880
rect 25485 7846 25491 7880
rect 25491 7846 25519 7880
rect 25557 7846 25559 7880
rect 25559 7846 25591 7880
rect 25629 7846 25661 7880
rect 25661 7846 25663 7880
rect 25701 7846 25729 7880
rect 25729 7846 25735 7880
rect 25773 7846 25797 7880
rect 25797 7846 25807 7880
rect 25845 7846 25865 7880
rect 25865 7846 25879 7880
rect 25917 7846 25933 7880
rect 25933 7846 25951 7880
rect 25989 7846 26001 7880
rect 26001 7846 26023 7880
rect 26061 7846 26069 7880
rect 26069 7846 26095 7880
rect 25038 7759 25072 7783
rect 25038 7749 25072 7759
rect 25038 7691 25072 7711
rect 25038 7677 25072 7691
rect 25038 7623 25072 7639
rect 25038 7605 25072 7623
rect 25038 7555 25072 7567
rect 25038 7533 25072 7555
rect 25038 7487 25072 7495
rect 25038 7461 25072 7487
rect 25038 7419 25072 7423
rect 25038 7389 25072 7419
rect 25038 7317 25072 7351
rect 25038 7249 25072 7279
rect 25038 7245 25072 7249
rect 25038 7181 25072 7207
rect 25038 7173 25072 7181
rect 25038 7113 25072 7135
rect 25038 7101 25072 7113
rect 25038 7045 25072 7063
rect 25038 7029 25072 7045
rect 25038 6977 25072 6991
rect 25038 6957 25072 6977
rect 25038 6909 25072 6919
rect 25038 6885 25072 6909
rect 26148 7759 26182 7783
rect 26148 7749 26182 7759
rect 26148 7691 26182 7711
rect 26148 7677 26182 7691
rect 26148 7623 26182 7639
rect 26148 7605 26182 7623
rect 26148 7555 26182 7567
rect 26148 7533 26182 7555
rect 26148 7487 26182 7495
rect 26148 7461 26182 7487
rect 26148 7419 26182 7423
rect 26148 7389 26182 7419
rect 26148 7317 26182 7351
rect 26148 7249 26182 7279
rect 26148 7245 26182 7249
rect 26148 7181 26182 7207
rect 26148 7173 26182 7181
rect 26148 7113 26182 7135
rect 26148 7101 26182 7113
rect 26148 7045 26182 7063
rect 26148 7029 26182 7045
rect 26148 6977 26182 6991
rect 26148 6957 26182 6977
rect 26148 6909 26182 6919
rect 26148 6885 26182 6909
rect 25125 6788 25151 6822
rect 25151 6788 25159 6822
rect 25197 6788 25219 6822
rect 25219 6788 25231 6822
rect 25269 6788 25287 6822
rect 25287 6788 25303 6822
rect 25341 6788 25355 6822
rect 25355 6788 25375 6822
rect 25413 6788 25423 6822
rect 25423 6788 25447 6822
rect 25485 6788 25491 6822
rect 25491 6788 25519 6822
rect 25557 6788 25559 6822
rect 25559 6788 25591 6822
rect 25629 6788 25661 6822
rect 25661 6788 25663 6822
rect 25701 6788 25729 6822
rect 25729 6788 25735 6822
rect 25773 6788 25797 6822
rect 25797 6788 25807 6822
rect 25845 6788 25865 6822
rect 25865 6788 25879 6822
rect 25917 6788 25933 6822
rect 25933 6788 25951 6822
rect 25989 6788 26001 6822
rect 26001 6788 26023 6822
rect 26061 6788 26069 6822
rect 26069 6788 26095 6822
rect 25038 6701 25072 6725
rect 25038 6691 25072 6701
rect 25038 6633 25072 6653
rect 25038 6619 25072 6633
rect 25038 6565 25072 6581
rect 25038 6547 25072 6565
rect 25038 6497 25072 6509
rect 25038 6475 25072 6497
rect 25038 6429 25072 6437
rect 25038 6403 25072 6429
rect 25038 6361 25072 6365
rect 25038 6331 25072 6361
rect 25038 6259 25072 6293
rect 25038 6191 25072 6221
rect 25038 6187 25072 6191
rect 25038 6123 25072 6149
rect 25038 6115 25072 6123
rect 25038 6055 25072 6077
rect 25038 6043 25072 6055
rect 25038 5987 25072 6005
rect 25038 5971 25072 5987
rect 25038 5919 25072 5933
rect 25038 5899 25072 5919
rect 25038 5851 25072 5861
rect 25038 5827 25072 5851
rect 26148 6701 26182 6725
rect 26148 6691 26182 6701
rect 26148 6633 26182 6653
rect 26148 6619 26182 6633
rect 26148 6565 26182 6581
rect 26148 6547 26182 6565
rect 26148 6497 26182 6509
rect 26148 6475 26182 6497
rect 26148 6429 26182 6437
rect 26148 6403 26182 6429
rect 26148 6361 26182 6365
rect 26148 6331 26182 6361
rect 26148 6259 26182 6293
rect 26148 6191 26182 6221
rect 26148 6187 26182 6191
rect 26148 6123 26182 6149
rect 26148 6115 26182 6123
rect 26148 6055 26182 6077
rect 26148 6043 26182 6055
rect 26148 5987 26182 6005
rect 26148 5971 26182 5987
rect 26148 5919 26182 5933
rect 26148 5899 26182 5919
rect 26148 5851 26182 5861
rect 26148 5827 26182 5851
rect 25125 5730 25151 5764
rect 25151 5730 25159 5764
rect 25197 5730 25219 5764
rect 25219 5730 25231 5764
rect 25269 5730 25287 5764
rect 25287 5730 25303 5764
rect 25341 5730 25355 5764
rect 25355 5730 25375 5764
rect 25413 5730 25423 5764
rect 25423 5730 25447 5764
rect 25485 5730 25491 5764
rect 25491 5730 25519 5764
rect 25557 5730 25559 5764
rect 25559 5730 25591 5764
rect 25629 5730 25661 5764
rect 25661 5730 25663 5764
rect 25701 5730 25729 5764
rect 25729 5730 25735 5764
rect 25773 5730 25797 5764
rect 25797 5730 25807 5764
rect 25845 5730 25865 5764
rect 25865 5730 25879 5764
rect 25917 5730 25933 5764
rect 25933 5730 25951 5764
rect 25989 5730 26001 5764
rect 26001 5730 26023 5764
rect 26061 5730 26069 5764
rect 26069 5730 26095 5764
rect 25038 5643 25072 5667
rect 25038 5633 25072 5643
rect 25038 5575 25072 5595
rect 25038 5561 25072 5575
rect 25038 5507 25072 5523
rect 25038 5489 25072 5507
rect 25038 5439 25072 5451
rect 25038 5417 25072 5439
rect 25038 5371 25072 5379
rect 25038 5345 25072 5371
rect 25038 5303 25072 5307
rect 25038 5273 25072 5303
rect 25038 5201 25072 5235
rect 25038 5133 25072 5163
rect 25038 5129 25072 5133
rect 25038 5065 25072 5091
rect 25038 5057 25072 5065
rect 25038 4997 25072 5019
rect 25038 4985 25072 4997
rect 25038 4929 25072 4947
rect 25038 4913 25072 4929
rect 25038 4861 25072 4875
rect 25038 4841 25072 4861
rect 25038 4793 25072 4803
rect 25038 4769 25072 4793
rect 26148 5643 26182 5667
rect 26148 5633 26182 5643
rect 26148 5575 26182 5595
rect 26148 5561 26182 5575
rect 26148 5507 26182 5523
rect 26148 5489 26182 5507
rect 26148 5439 26182 5451
rect 26148 5417 26182 5439
rect 26148 5371 26182 5379
rect 26148 5345 26182 5371
rect 26148 5303 26182 5307
rect 26148 5273 26182 5303
rect 26148 5201 26182 5235
rect 26148 5133 26182 5163
rect 26148 5129 26182 5133
rect 26148 5065 26182 5091
rect 26148 5057 26182 5065
rect 26148 4997 26182 5019
rect 26148 4985 26182 4997
rect 26148 4929 26182 4947
rect 26148 4913 26182 4929
rect 26148 4861 26182 4875
rect 26148 4841 26182 4861
rect 26148 4793 26182 4803
rect 26148 4769 26182 4793
rect 25125 4672 25151 4706
rect 25151 4672 25159 4706
rect 25197 4672 25219 4706
rect 25219 4672 25231 4706
rect 25269 4672 25287 4706
rect 25287 4672 25303 4706
rect 25341 4672 25355 4706
rect 25355 4672 25375 4706
rect 25413 4672 25423 4706
rect 25423 4672 25447 4706
rect 25485 4672 25491 4706
rect 25491 4672 25519 4706
rect 25557 4672 25559 4706
rect 25559 4672 25591 4706
rect 25629 4672 25661 4706
rect 25661 4672 25663 4706
rect 25701 4672 25729 4706
rect 25729 4672 25735 4706
rect 25773 4672 25797 4706
rect 25797 4672 25807 4706
rect 25845 4672 25865 4706
rect 25865 4672 25879 4706
rect 25917 4672 25933 4706
rect 25933 4672 25951 4706
rect 25989 4672 26001 4706
rect 26001 4672 26023 4706
rect 26061 4672 26069 4706
rect 26069 4672 26095 4706
rect 25038 4585 25072 4609
rect 25038 4575 25072 4585
rect 25038 4517 25072 4537
rect 25038 4503 25072 4517
rect 25038 4449 25072 4465
rect 25038 4431 25072 4449
rect 25038 4381 25072 4393
rect 25038 4359 25072 4381
rect 25038 4313 25072 4321
rect 25038 4287 25072 4313
rect 25038 4245 25072 4249
rect 25038 4215 25072 4245
rect 25038 4143 25072 4177
rect 25038 4075 25072 4105
rect 25038 4071 25072 4075
rect 25038 4007 25072 4033
rect 25038 3999 25072 4007
rect 25038 3939 25072 3961
rect 25038 3927 25072 3939
rect 25038 3871 25072 3889
rect 25038 3855 25072 3871
rect 25038 3803 25072 3817
rect 25038 3783 25072 3803
rect 25038 3735 25072 3745
rect 25038 3711 25072 3735
rect 26148 4585 26182 4609
rect 26148 4575 26182 4585
rect 26148 4517 26182 4537
rect 26148 4503 26182 4517
rect 26148 4449 26182 4465
rect 26148 4431 26182 4449
rect 26148 4381 26182 4393
rect 26148 4359 26182 4381
rect 26148 4313 26182 4321
rect 26148 4287 26182 4313
rect 26148 4245 26182 4249
rect 26148 4215 26182 4245
rect 26148 4143 26182 4177
rect 26148 4075 26182 4105
rect 26148 4071 26182 4075
rect 26148 4007 26182 4033
rect 26148 3999 26182 4007
rect 26148 3939 26182 3961
rect 26148 3927 26182 3939
rect 26148 3871 26182 3889
rect 26148 3855 26182 3871
rect 26148 3803 26182 3817
rect 26148 3783 26182 3803
rect 26148 3735 26182 3745
rect 26148 3711 26182 3735
rect 25125 3614 25151 3648
rect 25151 3614 25159 3648
rect 25197 3614 25219 3648
rect 25219 3614 25231 3648
rect 25269 3614 25287 3648
rect 25287 3614 25303 3648
rect 25341 3614 25355 3648
rect 25355 3614 25375 3648
rect 25413 3614 25423 3648
rect 25423 3614 25447 3648
rect 25485 3614 25491 3648
rect 25491 3614 25519 3648
rect 25557 3614 25559 3648
rect 25559 3614 25591 3648
rect 25629 3614 25661 3648
rect 25661 3614 25663 3648
rect 25701 3614 25729 3648
rect 25729 3614 25735 3648
rect 25773 3614 25797 3648
rect 25797 3614 25807 3648
rect 25845 3614 25865 3648
rect 25865 3614 25879 3648
rect 25917 3614 25933 3648
rect 25933 3614 25951 3648
rect 25989 3614 26001 3648
rect 26001 3614 26023 3648
rect 26061 3614 26069 3648
rect 26069 3614 26095 3648
rect 28036 13274 28070 13308
rect 28036 13202 28070 13236
rect 28036 13130 28070 13164
rect 28036 13058 28070 13092
rect 28036 12986 28070 13020
rect 28036 12914 28070 12948
rect 28354 13274 28388 13308
rect 28354 13202 28388 13236
rect 28354 13130 28388 13164
rect 28354 13058 28388 13092
rect 28354 12986 28388 13020
rect 28354 12914 28388 12948
rect 28672 13274 28706 13308
rect 28672 13202 28706 13236
rect 28672 13130 28706 13164
rect 28672 13058 28706 13092
rect 28672 12986 28706 13020
rect 28672 12914 28706 12948
rect 28990 13274 29024 13308
rect 28990 13202 29024 13236
rect 28990 13130 29024 13164
rect 28990 13058 29024 13092
rect 28990 12986 29024 13020
rect 28990 12914 29024 12948
rect 29308 13274 29342 13308
rect 29308 13202 29342 13236
rect 29308 13130 29342 13164
rect 29308 13058 29342 13092
rect 29308 12986 29342 13020
rect 29308 12914 29342 12948
rect 38752 13474 38786 13508
rect 38824 13474 38858 13508
rect 39681 15520 39715 15538
rect 39681 15504 39715 15520
rect 39681 15452 39715 15466
rect 39681 15432 39715 15452
rect 39681 15384 39715 15394
rect 39681 15360 39715 15384
rect 39681 15316 39715 15322
rect 39681 15288 39715 15316
rect 39681 15248 39715 15250
rect 39681 15216 39715 15248
rect 39681 15146 39715 15178
rect 39681 15144 39715 15146
rect 39681 15078 39715 15106
rect 39681 15072 39715 15078
rect 39681 15010 39715 15034
rect 39681 15000 39715 15010
rect 39681 14942 39715 14962
rect 39681 14928 39715 14942
rect 39681 14874 39715 14890
rect 39681 14856 39715 14874
rect 39681 14806 39715 14818
rect 39681 14784 39715 14806
rect 39681 14738 39715 14746
rect 39681 14712 39715 14738
rect 39681 14670 39715 14674
rect 39681 14640 39715 14670
rect 39681 14568 39715 14602
rect 39681 14500 39715 14530
rect 39681 14496 39715 14500
rect 39681 14432 39715 14458
rect 39681 14424 39715 14432
rect 39681 14364 39715 14386
rect 39681 14352 39715 14364
rect 39681 14296 39715 14314
rect 39681 14280 39715 14296
rect 39681 14228 39715 14242
rect 39681 14208 39715 14228
rect 39681 14160 39715 14170
rect 39681 14136 39715 14160
rect 39681 14092 39715 14098
rect 39681 14064 39715 14092
rect 39681 14024 39715 14026
rect 39681 13992 39715 14024
rect 39681 13922 39715 13954
rect 39681 13920 39715 13922
rect 39681 13854 39715 13882
rect 39681 13848 39715 13854
rect 39681 13786 39715 13810
rect 39681 13776 39715 13786
rect 39681 13718 39715 13738
rect 39681 13704 39715 13718
rect 39681 13650 39715 13666
rect 39681 13632 39715 13650
rect 40156 15651 40190 15685
rect 40228 15651 40262 15685
rect 40300 15651 40334 15685
rect 39939 15520 39973 15538
rect 39939 15504 39973 15520
rect 39939 15452 39973 15466
rect 39939 15432 39973 15452
rect 39939 15384 39973 15394
rect 39939 15360 39973 15384
rect 39939 15316 39973 15322
rect 39939 15288 39973 15316
rect 39939 15248 39973 15250
rect 39939 15216 39973 15248
rect 39939 15146 39973 15178
rect 39939 15144 39973 15146
rect 39939 15078 39973 15106
rect 39939 15072 39973 15078
rect 39939 15010 39973 15034
rect 39939 15000 39973 15010
rect 39939 14942 39973 14962
rect 39939 14928 39973 14942
rect 39939 14874 39973 14890
rect 39939 14856 39973 14874
rect 39939 14806 39973 14818
rect 39939 14784 39973 14806
rect 39939 14738 39973 14746
rect 39939 14712 39973 14738
rect 39939 14670 39973 14674
rect 39939 14640 39973 14670
rect 39939 14568 39973 14602
rect 39939 14500 39973 14530
rect 39939 14496 39973 14500
rect 39939 14432 39973 14458
rect 39939 14424 39973 14432
rect 39939 14364 39973 14386
rect 39939 14352 39973 14364
rect 39939 14296 39973 14314
rect 39939 14280 39973 14296
rect 39939 14228 39973 14242
rect 39939 14208 39973 14228
rect 39939 14160 39973 14170
rect 39939 14136 39973 14160
rect 39939 14092 39973 14098
rect 39939 14064 39973 14092
rect 39939 14024 39973 14026
rect 39939 13992 39973 14024
rect 39939 13922 39973 13954
rect 39939 13920 39973 13922
rect 39939 13854 39973 13882
rect 39939 13848 39973 13854
rect 39939 13786 39973 13810
rect 39939 13776 39973 13786
rect 39939 13718 39973 13738
rect 39939 13704 39973 13718
rect 39939 13650 39973 13666
rect 39939 13632 39973 13650
rect 40197 15520 40231 15538
rect 40197 15504 40231 15520
rect 40197 15452 40231 15466
rect 40197 15432 40231 15452
rect 40197 15384 40231 15394
rect 40197 15360 40231 15384
rect 40197 15316 40231 15322
rect 40197 15288 40231 15316
rect 40197 15248 40231 15250
rect 40197 15216 40231 15248
rect 40197 15146 40231 15178
rect 40197 15144 40231 15146
rect 40197 15078 40231 15106
rect 40197 15072 40231 15078
rect 40197 15010 40231 15034
rect 40197 15000 40231 15010
rect 40197 14942 40231 14962
rect 40197 14928 40231 14942
rect 40197 14874 40231 14890
rect 40197 14856 40231 14874
rect 40197 14806 40231 14818
rect 40197 14784 40231 14806
rect 40197 14738 40231 14746
rect 40197 14712 40231 14738
rect 40197 14670 40231 14674
rect 40197 14640 40231 14670
rect 40197 14568 40231 14602
rect 40197 14500 40231 14530
rect 40197 14496 40231 14500
rect 40197 14432 40231 14458
rect 40197 14424 40231 14432
rect 40197 14364 40231 14386
rect 40197 14352 40231 14364
rect 40197 14296 40231 14314
rect 40197 14280 40231 14296
rect 40197 14228 40231 14242
rect 40197 14208 40231 14228
rect 40197 14160 40231 14170
rect 40197 14136 40231 14160
rect 40197 14092 40231 14098
rect 40197 14064 40231 14092
rect 40197 14024 40231 14026
rect 40197 13992 40231 14024
rect 40197 13922 40231 13954
rect 40197 13920 40231 13922
rect 40197 13854 40231 13882
rect 40197 13848 40231 13854
rect 40197 13786 40231 13810
rect 40197 13776 40231 13786
rect 40197 13718 40231 13738
rect 40197 13704 40231 13718
rect 40197 13650 40231 13666
rect 40197 13632 40231 13650
rect 40455 15520 40489 15538
rect 40455 15504 40489 15520
rect 40455 15452 40489 15466
rect 40455 15432 40489 15452
rect 40455 15384 40489 15394
rect 40455 15360 40489 15384
rect 40455 15316 40489 15322
rect 40455 15288 40489 15316
rect 40455 15248 40489 15250
rect 40455 15216 40489 15248
rect 40455 15146 40489 15178
rect 40455 15144 40489 15146
rect 40455 15078 40489 15106
rect 40455 15072 40489 15078
rect 40455 15010 40489 15034
rect 40455 15000 40489 15010
rect 40455 14942 40489 14962
rect 40455 14928 40489 14942
rect 40455 14874 40489 14890
rect 40455 14856 40489 14874
rect 40455 14806 40489 14818
rect 40455 14784 40489 14806
rect 40455 14738 40489 14746
rect 40455 14712 40489 14738
rect 40455 14670 40489 14674
rect 40455 14640 40489 14670
rect 40455 14568 40489 14602
rect 40455 14500 40489 14530
rect 40455 14496 40489 14500
rect 40455 14432 40489 14458
rect 40455 14424 40489 14432
rect 40455 14364 40489 14386
rect 40455 14352 40489 14364
rect 40455 14296 40489 14314
rect 40455 14280 40489 14296
rect 40455 14228 40489 14242
rect 40455 14208 40489 14228
rect 40455 14160 40489 14170
rect 40455 14136 40489 14160
rect 40455 14092 40489 14098
rect 40455 14064 40489 14092
rect 40455 14024 40489 14026
rect 40455 13992 40489 14024
rect 40455 13922 40489 13954
rect 40455 13920 40489 13922
rect 40455 13854 40489 13882
rect 40455 13848 40489 13854
rect 40455 13786 40489 13810
rect 40455 13776 40489 13786
rect 40455 13718 40489 13738
rect 40455 13704 40489 13718
rect 40455 13650 40489 13666
rect 40455 13632 40489 13650
rect 40713 15520 40747 15538
rect 40713 15504 40747 15520
rect 40713 15452 40747 15466
rect 40713 15432 40747 15452
rect 40713 15384 40747 15394
rect 40713 15360 40747 15384
rect 40713 15316 40747 15322
rect 40713 15288 40747 15316
rect 40713 15248 40747 15250
rect 40713 15216 40747 15248
rect 40713 15146 40747 15178
rect 40713 15144 40747 15146
rect 40713 15078 40747 15106
rect 40713 15072 40747 15078
rect 40713 15010 40747 15034
rect 40713 15000 40747 15010
rect 40713 14942 40747 14962
rect 40713 14928 40747 14942
rect 40713 14874 40747 14890
rect 40713 14856 40747 14874
rect 40713 14806 40747 14818
rect 40713 14784 40747 14806
rect 40713 14738 40747 14746
rect 40713 14712 40747 14738
rect 40713 14670 40747 14674
rect 40713 14640 40747 14670
rect 40713 14568 40747 14602
rect 40713 14500 40747 14530
rect 40713 14496 40747 14500
rect 40713 14432 40747 14458
rect 40713 14424 40747 14432
rect 40713 14364 40747 14386
rect 40713 14352 40747 14364
rect 40713 14296 40747 14314
rect 40713 14280 40747 14296
rect 40713 14228 40747 14242
rect 40713 14208 40747 14228
rect 40713 14160 40747 14170
rect 40713 14136 40747 14160
rect 40713 14092 40747 14098
rect 40713 14064 40747 14092
rect 40713 14024 40747 14026
rect 40713 13992 40747 14024
rect 40713 13922 40747 13954
rect 40713 13920 40747 13922
rect 40713 13854 40747 13882
rect 40713 13848 40747 13854
rect 40713 13786 40747 13810
rect 40713 13776 40747 13786
rect 40713 13718 40747 13738
rect 40713 13704 40747 13718
rect 40713 13650 40747 13666
rect 40713 13632 40747 13650
rect 29626 13274 29660 13308
rect 29626 13202 29660 13236
rect 29626 13130 29660 13164
rect 29626 13058 29660 13092
rect 29626 12986 29660 13020
rect 38253 13268 38287 13302
rect 38253 13196 38287 13230
rect 39042 13276 39076 13310
rect 39042 13204 39076 13238
rect 39282 13278 39316 13312
rect 39282 13206 39316 13240
rect 40061 13273 40095 13307
rect 40061 13201 40095 13235
rect 40330 13286 40364 13320
rect 40330 13214 40364 13248
rect 41730 15601 41764 15635
rect 41730 15529 41764 15563
rect 41730 15457 41764 15491
rect 41730 15385 41764 15419
rect 41730 15313 41764 15347
rect 41730 15241 41764 15275
rect 41730 13570 41764 13604
rect 41730 13498 41764 13532
rect 41730 13426 41764 13460
rect 41730 13354 41764 13388
rect 41730 13282 41764 13316
rect 41730 13210 41764 13244
rect 29626 12914 29660 12948
rect 36870 11952 36872 11986
rect 36872 11952 36904 11986
rect 36942 11952 36974 11986
rect 36974 11952 36976 11986
rect 37128 11952 37130 11986
rect 37130 11952 37162 11986
rect 37200 11952 37232 11986
rect 37232 11952 37234 11986
rect 37386 11952 37388 11986
rect 37388 11952 37420 11986
rect 37458 11952 37490 11986
rect 37490 11952 37492 11986
rect 37644 11952 37646 11986
rect 37646 11952 37678 11986
rect 37716 11952 37748 11986
rect 37748 11952 37750 11986
rect 37902 11952 37904 11986
rect 37904 11952 37936 11986
rect 37974 11952 38006 11986
rect 38006 11952 38008 11986
rect 38160 11952 38162 11986
rect 38162 11952 38194 11986
rect 38232 11952 38264 11986
rect 38264 11952 38266 11986
rect 38418 11952 38420 11986
rect 38420 11952 38452 11986
rect 38490 11952 38522 11986
rect 38522 11952 38524 11986
rect 38676 11952 38678 11986
rect 38678 11952 38710 11986
rect 38748 11952 38780 11986
rect 38780 11952 38782 11986
rect 38934 11952 38936 11986
rect 38936 11952 38968 11986
rect 39006 11952 39038 11986
rect 39038 11952 39040 11986
rect 39192 11952 39194 11986
rect 39194 11952 39226 11986
rect 39264 11952 39296 11986
rect 39296 11952 39298 11986
rect 39450 11952 39452 11986
rect 39452 11952 39484 11986
rect 39522 11952 39554 11986
rect 39554 11952 39556 11986
rect 39708 11952 39710 11986
rect 39710 11952 39742 11986
rect 39780 11952 39812 11986
rect 39812 11952 39814 11986
rect 39966 11952 39968 11986
rect 39968 11952 40000 11986
rect 40038 11952 40070 11986
rect 40070 11952 40072 11986
rect 40224 11952 40226 11986
rect 40226 11952 40258 11986
rect 40296 11952 40328 11986
rect 40328 11952 40330 11986
rect 40482 11952 40484 11986
rect 40484 11952 40516 11986
rect 40554 11952 40586 11986
rect 40586 11952 40588 11986
rect 40740 11952 40742 11986
rect 40742 11952 40774 11986
rect 40812 11952 40844 11986
rect 40844 11952 40846 11986
rect 40998 11952 41000 11986
rect 41000 11952 41032 11986
rect 41070 11952 41102 11986
rect 41102 11952 41104 11986
rect 41256 11952 41258 11986
rect 41258 11952 41290 11986
rect 41328 11952 41360 11986
rect 41360 11952 41362 11986
rect 41514 11952 41516 11986
rect 41516 11952 41548 11986
rect 41586 11952 41618 11986
rect 41618 11952 41620 11986
rect 41772 11952 41774 11986
rect 41774 11952 41806 11986
rect 41844 11952 41876 11986
rect 41876 11952 41878 11986
rect 36777 11873 36811 11899
rect 36777 11865 36811 11873
rect 36777 11805 36811 11827
rect 36777 11793 36811 11805
rect 36777 11737 36811 11755
rect 36777 11721 36811 11737
rect 36777 11669 36811 11683
rect 36777 11649 36811 11669
rect 36777 11601 36811 11611
rect 36777 11577 36811 11601
rect 36777 11533 36811 11539
rect 36777 11505 36811 11533
rect 36777 11465 36811 11467
rect 36777 11433 36811 11465
rect 36777 11363 36811 11395
rect 36777 11361 36811 11363
rect 36777 11295 36811 11323
rect 36777 11289 36811 11295
rect 36777 11227 36811 11251
rect 36777 11217 36811 11227
rect 36777 11159 36811 11179
rect 36777 11145 36811 11159
rect 36777 11091 36811 11107
rect 36777 11073 36811 11091
rect 36777 11023 36811 11035
rect 36777 11001 36811 11023
rect 36777 10955 36811 10963
rect 36777 10929 36811 10955
rect 37035 11873 37069 11899
rect 37035 11865 37069 11873
rect 37035 11805 37069 11827
rect 37035 11793 37069 11805
rect 37035 11737 37069 11755
rect 37035 11721 37069 11737
rect 37035 11669 37069 11683
rect 37035 11649 37069 11669
rect 37035 11601 37069 11611
rect 37035 11577 37069 11601
rect 37035 11533 37069 11539
rect 37035 11505 37069 11533
rect 37035 11465 37069 11467
rect 37035 11433 37069 11465
rect 37035 11363 37069 11395
rect 37035 11361 37069 11363
rect 37035 11295 37069 11323
rect 37035 11289 37069 11295
rect 37035 11227 37069 11251
rect 37035 11217 37069 11227
rect 37035 11159 37069 11179
rect 37035 11145 37069 11159
rect 37035 11091 37069 11107
rect 37035 11073 37069 11091
rect 37035 11023 37069 11035
rect 37035 11001 37069 11023
rect 37035 10955 37069 10963
rect 37035 10929 37069 10955
rect 37293 11873 37327 11899
rect 37293 11865 37327 11873
rect 37293 11805 37327 11827
rect 37293 11793 37327 11805
rect 37293 11737 37327 11755
rect 37293 11721 37327 11737
rect 37293 11669 37327 11683
rect 37293 11649 37327 11669
rect 37293 11601 37327 11611
rect 37293 11577 37327 11601
rect 37293 11533 37327 11539
rect 37293 11505 37327 11533
rect 37293 11465 37327 11467
rect 37293 11433 37327 11465
rect 37293 11363 37327 11395
rect 37293 11361 37327 11363
rect 37293 11295 37327 11323
rect 37293 11289 37327 11295
rect 37293 11227 37327 11251
rect 37293 11217 37327 11227
rect 37293 11159 37327 11179
rect 37293 11145 37327 11159
rect 37293 11091 37327 11107
rect 37293 11073 37327 11091
rect 37293 11023 37327 11035
rect 37293 11001 37327 11023
rect 37293 10955 37327 10963
rect 37293 10929 37327 10955
rect 37551 11873 37585 11899
rect 37551 11865 37585 11873
rect 37551 11805 37585 11827
rect 37551 11793 37585 11805
rect 37551 11737 37585 11755
rect 37551 11721 37585 11737
rect 37551 11669 37585 11683
rect 37551 11649 37585 11669
rect 37551 11601 37585 11611
rect 37551 11577 37585 11601
rect 37551 11533 37585 11539
rect 37551 11505 37585 11533
rect 37551 11465 37585 11467
rect 37551 11433 37585 11465
rect 37551 11363 37585 11395
rect 37551 11361 37585 11363
rect 37551 11295 37585 11323
rect 37551 11289 37585 11295
rect 37551 11227 37585 11251
rect 37551 11217 37585 11227
rect 37551 11159 37585 11179
rect 37551 11145 37585 11159
rect 37551 11091 37585 11107
rect 37551 11073 37585 11091
rect 37551 11023 37585 11035
rect 37551 11001 37585 11023
rect 37551 10955 37585 10963
rect 37551 10929 37585 10955
rect 37809 11873 37843 11899
rect 37809 11865 37843 11873
rect 37809 11805 37843 11827
rect 37809 11793 37843 11805
rect 37809 11737 37843 11755
rect 37809 11721 37843 11737
rect 37809 11669 37843 11683
rect 37809 11649 37843 11669
rect 37809 11601 37843 11611
rect 37809 11577 37843 11601
rect 37809 11533 37843 11539
rect 37809 11505 37843 11533
rect 37809 11465 37843 11467
rect 37809 11433 37843 11465
rect 37809 11363 37843 11395
rect 37809 11361 37843 11363
rect 37809 11295 37843 11323
rect 37809 11289 37843 11295
rect 37809 11227 37843 11251
rect 37809 11217 37843 11227
rect 37809 11159 37843 11179
rect 37809 11145 37843 11159
rect 37809 11091 37843 11107
rect 37809 11073 37843 11091
rect 37809 11023 37843 11035
rect 37809 11001 37843 11023
rect 37809 10955 37843 10963
rect 37809 10929 37843 10955
rect 38067 11873 38101 11899
rect 38067 11865 38101 11873
rect 38067 11805 38101 11827
rect 38067 11793 38101 11805
rect 38067 11737 38101 11755
rect 38067 11721 38101 11737
rect 38067 11669 38101 11683
rect 38067 11649 38101 11669
rect 38067 11601 38101 11611
rect 38067 11577 38101 11601
rect 38067 11533 38101 11539
rect 38067 11505 38101 11533
rect 38067 11465 38101 11467
rect 38067 11433 38101 11465
rect 38067 11363 38101 11395
rect 38067 11361 38101 11363
rect 38067 11295 38101 11323
rect 38067 11289 38101 11295
rect 38067 11227 38101 11251
rect 38067 11217 38101 11227
rect 38067 11159 38101 11179
rect 38067 11145 38101 11159
rect 38067 11091 38101 11107
rect 38067 11073 38101 11091
rect 38067 11023 38101 11035
rect 38067 11001 38101 11023
rect 38067 10955 38101 10963
rect 38067 10929 38101 10955
rect 38325 11873 38359 11899
rect 38325 11865 38359 11873
rect 38325 11805 38359 11827
rect 38325 11793 38359 11805
rect 38325 11737 38359 11755
rect 38325 11721 38359 11737
rect 38325 11669 38359 11683
rect 38325 11649 38359 11669
rect 38325 11601 38359 11611
rect 38325 11577 38359 11601
rect 38325 11533 38359 11539
rect 38325 11505 38359 11533
rect 38325 11465 38359 11467
rect 38325 11433 38359 11465
rect 38325 11363 38359 11395
rect 38325 11361 38359 11363
rect 38325 11295 38359 11323
rect 38325 11289 38359 11295
rect 38325 11227 38359 11251
rect 38325 11217 38359 11227
rect 38325 11159 38359 11179
rect 38325 11145 38359 11159
rect 38325 11091 38359 11107
rect 38325 11073 38359 11091
rect 38325 11023 38359 11035
rect 38325 11001 38359 11023
rect 38325 10955 38359 10963
rect 38325 10929 38359 10955
rect 38583 11873 38617 11899
rect 38583 11865 38617 11873
rect 38583 11805 38617 11827
rect 38583 11793 38617 11805
rect 38583 11737 38617 11755
rect 38583 11721 38617 11737
rect 38583 11669 38617 11683
rect 38583 11649 38617 11669
rect 38583 11601 38617 11611
rect 38583 11577 38617 11601
rect 38583 11533 38617 11539
rect 38583 11505 38617 11533
rect 38583 11465 38617 11467
rect 38583 11433 38617 11465
rect 38583 11363 38617 11395
rect 38583 11361 38617 11363
rect 38583 11295 38617 11323
rect 38583 11289 38617 11295
rect 38583 11227 38617 11251
rect 38583 11217 38617 11227
rect 38583 11159 38617 11179
rect 38583 11145 38617 11159
rect 38583 11091 38617 11107
rect 38583 11073 38617 11091
rect 38583 11023 38617 11035
rect 38583 11001 38617 11023
rect 38583 10955 38617 10963
rect 38583 10929 38617 10955
rect 38841 11873 38875 11899
rect 38841 11865 38875 11873
rect 38841 11805 38875 11827
rect 38841 11793 38875 11805
rect 38841 11737 38875 11755
rect 38841 11721 38875 11737
rect 38841 11669 38875 11683
rect 38841 11649 38875 11669
rect 38841 11601 38875 11611
rect 38841 11577 38875 11601
rect 38841 11533 38875 11539
rect 38841 11505 38875 11533
rect 38841 11465 38875 11467
rect 38841 11433 38875 11465
rect 38841 11363 38875 11395
rect 38841 11361 38875 11363
rect 38841 11295 38875 11323
rect 38841 11289 38875 11295
rect 38841 11227 38875 11251
rect 38841 11217 38875 11227
rect 38841 11159 38875 11179
rect 38841 11145 38875 11159
rect 38841 11091 38875 11107
rect 38841 11073 38875 11091
rect 38841 11023 38875 11035
rect 38841 11001 38875 11023
rect 38841 10955 38875 10963
rect 38841 10929 38875 10955
rect 39099 11873 39133 11899
rect 39099 11865 39133 11873
rect 39099 11805 39133 11827
rect 39099 11793 39133 11805
rect 39099 11737 39133 11755
rect 39099 11721 39133 11737
rect 39099 11669 39133 11683
rect 39099 11649 39133 11669
rect 39099 11601 39133 11611
rect 39099 11577 39133 11601
rect 39099 11533 39133 11539
rect 39099 11505 39133 11533
rect 39099 11465 39133 11467
rect 39099 11433 39133 11465
rect 39099 11363 39133 11395
rect 39099 11361 39133 11363
rect 39099 11295 39133 11323
rect 39099 11289 39133 11295
rect 39099 11227 39133 11251
rect 39099 11217 39133 11227
rect 39099 11159 39133 11179
rect 39099 11145 39133 11159
rect 39099 11091 39133 11107
rect 39099 11073 39133 11091
rect 39099 11023 39133 11035
rect 39099 11001 39133 11023
rect 39099 10955 39133 10963
rect 39099 10929 39133 10955
rect 39357 11873 39391 11899
rect 39357 11865 39391 11873
rect 39357 11805 39391 11827
rect 39357 11793 39391 11805
rect 39357 11737 39391 11755
rect 39357 11721 39391 11737
rect 39357 11669 39391 11683
rect 39357 11649 39391 11669
rect 39357 11601 39391 11611
rect 39357 11577 39391 11601
rect 39357 11533 39391 11539
rect 39357 11505 39391 11533
rect 39357 11465 39391 11467
rect 39357 11433 39391 11465
rect 39357 11363 39391 11395
rect 39357 11361 39391 11363
rect 39357 11295 39391 11323
rect 39357 11289 39391 11295
rect 39357 11227 39391 11251
rect 39357 11217 39391 11227
rect 39357 11159 39391 11179
rect 39357 11145 39391 11159
rect 39357 11091 39391 11107
rect 39357 11073 39391 11091
rect 39357 11023 39391 11035
rect 39357 11001 39391 11023
rect 39357 10955 39391 10963
rect 39357 10929 39391 10955
rect 39615 11873 39649 11899
rect 39615 11865 39649 11873
rect 39615 11805 39649 11827
rect 39615 11793 39649 11805
rect 39615 11737 39649 11755
rect 39615 11721 39649 11737
rect 39615 11669 39649 11683
rect 39615 11649 39649 11669
rect 39615 11601 39649 11611
rect 39615 11577 39649 11601
rect 39615 11533 39649 11539
rect 39615 11505 39649 11533
rect 39615 11465 39649 11467
rect 39615 11433 39649 11465
rect 39615 11363 39649 11395
rect 39615 11361 39649 11363
rect 39615 11295 39649 11323
rect 39615 11289 39649 11295
rect 39615 11227 39649 11251
rect 39615 11217 39649 11227
rect 39615 11159 39649 11179
rect 39615 11145 39649 11159
rect 39615 11091 39649 11107
rect 39615 11073 39649 11091
rect 39615 11023 39649 11035
rect 39615 11001 39649 11023
rect 39615 10955 39649 10963
rect 39615 10929 39649 10955
rect 39873 11873 39907 11899
rect 39873 11865 39907 11873
rect 39873 11805 39907 11827
rect 39873 11793 39907 11805
rect 39873 11737 39907 11755
rect 39873 11721 39907 11737
rect 39873 11669 39907 11683
rect 39873 11649 39907 11669
rect 39873 11601 39907 11611
rect 39873 11577 39907 11601
rect 39873 11533 39907 11539
rect 39873 11505 39907 11533
rect 39873 11465 39907 11467
rect 39873 11433 39907 11465
rect 39873 11363 39907 11395
rect 39873 11361 39907 11363
rect 39873 11295 39907 11323
rect 39873 11289 39907 11295
rect 39873 11227 39907 11251
rect 39873 11217 39907 11227
rect 39873 11159 39907 11179
rect 39873 11145 39907 11159
rect 39873 11091 39907 11107
rect 39873 11073 39907 11091
rect 39873 11023 39907 11035
rect 39873 11001 39907 11023
rect 39873 10955 39907 10963
rect 39873 10929 39907 10955
rect 40131 11873 40165 11899
rect 40131 11865 40165 11873
rect 40131 11805 40165 11827
rect 40131 11793 40165 11805
rect 40131 11737 40165 11755
rect 40131 11721 40165 11737
rect 40131 11669 40165 11683
rect 40131 11649 40165 11669
rect 40131 11601 40165 11611
rect 40131 11577 40165 11601
rect 40131 11533 40165 11539
rect 40131 11505 40165 11533
rect 40131 11465 40165 11467
rect 40131 11433 40165 11465
rect 40131 11363 40165 11395
rect 40131 11361 40165 11363
rect 40131 11295 40165 11323
rect 40131 11289 40165 11295
rect 40131 11227 40165 11251
rect 40131 11217 40165 11227
rect 40131 11159 40165 11179
rect 40131 11145 40165 11159
rect 40131 11091 40165 11107
rect 40131 11073 40165 11091
rect 40131 11023 40165 11035
rect 40131 11001 40165 11023
rect 40131 10955 40165 10963
rect 40131 10929 40165 10955
rect 40389 11873 40423 11899
rect 40389 11865 40423 11873
rect 40389 11805 40423 11827
rect 40389 11793 40423 11805
rect 40389 11737 40423 11755
rect 40389 11721 40423 11737
rect 40389 11669 40423 11683
rect 40389 11649 40423 11669
rect 40389 11601 40423 11611
rect 40389 11577 40423 11601
rect 40389 11533 40423 11539
rect 40389 11505 40423 11533
rect 40389 11465 40423 11467
rect 40389 11433 40423 11465
rect 40389 11363 40423 11395
rect 40389 11361 40423 11363
rect 40389 11295 40423 11323
rect 40389 11289 40423 11295
rect 40389 11227 40423 11251
rect 40389 11217 40423 11227
rect 40389 11159 40423 11179
rect 40389 11145 40423 11159
rect 40389 11091 40423 11107
rect 40389 11073 40423 11091
rect 40389 11023 40423 11035
rect 40389 11001 40423 11023
rect 40389 10955 40423 10963
rect 40389 10929 40423 10955
rect 40647 11873 40681 11899
rect 40647 11865 40681 11873
rect 40647 11805 40681 11827
rect 40647 11793 40681 11805
rect 40647 11737 40681 11755
rect 40647 11721 40681 11737
rect 40647 11669 40681 11683
rect 40647 11649 40681 11669
rect 40647 11601 40681 11611
rect 40647 11577 40681 11601
rect 40647 11533 40681 11539
rect 40647 11505 40681 11533
rect 40647 11465 40681 11467
rect 40647 11433 40681 11465
rect 40647 11363 40681 11395
rect 40647 11361 40681 11363
rect 40647 11295 40681 11323
rect 40647 11289 40681 11295
rect 40647 11227 40681 11251
rect 40647 11217 40681 11227
rect 40647 11159 40681 11179
rect 40647 11145 40681 11159
rect 40647 11091 40681 11107
rect 40647 11073 40681 11091
rect 40647 11023 40681 11035
rect 40647 11001 40681 11023
rect 40647 10955 40681 10963
rect 40647 10929 40681 10955
rect 40905 11873 40939 11899
rect 40905 11865 40939 11873
rect 40905 11805 40939 11827
rect 40905 11793 40939 11805
rect 40905 11737 40939 11755
rect 40905 11721 40939 11737
rect 40905 11669 40939 11683
rect 40905 11649 40939 11669
rect 40905 11601 40939 11611
rect 40905 11577 40939 11601
rect 40905 11533 40939 11539
rect 40905 11505 40939 11533
rect 40905 11465 40939 11467
rect 40905 11433 40939 11465
rect 40905 11363 40939 11395
rect 40905 11361 40939 11363
rect 40905 11295 40939 11323
rect 40905 11289 40939 11295
rect 40905 11227 40939 11251
rect 40905 11217 40939 11227
rect 40905 11159 40939 11179
rect 40905 11145 40939 11159
rect 40905 11091 40939 11107
rect 40905 11073 40939 11091
rect 40905 11023 40939 11035
rect 40905 11001 40939 11023
rect 40905 10955 40939 10963
rect 40905 10929 40939 10955
rect 41163 11873 41197 11899
rect 41163 11865 41197 11873
rect 41163 11805 41197 11827
rect 41163 11793 41197 11805
rect 41163 11737 41197 11755
rect 41163 11721 41197 11737
rect 41163 11669 41197 11683
rect 41163 11649 41197 11669
rect 41163 11601 41197 11611
rect 41163 11577 41197 11601
rect 41163 11533 41197 11539
rect 41163 11505 41197 11533
rect 41163 11465 41197 11467
rect 41163 11433 41197 11465
rect 41163 11363 41197 11395
rect 41163 11361 41197 11363
rect 41163 11295 41197 11323
rect 41163 11289 41197 11295
rect 41163 11227 41197 11251
rect 41163 11217 41197 11227
rect 41163 11159 41197 11179
rect 41163 11145 41197 11159
rect 41163 11091 41197 11107
rect 41163 11073 41197 11091
rect 41163 11023 41197 11035
rect 41163 11001 41197 11023
rect 41163 10955 41197 10963
rect 41163 10929 41197 10955
rect 41421 11873 41455 11899
rect 41421 11865 41455 11873
rect 41421 11805 41455 11827
rect 41421 11793 41455 11805
rect 41421 11737 41455 11755
rect 41421 11721 41455 11737
rect 41421 11669 41455 11683
rect 41421 11649 41455 11669
rect 41421 11601 41455 11611
rect 41421 11577 41455 11601
rect 41421 11533 41455 11539
rect 41421 11505 41455 11533
rect 41421 11465 41455 11467
rect 41421 11433 41455 11465
rect 41421 11363 41455 11395
rect 41421 11361 41455 11363
rect 41421 11295 41455 11323
rect 41421 11289 41455 11295
rect 41421 11227 41455 11251
rect 41421 11217 41455 11227
rect 41421 11159 41455 11179
rect 41421 11145 41455 11159
rect 41421 11091 41455 11107
rect 41421 11073 41455 11091
rect 41421 11023 41455 11035
rect 41421 11001 41455 11023
rect 41421 10955 41455 10963
rect 41421 10929 41455 10955
rect 41679 11873 41713 11899
rect 41679 11865 41713 11873
rect 41679 11805 41713 11827
rect 41679 11793 41713 11805
rect 41679 11737 41713 11755
rect 41679 11721 41713 11737
rect 41679 11669 41713 11683
rect 41679 11649 41713 11669
rect 41679 11601 41713 11611
rect 41679 11577 41713 11601
rect 41679 11533 41713 11539
rect 41679 11505 41713 11533
rect 41679 11465 41713 11467
rect 41679 11433 41713 11465
rect 41679 11363 41713 11395
rect 41679 11361 41713 11363
rect 41679 11295 41713 11323
rect 41679 11289 41713 11295
rect 41679 11227 41713 11251
rect 41679 11217 41713 11227
rect 41679 11159 41713 11179
rect 41679 11145 41713 11159
rect 41679 11091 41713 11107
rect 41679 11073 41713 11091
rect 41679 11023 41713 11035
rect 41679 11001 41713 11023
rect 41679 10955 41713 10963
rect 41679 10929 41713 10955
rect 41937 11873 41971 11899
rect 41937 11865 41971 11873
rect 41937 11805 41971 11827
rect 41937 11793 41971 11805
rect 41937 11737 41971 11755
rect 41937 11721 41971 11737
rect 41937 11669 41971 11683
rect 41937 11649 41971 11669
rect 41937 11601 41971 11611
rect 41937 11577 41971 11601
rect 41937 11533 41971 11539
rect 41937 11505 41971 11533
rect 41937 11465 41971 11467
rect 41937 11433 41971 11465
rect 41937 11363 41971 11395
rect 41937 11361 41971 11363
rect 41937 11295 41971 11323
rect 41937 11289 41971 11295
rect 41937 11227 41971 11251
rect 41937 11217 41971 11227
rect 41937 11159 41971 11179
rect 41937 11145 41971 11159
rect 41937 11091 41971 11107
rect 41937 11073 41971 11091
rect 41937 11023 41971 11035
rect 41937 11001 41971 11023
rect 41937 10955 41971 10963
rect 41937 10929 41971 10955
rect 36870 10842 36872 10876
rect 36872 10842 36904 10876
rect 36942 10842 36974 10876
rect 36974 10842 36976 10876
rect 37128 10842 37130 10876
rect 37130 10842 37162 10876
rect 37200 10842 37232 10876
rect 37232 10842 37234 10876
rect 37386 10842 37388 10876
rect 37388 10842 37420 10876
rect 37458 10842 37490 10876
rect 37490 10842 37492 10876
rect 37644 10842 37646 10876
rect 37646 10842 37678 10876
rect 37716 10842 37748 10876
rect 37748 10842 37750 10876
rect 37902 10842 37904 10876
rect 37904 10842 37936 10876
rect 37974 10842 38006 10876
rect 38006 10842 38008 10876
rect 38160 10842 38162 10876
rect 38162 10842 38194 10876
rect 38232 10842 38264 10876
rect 38264 10842 38266 10876
rect 38418 10842 38420 10876
rect 38420 10842 38452 10876
rect 38490 10842 38522 10876
rect 38522 10842 38524 10876
rect 38676 10842 38678 10876
rect 38678 10842 38710 10876
rect 38748 10842 38780 10876
rect 38780 10842 38782 10876
rect 38934 10842 38936 10876
rect 38936 10842 38968 10876
rect 39006 10842 39038 10876
rect 39038 10842 39040 10876
rect 39192 10842 39194 10876
rect 39194 10842 39226 10876
rect 39264 10842 39296 10876
rect 39296 10842 39298 10876
rect 39450 10842 39452 10876
rect 39452 10842 39484 10876
rect 39522 10842 39554 10876
rect 39554 10842 39556 10876
rect 39708 10842 39710 10876
rect 39710 10842 39742 10876
rect 39780 10842 39812 10876
rect 39812 10842 39814 10876
rect 39966 10842 39968 10876
rect 39968 10842 40000 10876
rect 40038 10842 40070 10876
rect 40070 10842 40072 10876
rect 40224 10842 40226 10876
rect 40226 10842 40258 10876
rect 40296 10842 40328 10876
rect 40328 10842 40330 10876
rect 40482 10842 40484 10876
rect 40484 10842 40516 10876
rect 40554 10842 40586 10876
rect 40586 10842 40588 10876
rect 40740 10842 40742 10876
rect 40742 10842 40774 10876
rect 40812 10842 40844 10876
rect 40844 10842 40846 10876
rect 40998 10842 41000 10876
rect 41000 10842 41032 10876
rect 41070 10842 41102 10876
rect 41102 10842 41104 10876
rect 41256 10842 41258 10876
rect 41258 10842 41290 10876
rect 41328 10842 41360 10876
rect 41360 10842 41362 10876
rect 41514 10842 41516 10876
rect 41516 10842 41548 10876
rect 41586 10842 41618 10876
rect 41618 10842 41620 10876
rect 41772 10842 41774 10876
rect 41774 10842 41806 10876
rect 41844 10842 41876 10876
rect 41876 10842 41878 10876
rect 37905 10587 37907 10621
rect 37907 10587 37939 10621
rect 37977 10587 38009 10621
rect 38009 10587 38011 10621
rect 38371 10587 38373 10621
rect 38373 10587 38405 10621
rect 38443 10587 38475 10621
rect 38475 10587 38477 10621
rect 38629 10587 38631 10621
rect 38631 10587 38663 10621
rect 38701 10587 38733 10621
rect 38733 10587 38735 10621
rect 38887 10587 38889 10621
rect 38889 10587 38921 10621
rect 38959 10587 38991 10621
rect 38991 10587 38993 10621
rect 39145 10587 39147 10621
rect 39147 10587 39179 10621
rect 39217 10587 39249 10621
rect 39249 10587 39251 10621
rect 39403 10587 39405 10621
rect 39405 10587 39437 10621
rect 39475 10587 39507 10621
rect 39507 10587 39509 10621
rect 39661 10587 39663 10621
rect 39663 10587 39695 10621
rect 39733 10587 39765 10621
rect 39765 10587 39767 10621
rect 39919 10587 39921 10621
rect 39921 10587 39953 10621
rect 39991 10587 40023 10621
rect 40023 10587 40025 10621
rect 40177 10587 40179 10621
rect 40179 10587 40211 10621
rect 40249 10587 40281 10621
rect 40281 10587 40283 10621
rect 40435 10587 40437 10621
rect 40437 10587 40469 10621
rect 40507 10587 40539 10621
rect 40539 10587 40541 10621
rect 40693 10587 40695 10621
rect 40695 10587 40727 10621
rect 40765 10587 40797 10621
rect 40797 10587 40799 10621
rect 37812 10508 37846 10534
rect 37812 10500 37846 10508
rect 37812 10440 37846 10462
rect 37812 10428 37846 10440
rect 37812 10372 37846 10390
rect 37812 10356 37846 10372
rect 37812 10304 37846 10318
rect 37812 10284 37846 10304
rect 37812 10236 37846 10246
rect 37812 10212 37846 10236
rect 37812 10168 37846 10174
rect 37812 10140 37846 10168
rect 37812 10100 37846 10102
rect 37812 10068 37846 10100
rect 37812 9998 37846 10030
rect 37812 9996 37846 9998
rect 37812 9930 37846 9958
rect 37812 9924 37846 9930
rect 37812 9862 37846 9886
rect 37812 9852 37846 9862
rect 37812 9794 37846 9814
rect 37812 9780 37846 9794
rect 37812 9726 37846 9742
rect 37812 9708 37846 9726
rect 37812 9658 37846 9670
rect 37812 9636 37846 9658
rect 37812 9590 37846 9598
rect 37812 9564 37846 9590
rect 38070 10508 38104 10534
rect 38070 10500 38104 10508
rect 38070 10440 38104 10462
rect 38070 10428 38104 10440
rect 38070 10372 38104 10390
rect 38070 10356 38104 10372
rect 38070 10304 38104 10318
rect 38070 10284 38104 10304
rect 38070 10236 38104 10246
rect 38070 10212 38104 10236
rect 38070 10168 38104 10174
rect 38070 10140 38104 10168
rect 38070 10100 38104 10102
rect 38070 10068 38104 10100
rect 38070 9998 38104 10030
rect 38070 9996 38104 9998
rect 38070 9930 38104 9958
rect 38070 9924 38104 9930
rect 38070 9862 38104 9886
rect 38070 9852 38104 9862
rect 38070 9794 38104 9814
rect 38070 9780 38104 9794
rect 38070 9726 38104 9742
rect 38070 9708 38104 9726
rect 38070 9658 38104 9670
rect 38070 9636 38104 9658
rect 38070 9590 38104 9598
rect 38070 9564 38104 9590
rect 38278 10508 38312 10534
rect 38278 10500 38312 10508
rect 38278 10440 38312 10462
rect 38278 10428 38312 10440
rect 38278 10372 38312 10390
rect 38278 10356 38312 10372
rect 38278 10304 38312 10318
rect 38278 10284 38312 10304
rect 38278 10236 38312 10246
rect 38278 10212 38312 10236
rect 38278 10168 38312 10174
rect 38278 10140 38312 10168
rect 38278 10100 38312 10102
rect 38278 10068 38312 10100
rect 38278 9998 38312 10030
rect 38278 9996 38312 9998
rect 38278 9930 38312 9958
rect 38278 9924 38312 9930
rect 38278 9862 38312 9886
rect 38278 9852 38312 9862
rect 38278 9794 38312 9814
rect 38278 9780 38312 9794
rect 38278 9726 38312 9742
rect 38278 9708 38312 9726
rect 38278 9658 38312 9670
rect 38278 9636 38312 9658
rect 38278 9590 38312 9598
rect 38278 9564 38312 9590
rect 38536 10508 38570 10534
rect 38536 10500 38570 10508
rect 38536 10440 38570 10462
rect 38536 10428 38570 10440
rect 38536 10372 38570 10390
rect 38536 10356 38570 10372
rect 38536 10304 38570 10318
rect 38536 10284 38570 10304
rect 38536 10236 38570 10246
rect 38536 10212 38570 10236
rect 38536 10168 38570 10174
rect 38536 10140 38570 10168
rect 38536 10100 38570 10102
rect 38536 10068 38570 10100
rect 38536 9998 38570 10030
rect 38536 9996 38570 9998
rect 38536 9930 38570 9958
rect 38536 9924 38570 9930
rect 38536 9862 38570 9886
rect 38536 9852 38570 9862
rect 38536 9794 38570 9814
rect 38536 9780 38570 9794
rect 38536 9726 38570 9742
rect 38536 9708 38570 9726
rect 38536 9658 38570 9670
rect 38536 9636 38570 9658
rect 38536 9590 38570 9598
rect 38536 9564 38570 9590
rect 38794 10508 38828 10534
rect 38794 10500 38828 10508
rect 38794 10440 38828 10462
rect 38794 10428 38828 10440
rect 38794 10372 38828 10390
rect 38794 10356 38828 10372
rect 38794 10304 38828 10318
rect 38794 10284 38828 10304
rect 38794 10236 38828 10246
rect 38794 10212 38828 10236
rect 38794 10168 38828 10174
rect 38794 10140 38828 10168
rect 38794 10100 38828 10102
rect 38794 10068 38828 10100
rect 38794 9998 38828 10030
rect 38794 9996 38828 9998
rect 38794 9930 38828 9958
rect 38794 9924 38828 9930
rect 38794 9862 38828 9886
rect 38794 9852 38828 9862
rect 38794 9794 38828 9814
rect 38794 9780 38828 9794
rect 38794 9726 38828 9742
rect 38794 9708 38828 9726
rect 38794 9658 38828 9670
rect 38794 9636 38828 9658
rect 38794 9590 38828 9598
rect 38794 9564 38828 9590
rect 39052 10508 39086 10534
rect 39052 10500 39086 10508
rect 39052 10440 39086 10462
rect 39052 10428 39086 10440
rect 39052 10372 39086 10390
rect 39052 10356 39086 10372
rect 39052 10304 39086 10318
rect 39052 10284 39086 10304
rect 39052 10236 39086 10246
rect 39052 10212 39086 10236
rect 39052 10168 39086 10174
rect 39052 10140 39086 10168
rect 39052 10100 39086 10102
rect 39052 10068 39086 10100
rect 39052 9998 39086 10030
rect 39052 9996 39086 9998
rect 39052 9930 39086 9958
rect 39052 9924 39086 9930
rect 39052 9862 39086 9886
rect 39052 9852 39086 9862
rect 39052 9794 39086 9814
rect 39052 9780 39086 9794
rect 39052 9726 39086 9742
rect 39052 9708 39086 9726
rect 39052 9658 39086 9670
rect 39052 9636 39086 9658
rect 39052 9590 39086 9598
rect 39052 9564 39086 9590
rect 39310 10508 39344 10534
rect 39310 10500 39344 10508
rect 39310 10440 39344 10462
rect 39310 10428 39344 10440
rect 39310 10372 39344 10390
rect 39310 10356 39344 10372
rect 39310 10304 39344 10318
rect 39310 10284 39344 10304
rect 39310 10236 39344 10246
rect 39310 10212 39344 10236
rect 39310 10168 39344 10174
rect 39310 10140 39344 10168
rect 39310 10100 39344 10102
rect 39310 10068 39344 10100
rect 39310 9998 39344 10030
rect 39310 9996 39344 9998
rect 39310 9930 39344 9958
rect 39310 9924 39344 9930
rect 39310 9862 39344 9886
rect 39310 9852 39344 9862
rect 39310 9794 39344 9814
rect 39310 9780 39344 9794
rect 39310 9726 39344 9742
rect 39310 9708 39344 9726
rect 39310 9658 39344 9670
rect 39310 9636 39344 9658
rect 39310 9590 39344 9598
rect 39310 9564 39344 9590
rect 39568 10508 39602 10534
rect 39568 10500 39602 10508
rect 39568 10440 39602 10462
rect 39568 10428 39602 10440
rect 39568 10372 39602 10390
rect 39568 10356 39602 10372
rect 39568 10304 39602 10318
rect 39568 10284 39602 10304
rect 39568 10236 39602 10246
rect 39568 10212 39602 10236
rect 39568 10168 39602 10174
rect 39568 10140 39602 10168
rect 39568 10100 39602 10102
rect 39568 10068 39602 10100
rect 39568 9998 39602 10030
rect 39568 9996 39602 9998
rect 39568 9930 39602 9958
rect 39568 9924 39602 9930
rect 39568 9862 39602 9886
rect 39568 9852 39602 9862
rect 39568 9794 39602 9814
rect 39568 9780 39602 9794
rect 39568 9726 39602 9742
rect 39568 9708 39602 9726
rect 39568 9658 39602 9670
rect 39568 9636 39602 9658
rect 39568 9590 39602 9598
rect 39568 9564 39602 9590
rect 39826 10508 39860 10534
rect 39826 10500 39860 10508
rect 39826 10440 39860 10462
rect 39826 10428 39860 10440
rect 39826 10372 39860 10390
rect 39826 10356 39860 10372
rect 39826 10304 39860 10318
rect 39826 10284 39860 10304
rect 39826 10236 39860 10246
rect 39826 10212 39860 10236
rect 39826 10168 39860 10174
rect 39826 10140 39860 10168
rect 39826 10100 39860 10102
rect 39826 10068 39860 10100
rect 39826 9998 39860 10030
rect 39826 9996 39860 9998
rect 39826 9930 39860 9958
rect 39826 9924 39860 9930
rect 39826 9862 39860 9886
rect 39826 9852 39860 9862
rect 39826 9794 39860 9814
rect 39826 9780 39860 9794
rect 39826 9726 39860 9742
rect 39826 9708 39860 9726
rect 39826 9658 39860 9670
rect 39826 9636 39860 9658
rect 39826 9590 39860 9598
rect 39826 9564 39860 9590
rect 40084 10508 40118 10534
rect 40084 10500 40118 10508
rect 40084 10440 40118 10462
rect 40084 10428 40118 10440
rect 40084 10372 40118 10390
rect 40084 10356 40118 10372
rect 40084 10304 40118 10318
rect 40084 10284 40118 10304
rect 40084 10236 40118 10246
rect 40084 10212 40118 10236
rect 40084 10168 40118 10174
rect 40084 10140 40118 10168
rect 40084 10100 40118 10102
rect 40084 10068 40118 10100
rect 40084 9998 40118 10030
rect 40084 9996 40118 9998
rect 40084 9930 40118 9958
rect 40084 9924 40118 9930
rect 40084 9862 40118 9886
rect 40084 9852 40118 9862
rect 40084 9794 40118 9814
rect 40084 9780 40118 9794
rect 40084 9726 40118 9742
rect 40084 9708 40118 9726
rect 40084 9658 40118 9670
rect 40084 9636 40118 9658
rect 40084 9590 40118 9598
rect 40084 9564 40118 9590
rect 40342 10508 40376 10534
rect 40342 10500 40376 10508
rect 40342 10440 40376 10462
rect 40342 10428 40376 10440
rect 40342 10372 40376 10390
rect 40342 10356 40376 10372
rect 40342 10304 40376 10318
rect 40342 10284 40376 10304
rect 40342 10236 40376 10246
rect 40342 10212 40376 10236
rect 40342 10168 40376 10174
rect 40342 10140 40376 10168
rect 40342 10100 40376 10102
rect 40342 10068 40376 10100
rect 40342 9998 40376 10030
rect 40342 9996 40376 9998
rect 40342 9930 40376 9958
rect 40342 9924 40376 9930
rect 40342 9862 40376 9886
rect 40342 9852 40376 9862
rect 40342 9794 40376 9814
rect 40342 9780 40376 9794
rect 40342 9726 40376 9742
rect 40342 9708 40376 9726
rect 40342 9658 40376 9670
rect 40342 9636 40376 9658
rect 40342 9590 40376 9598
rect 40342 9564 40376 9590
rect 40600 10508 40634 10534
rect 40600 10500 40634 10508
rect 40600 10440 40634 10462
rect 40600 10428 40634 10440
rect 40600 10372 40634 10390
rect 40600 10356 40634 10372
rect 40600 10304 40634 10318
rect 40600 10284 40634 10304
rect 40600 10236 40634 10246
rect 40600 10212 40634 10236
rect 40600 10168 40634 10174
rect 40600 10140 40634 10168
rect 40600 10100 40634 10102
rect 40600 10068 40634 10100
rect 40600 9998 40634 10030
rect 40600 9996 40634 9998
rect 40600 9930 40634 9958
rect 40600 9924 40634 9930
rect 40600 9862 40634 9886
rect 40600 9852 40634 9862
rect 40600 9794 40634 9814
rect 40600 9780 40634 9794
rect 40600 9726 40634 9742
rect 40600 9708 40634 9726
rect 40600 9658 40634 9670
rect 40600 9636 40634 9658
rect 40600 9590 40634 9598
rect 40600 9564 40634 9590
rect 40858 10508 40892 10534
rect 40858 10500 40892 10508
rect 40858 10440 40892 10462
rect 40858 10428 40892 10440
rect 40858 10372 40892 10390
rect 40858 10356 40892 10372
rect 40858 10304 40892 10318
rect 40858 10284 40892 10304
rect 40858 10236 40892 10246
rect 40858 10212 40892 10236
rect 40858 10168 40892 10174
rect 40858 10140 40892 10168
rect 40858 10100 40892 10102
rect 40858 10068 40892 10100
rect 40858 9998 40892 10030
rect 40858 9996 40892 9998
rect 40858 9930 40892 9958
rect 40858 9924 40892 9930
rect 40858 9862 40892 9886
rect 40858 9852 40892 9862
rect 40858 9794 40892 9814
rect 40858 9780 40892 9794
rect 40858 9726 40892 9742
rect 40858 9708 40892 9726
rect 40858 9658 40892 9670
rect 40858 9636 40892 9658
rect 40858 9590 40892 9598
rect 40858 9564 40892 9590
rect 37905 9477 37907 9511
rect 37907 9477 37939 9511
rect 37977 9477 38009 9511
rect 38009 9477 38011 9511
rect 38371 9477 38373 9511
rect 38373 9477 38405 9511
rect 38443 9477 38475 9511
rect 38475 9477 38477 9511
rect 38629 9477 38631 9511
rect 38631 9477 38663 9511
rect 38701 9477 38733 9511
rect 38733 9477 38735 9511
rect 38887 9477 38889 9511
rect 38889 9477 38921 9511
rect 38959 9477 38991 9511
rect 38991 9477 38993 9511
rect 39145 9477 39147 9511
rect 39147 9477 39179 9511
rect 39217 9477 39249 9511
rect 39249 9477 39251 9511
rect 39403 9477 39405 9511
rect 39405 9477 39437 9511
rect 39475 9477 39507 9511
rect 39507 9477 39509 9511
rect 39661 9477 39663 9511
rect 39663 9477 39695 9511
rect 39733 9477 39765 9511
rect 39765 9477 39767 9511
rect 39919 9477 39921 9511
rect 39921 9477 39953 9511
rect 39991 9477 40023 9511
rect 40023 9477 40025 9511
rect 40177 9477 40179 9511
rect 40179 9477 40211 9511
rect 40249 9477 40281 9511
rect 40281 9477 40283 9511
rect 40435 9477 40437 9511
rect 40437 9477 40469 9511
rect 40507 9477 40539 9511
rect 40539 9477 40541 9511
rect 40693 9477 40695 9511
rect 40695 9477 40727 9511
rect 40765 9477 40797 9511
rect 40797 9477 40799 9511
rect 27718 6843 27752 6877
rect 27718 6771 27752 6805
rect 27718 6699 27752 6733
rect 27718 6627 27752 6661
rect 27718 6555 27752 6589
rect 24389 3480 24399 3504
rect 24399 3480 24423 3504
rect 24461 3480 24467 3504
rect 24467 3480 24495 3504
rect 27718 6483 27752 6517
rect 28036 6843 28070 6877
rect 28036 6771 28070 6805
rect 28036 6699 28070 6733
rect 28036 6627 28070 6661
rect 28036 6555 28070 6589
rect 28036 6483 28070 6517
rect 28354 6843 28388 6877
rect 28354 6771 28388 6805
rect 28354 6699 28388 6733
rect 28354 6627 28388 6661
rect 28354 6555 28388 6589
rect 28354 6483 28388 6517
rect 28672 6843 28706 6877
rect 28672 6771 28706 6805
rect 28672 6699 28706 6733
rect 28672 6627 28706 6661
rect 28672 6555 28706 6589
rect 28672 6483 28706 6517
rect 28990 6843 29024 6877
rect 28990 6771 29024 6805
rect 28990 6699 29024 6733
rect 28990 6627 29024 6661
rect 28990 6555 29024 6589
rect 28990 6483 29024 6517
rect 29308 6843 29342 6877
rect 29308 6771 29342 6805
rect 29308 6699 29342 6733
rect 29308 6627 29342 6661
rect 29308 6555 29342 6589
rect 29308 6483 29342 6517
rect 29626 6843 29660 6877
rect 29626 6771 29660 6805
rect 29626 6699 29660 6733
rect 29626 6627 29660 6661
rect 29626 6555 29660 6589
rect 29626 6483 29660 6517
rect 37905 8326 37907 8360
rect 37907 8326 37939 8360
rect 37977 8326 38009 8360
rect 38009 8326 38011 8360
rect 38163 8326 38165 8360
rect 38165 8326 38197 8360
rect 38235 8326 38267 8360
rect 38267 8326 38269 8360
rect 38421 8326 38423 8360
rect 38423 8326 38455 8360
rect 38493 8326 38525 8360
rect 38525 8326 38527 8360
rect 38679 8326 38681 8360
rect 38681 8326 38713 8360
rect 38751 8326 38783 8360
rect 38783 8326 38785 8360
rect 38937 8326 38939 8360
rect 38939 8326 38971 8360
rect 39009 8326 39041 8360
rect 39041 8326 39043 8360
rect 39195 8326 39197 8360
rect 39197 8326 39229 8360
rect 39267 8326 39299 8360
rect 39299 8326 39301 8360
rect 39453 8326 39455 8360
rect 39455 8326 39487 8360
rect 39525 8326 39557 8360
rect 39557 8326 39559 8360
rect 39711 8326 39713 8360
rect 39713 8326 39745 8360
rect 39783 8326 39815 8360
rect 39815 8326 39817 8360
rect 39969 8326 39971 8360
rect 39971 8326 40003 8360
rect 40041 8326 40073 8360
rect 40073 8326 40075 8360
rect 40227 8326 40229 8360
rect 40229 8326 40261 8360
rect 40299 8326 40331 8360
rect 40331 8326 40333 8360
rect 40485 8326 40487 8360
rect 40487 8326 40519 8360
rect 40557 8326 40589 8360
rect 40589 8326 40591 8360
rect 40743 8326 40745 8360
rect 40745 8326 40777 8360
rect 40815 8326 40847 8360
rect 40847 8326 40849 8360
rect 41001 8326 41003 8360
rect 41003 8326 41035 8360
rect 41073 8326 41105 8360
rect 41105 8326 41107 8360
rect 41259 8326 41261 8360
rect 41261 8326 41293 8360
rect 41331 8326 41363 8360
rect 41363 8326 41365 8360
rect 41517 8326 41519 8360
rect 41519 8326 41551 8360
rect 41589 8326 41621 8360
rect 41621 8326 41623 8360
rect 41775 8326 41777 8360
rect 41777 8326 41809 8360
rect 41847 8326 41879 8360
rect 41879 8326 41881 8360
rect 37623 6630 37624 6636
rect 37624 6630 37657 6636
rect 37623 6602 37657 6630
rect 37623 6562 37624 6564
rect 37624 6562 37657 6564
rect 37623 6530 37657 6562
rect 37623 6460 37657 6492
rect 37623 6458 37624 6460
rect 37624 6458 37657 6460
rect 37812 8223 37846 8241
rect 37812 8207 37846 8223
rect 37812 8155 37846 8169
rect 37812 8135 37846 8155
rect 37812 8087 37846 8097
rect 37812 8063 37846 8087
rect 37812 8019 37846 8025
rect 37812 7991 37846 8019
rect 37812 7951 37846 7953
rect 37812 7919 37846 7951
rect 37812 7849 37846 7881
rect 37812 7847 37846 7849
rect 37812 7781 37846 7809
rect 37812 7775 37846 7781
rect 37812 7713 37846 7737
rect 37812 7703 37846 7713
rect 37812 7645 37846 7665
rect 37812 7631 37846 7645
rect 37812 7577 37846 7593
rect 37812 7559 37846 7577
rect 37812 7509 37846 7521
rect 37812 7487 37846 7509
rect 37812 7441 37846 7449
rect 37812 7415 37846 7441
rect 37812 7373 37846 7377
rect 37812 7343 37846 7373
rect 37812 7271 37846 7305
rect 37812 7203 37846 7233
rect 37812 7199 37846 7203
rect 37812 7135 37846 7161
rect 37812 7127 37846 7135
rect 37812 7067 37846 7089
rect 37812 7055 37846 7067
rect 37812 6999 37846 7017
rect 37812 6983 37846 6999
rect 37812 6931 37846 6945
rect 37812 6911 37846 6931
rect 37812 6863 37846 6873
rect 37812 6839 37846 6863
rect 37812 6795 37846 6801
rect 37812 6767 37846 6795
rect 37812 6727 37846 6729
rect 37812 6695 37846 6727
rect 37812 6625 37846 6657
rect 37812 6623 37846 6625
rect 37812 6557 37846 6585
rect 37812 6551 37846 6557
rect 37812 6489 37846 6513
rect 37812 6479 37846 6489
rect 37812 6421 37846 6441
rect 37812 6407 37846 6421
rect 37812 6353 37846 6369
rect 37812 6335 37846 6353
rect 38070 8223 38104 8241
rect 38070 8207 38104 8223
rect 38070 8155 38104 8169
rect 38070 8135 38104 8155
rect 38070 8087 38104 8097
rect 38070 8063 38104 8087
rect 38070 8019 38104 8025
rect 38070 7991 38104 8019
rect 38070 7951 38104 7953
rect 38070 7919 38104 7951
rect 38070 7849 38104 7881
rect 38070 7847 38104 7849
rect 38070 7781 38104 7809
rect 38070 7775 38104 7781
rect 38070 7713 38104 7737
rect 38070 7703 38104 7713
rect 38070 7645 38104 7665
rect 38070 7631 38104 7645
rect 38070 7577 38104 7593
rect 38070 7559 38104 7577
rect 38070 7509 38104 7521
rect 38070 7487 38104 7509
rect 38070 7441 38104 7449
rect 38070 7415 38104 7441
rect 38070 7373 38104 7377
rect 38070 7343 38104 7373
rect 38070 7271 38104 7305
rect 38070 7203 38104 7233
rect 38070 7199 38104 7203
rect 38070 7135 38104 7161
rect 38070 7127 38104 7135
rect 38070 7067 38104 7089
rect 38070 7055 38104 7067
rect 38070 6999 38104 7017
rect 38070 6983 38104 6999
rect 38070 6931 38104 6945
rect 38070 6911 38104 6931
rect 38070 6863 38104 6873
rect 38070 6839 38104 6863
rect 38070 6795 38104 6801
rect 38070 6767 38104 6795
rect 38070 6727 38104 6729
rect 38070 6695 38104 6727
rect 38070 6625 38104 6657
rect 38070 6623 38104 6625
rect 38070 6557 38104 6585
rect 38070 6551 38104 6557
rect 38070 6489 38104 6513
rect 38070 6479 38104 6489
rect 38070 6421 38104 6441
rect 38070 6407 38104 6421
rect 38070 6353 38104 6369
rect 38070 6335 38104 6353
rect 38328 8223 38362 8241
rect 38328 8207 38362 8223
rect 38328 8155 38362 8169
rect 38328 8135 38362 8155
rect 38328 8087 38362 8097
rect 38328 8063 38362 8087
rect 38328 8019 38362 8025
rect 38328 7991 38362 8019
rect 38328 7951 38362 7953
rect 38328 7919 38362 7951
rect 38328 7849 38362 7881
rect 38328 7847 38362 7849
rect 38328 7781 38362 7809
rect 38328 7775 38362 7781
rect 38328 7713 38362 7737
rect 38328 7703 38362 7713
rect 38328 7645 38362 7665
rect 38328 7631 38362 7645
rect 38328 7577 38362 7593
rect 38328 7559 38362 7577
rect 38328 7509 38362 7521
rect 38328 7487 38362 7509
rect 38328 7441 38362 7449
rect 38328 7415 38362 7441
rect 38328 7373 38362 7377
rect 38328 7343 38362 7373
rect 38328 7271 38362 7305
rect 38328 7203 38362 7233
rect 38328 7199 38362 7203
rect 38328 7135 38362 7161
rect 38328 7127 38362 7135
rect 38328 7067 38362 7089
rect 38328 7055 38362 7067
rect 38328 6999 38362 7017
rect 38328 6983 38362 6999
rect 38328 6931 38362 6945
rect 38328 6911 38362 6931
rect 38328 6863 38362 6873
rect 38328 6839 38362 6863
rect 38328 6795 38362 6801
rect 38328 6767 38362 6795
rect 38328 6727 38362 6729
rect 38328 6695 38362 6727
rect 38328 6625 38362 6657
rect 38328 6623 38362 6625
rect 38328 6557 38362 6585
rect 38328 6551 38362 6557
rect 38328 6489 38362 6513
rect 38328 6479 38362 6489
rect 38328 6421 38362 6441
rect 38328 6407 38362 6421
rect 38328 6353 38362 6369
rect 38328 6335 38362 6353
rect 38586 8223 38620 8241
rect 38586 8207 38620 8223
rect 38586 8155 38620 8169
rect 38586 8135 38620 8155
rect 38586 8087 38620 8097
rect 38586 8063 38620 8087
rect 38586 8019 38620 8025
rect 38586 7991 38620 8019
rect 38586 7951 38620 7953
rect 38586 7919 38620 7951
rect 38586 7849 38620 7881
rect 38586 7847 38620 7849
rect 38586 7781 38620 7809
rect 38586 7775 38620 7781
rect 38586 7713 38620 7737
rect 38586 7703 38620 7713
rect 38586 7645 38620 7665
rect 38586 7631 38620 7645
rect 38586 7577 38620 7593
rect 38586 7559 38620 7577
rect 38586 7509 38620 7521
rect 38586 7487 38620 7509
rect 38586 7441 38620 7449
rect 38586 7415 38620 7441
rect 38586 7373 38620 7377
rect 38586 7343 38620 7373
rect 38586 7271 38620 7305
rect 38586 7203 38620 7233
rect 38586 7199 38620 7203
rect 38586 7135 38620 7161
rect 38586 7127 38620 7135
rect 38586 7067 38620 7089
rect 38586 7055 38620 7067
rect 38586 6999 38620 7017
rect 38586 6983 38620 6999
rect 38586 6931 38620 6945
rect 38586 6911 38620 6931
rect 38586 6863 38620 6873
rect 38586 6839 38620 6863
rect 38586 6795 38620 6801
rect 38586 6767 38620 6795
rect 38586 6727 38620 6729
rect 38586 6695 38620 6727
rect 38586 6625 38620 6657
rect 38586 6623 38620 6625
rect 38586 6557 38620 6585
rect 38586 6551 38620 6557
rect 38586 6489 38620 6513
rect 38586 6479 38620 6489
rect 38586 6421 38620 6441
rect 38586 6407 38620 6421
rect 38586 6353 38620 6369
rect 38586 6335 38620 6353
rect 38844 8223 38878 8241
rect 38844 8207 38878 8223
rect 38844 8155 38878 8169
rect 38844 8135 38878 8155
rect 38844 8087 38878 8097
rect 38844 8063 38878 8087
rect 38844 8019 38878 8025
rect 38844 7991 38878 8019
rect 38844 7951 38878 7953
rect 38844 7919 38878 7951
rect 38844 7849 38878 7881
rect 38844 7847 38878 7849
rect 38844 7781 38878 7809
rect 38844 7775 38878 7781
rect 38844 7713 38878 7737
rect 38844 7703 38878 7713
rect 38844 7645 38878 7665
rect 38844 7631 38878 7645
rect 38844 7577 38878 7593
rect 38844 7559 38878 7577
rect 38844 7509 38878 7521
rect 38844 7487 38878 7509
rect 38844 7441 38878 7449
rect 38844 7415 38878 7441
rect 38844 7373 38878 7377
rect 38844 7343 38878 7373
rect 38844 7271 38878 7305
rect 38844 7203 38878 7233
rect 38844 7199 38878 7203
rect 38844 7135 38878 7161
rect 38844 7127 38878 7135
rect 38844 7067 38878 7089
rect 38844 7055 38878 7067
rect 38844 6999 38878 7017
rect 38844 6983 38878 6999
rect 38844 6931 38878 6945
rect 38844 6911 38878 6931
rect 38844 6863 38878 6873
rect 38844 6839 38878 6863
rect 38844 6795 38878 6801
rect 38844 6767 38878 6795
rect 38844 6727 38878 6729
rect 38844 6695 38878 6727
rect 38844 6625 38878 6657
rect 38844 6623 38878 6625
rect 38844 6557 38878 6585
rect 38844 6551 38878 6557
rect 38844 6489 38878 6513
rect 38844 6479 38878 6489
rect 38844 6421 38878 6441
rect 38844 6407 38878 6421
rect 38844 6353 38878 6369
rect 38844 6335 38878 6353
rect 39102 8223 39136 8241
rect 39102 8207 39136 8223
rect 39102 8155 39136 8169
rect 39102 8135 39136 8155
rect 39102 8087 39136 8097
rect 39102 8063 39136 8087
rect 39102 8019 39136 8025
rect 39102 7991 39136 8019
rect 39102 7951 39136 7953
rect 39102 7919 39136 7951
rect 39102 7849 39136 7881
rect 39102 7847 39136 7849
rect 39102 7781 39136 7809
rect 39102 7775 39136 7781
rect 39102 7713 39136 7737
rect 39102 7703 39136 7713
rect 39102 7645 39136 7665
rect 39102 7631 39136 7645
rect 39102 7577 39136 7593
rect 39102 7559 39136 7577
rect 39102 7509 39136 7521
rect 39102 7487 39136 7509
rect 39102 7441 39136 7449
rect 39102 7415 39136 7441
rect 39102 7373 39136 7377
rect 39102 7343 39136 7373
rect 39102 7271 39136 7305
rect 39102 7203 39136 7233
rect 39102 7199 39136 7203
rect 39102 7135 39136 7161
rect 39102 7127 39136 7135
rect 39102 7067 39136 7089
rect 39102 7055 39136 7067
rect 39102 6999 39136 7017
rect 39102 6983 39136 6999
rect 39102 6931 39136 6945
rect 39102 6911 39136 6931
rect 39102 6863 39136 6873
rect 39102 6839 39136 6863
rect 39102 6795 39136 6801
rect 39102 6767 39136 6795
rect 39102 6727 39136 6729
rect 39102 6695 39136 6727
rect 39102 6625 39136 6657
rect 39102 6623 39136 6625
rect 39102 6557 39136 6585
rect 39102 6551 39136 6557
rect 39102 6489 39136 6513
rect 39102 6479 39136 6489
rect 39102 6421 39136 6441
rect 39102 6407 39136 6421
rect 39102 6353 39136 6369
rect 39102 6335 39136 6353
rect 39360 8223 39394 8241
rect 39360 8207 39394 8223
rect 39360 8155 39394 8169
rect 39360 8135 39394 8155
rect 39360 8087 39394 8097
rect 39360 8063 39394 8087
rect 39360 8019 39394 8025
rect 39360 7991 39394 8019
rect 39360 7951 39394 7953
rect 39360 7919 39394 7951
rect 39360 7849 39394 7881
rect 39360 7847 39394 7849
rect 39360 7781 39394 7809
rect 39360 7775 39394 7781
rect 39360 7713 39394 7737
rect 39360 7703 39394 7713
rect 39360 7645 39394 7665
rect 39360 7631 39394 7645
rect 39360 7577 39394 7593
rect 39360 7559 39394 7577
rect 39360 7509 39394 7521
rect 39360 7487 39394 7509
rect 39360 7441 39394 7449
rect 39360 7415 39394 7441
rect 39360 7373 39394 7377
rect 39360 7343 39394 7373
rect 39360 7271 39394 7305
rect 39360 7203 39394 7233
rect 39360 7199 39394 7203
rect 39360 7135 39394 7161
rect 39360 7127 39394 7135
rect 39360 7067 39394 7089
rect 39360 7055 39394 7067
rect 39360 6999 39394 7017
rect 39360 6983 39394 6999
rect 39360 6931 39394 6945
rect 39360 6911 39394 6931
rect 39360 6863 39394 6873
rect 39360 6839 39394 6863
rect 39360 6795 39394 6801
rect 39360 6767 39394 6795
rect 39360 6727 39394 6729
rect 39360 6695 39394 6727
rect 39360 6625 39394 6657
rect 39360 6623 39394 6625
rect 39360 6557 39394 6585
rect 39360 6551 39394 6557
rect 39360 6489 39394 6513
rect 39360 6479 39394 6489
rect 39360 6421 39394 6441
rect 39360 6407 39394 6421
rect 39360 6353 39394 6369
rect 39360 6335 39394 6353
rect 39618 8223 39652 8241
rect 39618 8207 39652 8223
rect 39618 8155 39652 8169
rect 39618 8135 39652 8155
rect 39618 8087 39652 8097
rect 39618 8063 39652 8087
rect 39618 8019 39652 8025
rect 39618 7991 39652 8019
rect 39618 7951 39652 7953
rect 39618 7919 39652 7951
rect 39618 7849 39652 7881
rect 39618 7847 39652 7849
rect 39618 7781 39652 7809
rect 39618 7775 39652 7781
rect 39618 7713 39652 7737
rect 39618 7703 39652 7713
rect 39618 7645 39652 7665
rect 39618 7631 39652 7645
rect 39618 7577 39652 7593
rect 39618 7559 39652 7577
rect 39618 7509 39652 7521
rect 39618 7487 39652 7509
rect 39618 7441 39652 7449
rect 39618 7415 39652 7441
rect 39618 7373 39652 7377
rect 39618 7343 39652 7373
rect 39618 7271 39652 7305
rect 39618 7203 39652 7233
rect 39618 7199 39652 7203
rect 39618 7135 39652 7161
rect 39618 7127 39652 7135
rect 39618 7067 39652 7089
rect 39618 7055 39652 7067
rect 39618 6999 39652 7017
rect 39618 6983 39652 6999
rect 39618 6931 39652 6945
rect 39618 6911 39652 6931
rect 39618 6863 39652 6873
rect 39618 6839 39652 6863
rect 39618 6795 39652 6801
rect 39618 6767 39652 6795
rect 39618 6727 39652 6729
rect 39618 6695 39652 6727
rect 39618 6625 39652 6657
rect 39618 6623 39652 6625
rect 39618 6557 39652 6585
rect 39618 6551 39652 6557
rect 39618 6489 39652 6513
rect 39618 6479 39652 6489
rect 39618 6421 39652 6441
rect 39618 6407 39652 6421
rect 39618 6353 39652 6369
rect 39618 6335 39652 6353
rect 39876 8223 39910 8241
rect 39876 8207 39910 8223
rect 39876 8155 39910 8169
rect 39876 8135 39910 8155
rect 39876 8087 39910 8097
rect 39876 8063 39910 8087
rect 39876 8019 39910 8025
rect 39876 7991 39910 8019
rect 39876 7951 39910 7953
rect 39876 7919 39910 7951
rect 39876 7849 39910 7881
rect 39876 7847 39910 7849
rect 39876 7781 39910 7809
rect 39876 7775 39910 7781
rect 39876 7713 39910 7737
rect 39876 7703 39910 7713
rect 39876 7645 39910 7665
rect 39876 7631 39910 7645
rect 39876 7577 39910 7593
rect 39876 7559 39910 7577
rect 39876 7509 39910 7521
rect 39876 7487 39910 7509
rect 39876 7441 39910 7449
rect 39876 7415 39910 7441
rect 39876 7373 39910 7377
rect 39876 7343 39910 7373
rect 39876 7271 39910 7305
rect 39876 7203 39910 7233
rect 39876 7199 39910 7203
rect 39876 7135 39910 7161
rect 39876 7127 39910 7135
rect 39876 7067 39910 7089
rect 39876 7055 39910 7067
rect 39876 6999 39910 7017
rect 39876 6983 39910 6999
rect 39876 6931 39910 6945
rect 39876 6911 39910 6931
rect 39876 6863 39910 6873
rect 39876 6839 39910 6863
rect 39876 6795 39910 6801
rect 39876 6767 39910 6795
rect 39876 6727 39910 6729
rect 39876 6695 39910 6727
rect 39876 6625 39910 6657
rect 39876 6623 39910 6625
rect 39876 6557 39910 6585
rect 39876 6551 39910 6557
rect 39876 6489 39910 6513
rect 39876 6479 39910 6489
rect 39876 6421 39910 6441
rect 39876 6407 39910 6421
rect 39876 6353 39910 6369
rect 39876 6335 39910 6353
rect 40134 8223 40168 8241
rect 40134 8207 40168 8223
rect 40134 8155 40168 8169
rect 40134 8135 40168 8155
rect 40134 8087 40168 8097
rect 40134 8063 40168 8087
rect 40134 8019 40168 8025
rect 40134 7991 40168 8019
rect 40134 7951 40168 7953
rect 40134 7919 40168 7951
rect 40134 7849 40168 7881
rect 40134 7847 40168 7849
rect 40134 7781 40168 7809
rect 40134 7775 40168 7781
rect 40134 7713 40168 7737
rect 40134 7703 40168 7713
rect 40134 7645 40168 7665
rect 40134 7631 40168 7645
rect 40134 7577 40168 7593
rect 40134 7559 40168 7577
rect 40134 7509 40168 7521
rect 40134 7487 40168 7509
rect 40134 7441 40168 7449
rect 40134 7415 40168 7441
rect 40134 7373 40168 7377
rect 40134 7343 40168 7373
rect 40134 7271 40168 7305
rect 40134 7203 40168 7233
rect 40134 7199 40168 7203
rect 40134 7135 40168 7161
rect 40134 7127 40168 7135
rect 40134 7067 40168 7089
rect 40134 7055 40168 7067
rect 40134 6999 40168 7017
rect 40134 6983 40168 6999
rect 40134 6931 40168 6945
rect 40134 6911 40168 6931
rect 40134 6863 40168 6873
rect 40134 6839 40168 6863
rect 40134 6795 40168 6801
rect 40134 6767 40168 6795
rect 40134 6727 40168 6729
rect 40134 6695 40168 6727
rect 40134 6625 40168 6657
rect 40134 6623 40168 6625
rect 40134 6557 40168 6585
rect 40134 6551 40168 6557
rect 40134 6489 40168 6513
rect 40134 6479 40168 6489
rect 40134 6421 40168 6441
rect 40134 6407 40168 6421
rect 40134 6353 40168 6369
rect 40134 6335 40168 6353
rect 40392 8223 40426 8241
rect 40392 8207 40426 8223
rect 40392 8155 40426 8169
rect 40392 8135 40426 8155
rect 40392 8087 40426 8097
rect 40392 8063 40426 8087
rect 40392 8019 40426 8025
rect 40392 7991 40426 8019
rect 40392 7951 40426 7953
rect 40392 7919 40426 7951
rect 40392 7849 40426 7881
rect 40392 7847 40426 7849
rect 40392 7781 40426 7809
rect 40392 7775 40426 7781
rect 40392 7713 40426 7737
rect 40392 7703 40426 7713
rect 40392 7645 40426 7665
rect 40392 7631 40426 7645
rect 40392 7577 40426 7593
rect 40392 7559 40426 7577
rect 40392 7509 40426 7521
rect 40392 7487 40426 7509
rect 40392 7441 40426 7449
rect 40392 7415 40426 7441
rect 40392 7373 40426 7377
rect 40392 7343 40426 7373
rect 40392 7271 40426 7305
rect 40392 7203 40426 7233
rect 40392 7199 40426 7203
rect 40392 7135 40426 7161
rect 40392 7127 40426 7135
rect 40392 7067 40426 7089
rect 40392 7055 40426 7067
rect 40392 6999 40426 7017
rect 40392 6983 40426 6999
rect 40392 6931 40426 6945
rect 40392 6911 40426 6931
rect 40392 6863 40426 6873
rect 40392 6839 40426 6863
rect 40392 6795 40426 6801
rect 40392 6767 40426 6795
rect 40392 6727 40426 6729
rect 40392 6695 40426 6727
rect 40392 6625 40426 6657
rect 40392 6623 40426 6625
rect 40392 6557 40426 6585
rect 40392 6551 40426 6557
rect 40392 6489 40426 6513
rect 40392 6479 40426 6489
rect 40392 6421 40426 6441
rect 40392 6407 40426 6421
rect 40392 6353 40426 6369
rect 40392 6335 40426 6353
rect 40650 8223 40684 8241
rect 40650 8207 40684 8223
rect 40650 8155 40684 8169
rect 40650 8135 40684 8155
rect 40650 8087 40684 8097
rect 40650 8063 40684 8087
rect 40650 8019 40684 8025
rect 40650 7991 40684 8019
rect 40650 7951 40684 7953
rect 40650 7919 40684 7951
rect 40650 7849 40684 7881
rect 40650 7847 40684 7849
rect 40650 7781 40684 7809
rect 40650 7775 40684 7781
rect 40650 7713 40684 7737
rect 40650 7703 40684 7713
rect 40650 7645 40684 7665
rect 40650 7631 40684 7645
rect 40650 7577 40684 7593
rect 40650 7559 40684 7577
rect 40650 7509 40684 7521
rect 40650 7487 40684 7509
rect 40650 7441 40684 7449
rect 40650 7415 40684 7441
rect 40650 7373 40684 7377
rect 40650 7343 40684 7373
rect 40650 7271 40684 7305
rect 40650 7203 40684 7233
rect 40650 7199 40684 7203
rect 40650 7135 40684 7161
rect 40650 7127 40684 7135
rect 40650 7067 40684 7089
rect 40650 7055 40684 7067
rect 40650 6999 40684 7017
rect 40650 6983 40684 6999
rect 40650 6931 40684 6945
rect 40650 6911 40684 6931
rect 40650 6863 40684 6873
rect 40650 6839 40684 6863
rect 40650 6795 40684 6801
rect 40650 6767 40684 6795
rect 40650 6727 40684 6729
rect 40650 6695 40684 6727
rect 40650 6625 40684 6657
rect 40650 6623 40684 6625
rect 40650 6557 40684 6585
rect 40650 6551 40684 6557
rect 40650 6489 40684 6513
rect 40650 6479 40684 6489
rect 40650 6421 40684 6441
rect 40650 6407 40684 6421
rect 40650 6353 40684 6369
rect 40650 6335 40684 6353
rect 40908 8223 40942 8241
rect 40908 8207 40942 8223
rect 40908 8155 40942 8169
rect 40908 8135 40942 8155
rect 40908 8087 40942 8097
rect 40908 8063 40942 8087
rect 40908 8019 40942 8025
rect 40908 7991 40942 8019
rect 40908 7951 40942 7953
rect 40908 7919 40942 7951
rect 40908 7849 40942 7881
rect 40908 7847 40942 7849
rect 40908 7781 40942 7809
rect 40908 7775 40942 7781
rect 40908 7713 40942 7737
rect 40908 7703 40942 7713
rect 40908 7645 40942 7665
rect 40908 7631 40942 7645
rect 40908 7577 40942 7593
rect 40908 7559 40942 7577
rect 40908 7509 40942 7521
rect 40908 7487 40942 7509
rect 40908 7441 40942 7449
rect 40908 7415 40942 7441
rect 40908 7373 40942 7377
rect 40908 7343 40942 7373
rect 40908 7271 40942 7305
rect 40908 7203 40942 7233
rect 40908 7199 40942 7203
rect 40908 7135 40942 7161
rect 40908 7127 40942 7135
rect 40908 7067 40942 7089
rect 40908 7055 40942 7067
rect 40908 6999 40942 7017
rect 40908 6983 40942 6999
rect 40908 6931 40942 6945
rect 40908 6911 40942 6931
rect 40908 6863 40942 6873
rect 40908 6839 40942 6863
rect 40908 6795 40942 6801
rect 40908 6767 40942 6795
rect 40908 6727 40942 6729
rect 40908 6695 40942 6727
rect 40908 6625 40942 6657
rect 40908 6623 40942 6625
rect 40908 6557 40942 6585
rect 40908 6551 40942 6557
rect 40908 6489 40942 6513
rect 40908 6479 40942 6489
rect 40908 6421 40942 6441
rect 40908 6407 40942 6421
rect 40908 6353 40942 6369
rect 40908 6335 40942 6353
rect 41166 8223 41200 8241
rect 41166 8207 41200 8223
rect 41166 8155 41200 8169
rect 41166 8135 41200 8155
rect 41166 8087 41200 8097
rect 41166 8063 41200 8087
rect 41166 8019 41200 8025
rect 41166 7991 41200 8019
rect 41166 7951 41200 7953
rect 41166 7919 41200 7951
rect 41166 7849 41200 7881
rect 41166 7847 41200 7849
rect 41166 7781 41200 7809
rect 41166 7775 41200 7781
rect 41166 7713 41200 7737
rect 41166 7703 41200 7713
rect 41166 7645 41200 7665
rect 41166 7631 41200 7645
rect 41166 7577 41200 7593
rect 41166 7559 41200 7577
rect 41166 7509 41200 7521
rect 41166 7487 41200 7509
rect 41166 7441 41200 7449
rect 41166 7415 41200 7441
rect 41166 7373 41200 7377
rect 41166 7343 41200 7373
rect 41166 7271 41200 7305
rect 41166 7203 41200 7233
rect 41166 7199 41200 7203
rect 41166 7135 41200 7161
rect 41166 7127 41200 7135
rect 41166 7067 41200 7089
rect 41166 7055 41200 7067
rect 41166 6999 41200 7017
rect 41166 6983 41200 6999
rect 41166 6931 41200 6945
rect 41166 6911 41200 6931
rect 41166 6863 41200 6873
rect 41166 6839 41200 6863
rect 41166 6795 41200 6801
rect 41166 6767 41200 6795
rect 41166 6727 41200 6729
rect 41166 6695 41200 6727
rect 41166 6625 41200 6657
rect 41166 6623 41200 6625
rect 41166 6557 41200 6585
rect 41166 6551 41200 6557
rect 41166 6489 41200 6513
rect 41166 6479 41200 6489
rect 41166 6421 41200 6441
rect 41166 6407 41200 6421
rect 41166 6353 41200 6369
rect 41166 6335 41200 6353
rect 41424 8223 41458 8241
rect 41424 8207 41458 8223
rect 41424 8155 41458 8169
rect 41424 8135 41458 8155
rect 41424 8087 41458 8097
rect 41424 8063 41458 8087
rect 41424 8019 41458 8025
rect 41424 7991 41458 8019
rect 41424 7951 41458 7953
rect 41424 7919 41458 7951
rect 41424 7849 41458 7881
rect 41424 7847 41458 7849
rect 41424 7781 41458 7809
rect 41424 7775 41458 7781
rect 41424 7713 41458 7737
rect 41424 7703 41458 7713
rect 41424 7645 41458 7665
rect 41424 7631 41458 7645
rect 41424 7577 41458 7593
rect 41424 7559 41458 7577
rect 41424 7509 41458 7521
rect 41424 7487 41458 7509
rect 41424 7441 41458 7449
rect 41424 7415 41458 7441
rect 41424 7373 41458 7377
rect 41424 7343 41458 7373
rect 41424 7271 41458 7305
rect 41424 7203 41458 7233
rect 41424 7199 41458 7203
rect 41424 7135 41458 7161
rect 41424 7127 41458 7135
rect 41424 7067 41458 7089
rect 41424 7055 41458 7067
rect 41424 6999 41458 7017
rect 41424 6983 41458 6999
rect 41424 6931 41458 6945
rect 41424 6911 41458 6931
rect 41424 6863 41458 6873
rect 41424 6839 41458 6863
rect 41424 6795 41458 6801
rect 41424 6767 41458 6795
rect 41424 6727 41458 6729
rect 41424 6695 41458 6727
rect 41424 6625 41458 6657
rect 41424 6623 41458 6625
rect 41424 6557 41458 6585
rect 41424 6551 41458 6557
rect 41424 6489 41458 6513
rect 41424 6479 41458 6489
rect 41424 6421 41458 6441
rect 41424 6407 41458 6421
rect 41424 6353 41458 6369
rect 41424 6335 41458 6353
rect 41682 8223 41716 8241
rect 41682 8207 41716 8223
rect 41682 8155 41716 8169
rect 41682 8135 41716 8155
rect 41682 8087 41716 8097
rect 41682 8063 41716 8087
rect 41682 8019 41716 8025
rect 41682 7991 41716 8019
rect 41682 7951 41716 7953
rect 41682 7919 41716 7951
rect 41682 7849 41716 7881
rect 41682 7847 41716 7849
rect 41682 7781 41716 7809
rect 41682 7775 41716 7781
rect 41682 7713 41716 7737
rect 41682 7703 41716 7713
rect 41682 7645 41716 7665
rect 41682 7631 41716 7645
rect 41682 7577 41716 7593
rect 41682 7559 41716 7577
rect 41682 7509 41716 7521
rect 41682 7487 41716 7509
rect 41682 7441 41716 7449
rect 41682 7415 41716 7441
rect 41682 7373 41716 7377
rect 41682 7343 41716 7373
rect 41682 7271 41716 7305
rect 41682 7203 41716 7233
rect 41682 7199 41716 7203
rect 41682 7135 41716 7161
rect 41682 7127 41716 7135
rect 41682 7067 41716 7089
rect 41682 7055 41716 7067
rect 41682 6999 41716 7017
rect 41682 6983 41716 6999
rect 41682 6931 41716 6945
rect 41682 6911 41716 6931
rect 41682 6863 41716 6873
rect 41682 6839 41716 6863
rect 41682 6795 41716 6801
rect 41682 6767 41716 6795
rect 41682 6727 41716 6729
rect 41682 6695 41716 6727
rect 41682 6625 41716 6657
rect 41682 6623 41716 6625
rect 41682 6557 41716 6585
rect 41682 6551 41716 6557
rect 41682 6489 41716 6513
rect 41682 6479 41716 6489
rect 41682 6421 41716 6441
rect 41682 6407 41716 6421
rect 41682 6353 41716 6369
rect 41682 6335 41716 6353
rect 41940 8223 41974 8241
rect 41940 8207 41974 8223
rect 41940 8155 41974 8169
rect 41940 8135 41974 8155
rect 41940 8087 41974 8097
rect 41940 8063 41974 8087
rect 41940 8019 41974 8025
rect 41940 7991 41974 8019
rect 41940 7951 41974 7953
rect 41940 7919 41974 7951
rect 41940 7849 41974 7881
rect 41940 7847 41974 7849
rect 41940 7781 41974 7809
rect 41940 7775 41974 7781
rect 41940 7713 41974 7737
rect 41940 7703 41974 7713
rect 41940 7645 41974 7665
rect 41940 7631 41974 7645
rect 41940 7577 41974 7593
rect 41940 7559 41974 7577
rect 41940 7509 41974 7521
rect 41940 7487 41974 7509
rect 41940 7441 41974 7449
rect 41940 7415 41974 7441
rect 41940 7373 41974 7377
rect 41940 7343 41974 7373
rect 41940 7271 41974 7305
rect 41940 7203 41974 7233
rect 41940 7199 41974 7203
rect 41940 7135 41974 7161
rect 41940 7127 41974 7135
rect 41940 7067 41974 7089
rect 41940 7055 41974 7067
rect 41940 6999 41974 7017
rect 41940 6983 41974 6999
rect 41940 6931 41974 6945
rect 41940 6911 41974 6931
rect 41940 6863 41974 6873
rect 41940 6839 41974 6863
rect 41940 6795 41974 6801
rect 41940 6767 41974 6795
rect 41940 6727 41974 6729
rect 41940 6695 41974 6727
rect 41940 6625 41974 6657
rect 41940 6623 41974 6625
rect 41940 6557 41974 6585
rect 41940 6551 41974 6557
rect 41940 6489 41974 6513
rect 41940 6479 41974 6489
rect 41940 6421 41974 6441
rect 41940 6407 41974 6421
rect 41940 6353 41974 6369
rect 41940 6335 41974 6353
rect 42136 6608 42170 6635
rect 42136 6601 42170 6608
rect 42136 6540 42170 6563
rect 42136 6529 42170 6540
rect 42136 6472 42170 6491
rect 42136 6457 42170 6472
rect 37905 6216 37907 6250
rect 37907 6216 37939 6250
rect 37977 6216 38009 6250
rect 38009 6216 38011 6250
rect 38163 6216 38165 6250
rect 38165 6216 38197 6250
rect 38235 6216 38267 6250
rect 38267 6216 38269 6250
rect 38421 6216 38423 6250
rect 38423 6216 38455 6250
rect 38493 6216 38525 6250
rect 38525 6216 38527 6250
rect 38679 6216 38681 6250
rect 38681 6216 38713 6250
rect 38751 6216 38783 6250
rect 38783 6216 38785 6250
rect 38937 6216 38939 6250
rect 38939 6216 38971 6250
rect 39009 6216 39041 6250
rect 39041 6216 39043 6250
rect 39195 6216 39197 6250
rect 39197 6216 39229 6250
rect 39267 6216 39299 6250
rect 39299 6216 39301 6250
rect 39453 6216 39455 6250
rect 39455 6216 39487 6250
rect 39525 6216 39557 6250
rect 39557 6216 39559 6250
rect 39711 6216 39713 6250
rect 39713 6216 39745 6250
rect 39783 6216 39815 6250
rect 39815 6216 39817 6250
rect 39969 6216 39971 6250
rect 39971 6216 40003 6250
rect 40041 6216 40073 6250
rect 40073 6216 40075 6250
rect 40227 6216 40229 6250
rect 40229 6216 40261 6250
rect 40299 6216 40331 6250
rect 40331 6216 40333 6250
rect 40485 6216 40487 6250
rect 40487 6216 40519 6250
rect 40557 6216 40589 6250
rect 40589 6216 40591 6250
rect 40743 6216 40745 6250
rect 40745 6216 40777 6250
rect 40815 6216 40847 6250
rect 40847 6216 40849 6250
rect 41001 6216 41003 6250
rect 41003 6216 41035 6250
rect 41073 6216 41105 6250
rect 41105 6216 41107 6250
rect 41259 6216 41261 6250
rect 41261 6216 41293 6250
rect 41331 6216 41363 6250
rect 41363 6216 41365 6250
rect 41517 6216 41519 6250
rect 41519 6216 41551 6250
rect 41589 6216 41621 6250
rect 41621 6216 41623 6250
rect 41775 6216 41777 6250
rect 41777 6216 41809 6250
rect 41847 6216 41879 6250
rect 41879 6216 41881 6250
rect 24389 3470 24423 3480
rect 24461 3470 24495 3480
rect 26546 3459 26580 3493
rect 26546 3387 26580 3421
rect 26546 3315 26580 3349
rect 26546 3243 26580 3277
rect 26546 3171 26580 3205
rect 26546 3099 26580 3133
rect 26864 3459 26898 3493
rect 26864 3387 26898 3421
rect 26864 3315 26898 3349
rect 26864 3243 26898 3277
rect 26864 3171 26898 3205
rect 26864 3099 26898 3133
rect 27182 3459 27216 3493
rect 27182 3387 27216 3421
rect 27182 3315 27216 3349
rect 27182 3243 27216 3277
rect 27182 3171 27216 3205
rect 27182 3099 27216 3133
rect -6980 -39 -5434 787
rect 38612 711 40158 1537
<< metal1 >>
rect 8036 24833 52616 24867
rect 8036 24117 8103 24833
rect -15372 23971 8103 24117
rect -15372 23151 -15293 23971
rect -14217 23963 8103 23971
rect -14217 23207 5874 23963
rect 6886 23885 8103 23963
rect 8987 24721 52616 24833
rect 8987 23901 30299 24721
rect 31375 24713 52616 24721
rect 31375 23957 51466 24713
rect 52478 23957 52616 24713
rect 31375 23901 52616 23957
rect 8987 23885 52616 23901
rect 6886 23843 52616 23885
rect 6886 23207 9062 23843
rect -14217 23151 9062 23207
rect -15372 23093 9062 23151
rect 10298 23028 50454 23039
rect 10282 23002 50454 23028
rect 10282 22289 10363 23002
rect -13158 22198 10363 22289
rect -13158 22185 3696 22198
rect -13158 22182 -4261 22185
rect -3579 22182 3696 22185
rect -13158 22132 -4266 22182
rect -13158 21376 -13012 22132
rect -12000 21376 -4266 22132
rect -13158 21362 -4266 21376
rect -3574 21378 3696 22182
rect 4772 22054 10363 22198
rect 11247 22948 50454 23002
rect 11247 22935 49288 22948
rect 11247 22932 41331 22935
rect 42013 22932 49288 22935
rect 11247 22882 41326 22932
rect 11247 22126 32580 22882
rect 33592 22126 41326 22882
rect 11247 22112 41326 22126
rect 42018 22128 49288 22932
rect 50364 22128 50454 22948
rect 42018 22112 50454 22128
rect 11247 22109 41331 22112
rect 42013 22109 50454 22112
rect 11247 22054 50454 22109
rect 4772 22015 50454 22054
rect 4772 21378 11306 22015
rect -3574 21362 11306 21378
rect -13158 21359 -4261 21362
rect -3579 21359 11306 21362
rect -13158 21265 11306 21359
rect 41500 19216 41794 19249
rect 41500 19215 41523 19216
rect 41767 19215 41794 19216
rect 41500 19037 41520 19215
rect 41770 19037 41794 19215
rect 43556 19204 43762 19252
rect 43556 19088 43599 19204
rect 43715 19088 43762 19204
rect 43556 19046 43762 19088
rect 41500 19036 41523 19037
rect 41767 19036 41794 19037
rect 41500 19003 41794 19036
rect 42690 18930 45215 18947
rect 42662 18924 45215 18930
rect 23225 18844 27838 18916
rect 42662 18890 42705 18924
rect 42739 18890 42777 18924
rect 42811 18897 42963 18924
rect 42811 18890 42854 18897
rect 42662 18884 42854 18890
rect 42920 18890 42963 18897
rect 42997 18890 43035 18924
rect 43069 18897 43221 18924
rect 43069 18890 43112 18897
rect 42920 18884 43112 18890
rect 43178 18890 43221 18897
rect 43255 18890 43293 18924
rect 43327 18897 43479 18924
rect 43327 18890 43370 18897
rect 43178 18884 43370 18890
rect 43436 18890 43479 18897
rect 43513 18890 43551 18924
rect 43585 18897 43737 18924
rect 43585 18890 43628 18897
rect 43436 18884 43628 18890
rect 43694 18890 43737 18897
rect 43771 18890 43809 18924
rect 43843 18897 43995 18924
rect 43843 18890 43886 18897
rect 43694 18884 43886 18890
rect 43952 18890 43995 18897
rect 44029 18890 44067 18924
rect 44101 18897 44253 18924
rect 44101 18890 44144 18897
rect 43952 18884 44144 18890
rect 44210 18890 44253 18897
rect 44287 18890 44325 18924
rect 44359 18897 44511 18924
rect 44359 18890 44402 18897
rect 44210 18884 44402 18890
rect 44468 18890 44511 18897
rect 44545 18890 44583 18924
rect 44617 18897 44769 18924
rect 44617 18890 44660 18897
rect 44468 18884 44660 18890
rect 44726 18890 44769 18897
rect 44803 18890 44841 18924
rect 44875 18897 45027 18924
rect 44875 18890 44918 18897
rect 44726 18884 44918 18890
rect 44984 18890 45027 18897
rect 45061 18890 45099 18924
rect 45133 18897 45215 18924
rect 45133 18890 45176 18897
rect 44984 18884 45176 18890
rect 23225 18828 24280 18844
rect 23225 18794 23273 18828
rect 23307 18794 23345 18828
rect 23379 18794 23417 18828
rect 23451 18794 23489 18828
rect 23523 18794 23561 18828
rect 23595 18794 23633 18828
rect 23667 18794 23705 18828
rect 23739 18794 23777 18828
rect 23811 18794 23849 18828
rect 23883 18794 23921 18828
rect 23955 18794 23993 18828
rect 24027 18794 24065 18828
rect 24099 18794 24137 18828
rect 24171 18794 24280 18828
rect 23225 18788 24280 18794
rect 24742 18828 25734 18844
rect 24742 18794 24789 18828
rect 24823 18794 24861 18828
rect 24895 18794 24933 18828
rect 24967 18794 25005 18828
rect 25039 18794 25077 18828
rect 25111 18794 25149 18828
rect 25183 18794 25221 18828
rect 25255 18794 25293 18828
rect 25327 18794 25365 18828
rect 25399 18794 25437 18828
rect 25471 18794 25509 18828
rect 25543 18794 25581 18828
rect 25615 18794 25653 18828
rect 25687 18794 25734 18828
rect 24742 18788 25734 18794
rect 25800 18828 26792 18844
rect 25800 18794 25847 18828
rect 25881 18794 25919 18828
rect 25953 18794 25991 18828
rect 26025 18794 26063 18828
rect 26097 18794 26135 18828
rect 26169 18794 26207 18828
rect 26241 18794 26279 18828
rect 26313 18794 26351 18828
rect 26385 18794 26423 18828
rect 26457 18794 26495 18828
rect 26529 18794 26567 18828
rect 26601 18794 26639 18828
rect 26673 18794 26711 18828
rect 26745 18794 26792 18828
rect 25800 18788 26792 18794
rect 26858 18834 27838 18844
rect 42873 18843 43003 18855
rect 43382 18843 43512 18855
rect 43897 18843 44027 18851
rect 26858 18828 27850 18834
rect 26858 18794 26905 18828
rect 26939 18794 26977 18828
rect 27011 18794 27049 18828
rect 27083 18794 27121 18828
rect 27155 18794 27193 18828
rect 27227 18794 27265 18828
rect 27299 18794 27337 18828
rect 27371 18794 27409 18828
rect 27443 18794 27481 18828
rect 27515 18794 27553 18828
rect 27587 18794 27625 18828
rect 27659 18794 27697 18828
rect 27731 18794 27769 18828
rect 27803 18794 27850 18828
rect 26858 18788 27850 18794
rect 42606 18796 42652 18843
rect 23170 18732 23216 18747
rect 23170 18698 23176 18732
rect 23210 18698 23216 18732
rect 23170 18660 23216 18698
rect 23170 18626 23176 18660
rect 23210 18626 23216 18660
rect 24222 18732 24280 18788
rect 42606 18762 42612 18796
rect 42646 18762 42652 18796
rect 24222 18698 24234 18732
rect 24268 18698 24280 18732
rect 24686 18720 24732 18747
rect 24686 18698 24692 18720
rect 24222 18660 24280 18698
rect 24222 18629 24234 18660
rect 23170 18588 23216 18626
rect 23170 18554 23176 18588
rect 23210 18554 23216 18588
rect 23170 18516 23216 18554
rect -4092 18466 -3798 18499
rect -4092 18465 -4069 18466
rect -3825 18465 -3798 18466
rect -4092 18287 -4072 18465
rect -3822 18287 -3798 18465
rect -2036 18454 -1830 18502
rect -2036 18338 -1993 18454
rect -1877 18338 -1830 18454
rect -2036 18296 -1830 18338
rect 23170 18482 23176 18516
rect 23210 18482 23216 18516
rect 23170 18444 23216 18482
rect 23170 18410 23176 18444
rect 23210 18410 23216 18444
rect 23170 18372 23216 18410
rect 23170 18338 23176 18372
rect 23210 18338 23216 18372
rect 23170 18300 23216 18338
rect -4092 18286 -4069 18287
rect -3825 18286 -3798 18287
rect -4092 18253 -3798 18286
rect 23170 18266 23176 18300
rect 23210 18266 23216 18300
rect 23170 18228 23216 18266
rect -2902 18180 -377 18197
rect -2930 18174 -377 18180
rect -2930 18140 -2887 18174
rect -2853 18140 -2815 18174
rect -2781 18147 -2629 18174
rect -2781 18140 -2738 18147
rect -2930 18134 -2738 18140
rect -2672 18140 -2629 18147
rect -2595 18140 -2557 18174
rect -2523 18147 -2371 18174
rect -2523 18140 -2480 18147
rect -2672 18134 -2480 18140
rect -2414 18140 -2371 18147
rect -2337 18140 -2299 18174
rect -2265 18147 -2113 18174
rect -2265 18140 -2222 18147
rect -2414 18134 -2222 18140
rect -2156 18140 -2113 18147
rect -2079 18140 -2041 18174
rect -2007 18147 -1855 18174
rect -2007 18140 -1964 18147
rect -2156 18134 -1964 18140
rect -1898 18140 -1855 18147
rect -1821 18140 -1783 18174
rect -1749 18147 -1597 18174
rect -1749 18140 -1706 18147
rect -1898 18134 -1706 18140
rect -1640 18140 -1597 18147
rect -1563 18140 -1525 18174
rect -1491 18147 -1339 18174
rect -1491 18140 -1448 18147
rect -1640 18134 -1448 18140
rect -1382 18140 -1339 18147
rect -1305 18140 -1267 18174
rect -1233 18147 -1081 18174
rect -1233 18140 -1190 18147
rect -1382 18134 -1190 18140
rect -1124 18140 -1081 18147
rect -1047 18140 -1009 18174
rect -975 18147 -823 18174
rect -975 18140 -932 18147
rect -1124 18134 -932 18140
rect -866 18140 -823 18147
rect -789 18140 -751 18174
rect -717 18147 -565 18174
rect -717 18140 -674 18147
rect -866 18134 -674 18140
rect -608 18140 -565 18147
rect -531 18140 -493 18174
rect -459 18147 -377 18174
rect 23170 18194 23176 18228
rect 23210 18194 23216 18228
rect 23170 18156 23216 18194
rect -459 18140 -416 18147
rect -608 18134 -416 18140
rect 23170 18122 23176 18156
rect 23210 18122 23216 18156
rect -2719 18093 -2589 18105
rect -2210 18093 -2080 18105
rect -1695 18093 -1565 18101
rect -2986 18046 -2940 18093
rect -2986 18012 -2980 18046
rect -2946 18012 -2940 18046
rect -2986 17974 -2940 18012
rect -2986 17940 -2980 17974
rect -2946 17940 -2940 17974
rect -2986 17902 -2940 17940
rect -2986 17868 -2980 17902
rect -2946 17868 -2940 17902
rect -2986 17830 -2940 17868
rect -2986 17796 -2980 17830
rect -2946 17796 -2940 17830
rect -2986 17758 -2940 17796
rect -2986 17724 -2980 17758
rect -2946 17724 -2940 17758
rect -2986 17686 -2940 17724
rect -2986 17652 -2980 17686
rect -2946 17652 -2940 17686
rect -2986 17614 -2940 17652
rect -6276 17550 -6096 17594
rect -6276 17498 -6244 17550
rect -6192 17498 -6180 17550
rect -6128 17498 -6096 17550
rect -6276 17454 -6096 17498
rect -2986 17580 -2980 17614
rect -2946 17580 -2940 17614
rect -2986 17542 -2940 17580
rect -2986 17508 -2980 17542
rect -2946 17508 -2940 17542
rect -2986 17470 -2940 17508
rect -2986 17436 -2980 17470
rect -2946 17436 -2940 17470
rect -2986 17398 -2940 17436
rect -2986 17364 -2980 17398
rect -2946 17364 -2940 17398
rect -2986 17326 -2940 17364
rect -6398 17305 -6206 17311
rect -6398 17271 -6355 17305
rect -6321 17271 -6283 17305
rect -6249 17271 -6206 17305
rect -6398 17265 -6206 17271
rect -6140 17305 -5948 17311
rect -6140 17271 -6097 17305
rect -6063 17271 -6025 17305
rect -5991 17271 -5948 17305
rect -6140 17265 -5948 17271
rect -2986 17292 -2980 17326
rect -2946 17292 -2940 17326
rect -2986 17254 -2940 17292
rect -6454 17209 -6408 17224
rect -6196 17214 -6150 17224
rect -6454 17175 -6448 17209
rect -6414 17175 -6408 17209
rect -6454 17137 -6408 17175
rect -6454 17103 -6448 17137
rect -6414 17103 -6408 17137
rect -6454 17065 -6408 17103
rect -6246 17209 -6116 17214
rect -6246 17175 -6190 17209
rect -6156 17175 -6116 17209
rect -6246 17123 -6207 17175
rect -6155 17123 -6116 17175
rect -6246 17103 -6190 17123
rect -6156 17103 -6116 17123
rect -6246 17084 -6116 17103
rect -5938 17209 -5892 17224
rect -5938 17175 -5932 17209
rect -5898 17175 -5892 17209
rect -5938 17137 -5892 17175
rect -5938 17103 -5932 17137
rect -5898 17103 -5892 17137
rect -6454 17031 -6448 17065
rect -6414 17031 -6408 17065
rect -6454 16993 -6408 17031
rect -6454 16959 -6448 16993
rect -6414 16959 -6408 16993
rect -6454 16921 -6408 16959
rect -6454 16887 -6448 16921
rect -6414 16887 -6408 16921
rect -6454 16849 -6408 16887
rect -6454 16815 -6448 16849
rect -6414 16815 -6408 16849
rect -6454 16777 -6408 16815
rect -6454 16743 -6448 16777
rect -6414 16743 -6408 16777
rect -6454 16705 -6408 16743
rect -6454 16671 -6448 16705
rect -6414 16671 -6408 16705
rect -6454 16633 -6408 16671
rect -6454 16599 -6448 16633
rect -6414 16599 -6408 16633
rect -6454 16561 -6408 16599
rect -6454 16527 -6448 16561
rect -6414 16527 -6408 16561
rect -6454 16489 -6408 16527
rect -6454 16455 -6448 16489
rect -6414 16455 -6408 16489
rect -6454 16417 -6408 16455
rect -6454 16383 -6448 16417
rect -6414 16383 -6408 16417
rect -6454 16345 -6408 16383
rect -6454 16311 -6448 16345
rect -6414 16311 -6408 16345
rect -6454 16273 -6408 16311
rect -6454 16254 -6448 16273
rect -6456 16239 -6448 16254
rect -6414 16254 -6408 16273
rect -6196 17065 -6150 17084
rect -6196 17031 -6190 17065
rect -6156 17031 -6150 17065
rect -6196 16993 -6150 17031
rect -6196 16959 -6190 16993
rect -6156 16959 -6150 16993
rect -6196 16921 -6150 16959
rect -6196 16887 -6190 16921
rect -6156 16887 -6150 16921
rect -6196 16849 -6150 16887
rect -6196 16815 -6190 16849
rect -6156 16815 -6150 16849
rect -6196 16777 -6150 16815
rect -6196 16743 -6190 16777
rect -6156 16743 -6150 16777
rect -6196 16705 -6150 16743
rect -6196 16671 -6190 16705
rect -6156 16671 -6150 16705
rect -6196 16633 -6150 16671
rect -6196 16599 -6190 16633
rect -6156 16599 -6150 16633
rect -6196 16561 -6150 16599
rect -6196 16527 -6190 16561
rect -6156 16527 -6150 16561
rect -6196 16489 -6150 16527
rect -6196 16455 -6190 16489
rect -6156 16455 -6150 16489
rect -6196 16417 -6150 16455
rect -6196 16383 -6190 16417
rect -6156 16383 -6150 16417
rect -6196 16345 -6150 16383
rect -6196 16311 -6190 16345
rect -6156 16311 -6150 16345
rect -6196 16273 -6150 16311
rect -6414 16239 -6396 16254
rect -6456 16184 -6396 16239
rect -6196 16239 -6190 16273
rect -6156 16239 -6150 16273
rect -6196 16224 -6150 16239
rect -5938 17065 -5892 17103
rect -5938 17031 -5932 17065
rect -5898 17031 -5892 17065
rect -5938 16993 -5892 17031
rect -5938 16959 -5932 16993
rect -5898 16959 -5892 16993
rect -5938 16921 -5892 16959
rect -5938 16887 -5932 16921
rect -5898 16887 -5892 16921
rect -5938 16849 -5892 16887
rect -5938 16815 -5932 16849
rect -5898 16815 -5892 16849
rect -5938 16777 -5892 16815
rect -5938 16743 -5932 16777
rect -5898 16743 -5892 16777
rect -5938 16705 -5892 16743
rect -5938 16671 -5932 16705
rect -5898 16671 -5892 16705
rect -5938 16633 -5892 16671
rect -5938 16599 -5932 16633
rect -5898 16599 -5892 16633
rect -5938 16561 -5892 16599
rect -5938 16527 -5932 16561
rect -5898 16527 -5892 16561
rect -5938 16489 -5892 16527
rect -5938 16455 -5932 16489
rect -5898 16455 -5892 16489
rect -5938 16417 -5892 16455
rect -5938 16383 -5932 16417
rect -5898 16394 -5892 16417
rect -2986 17220 -2980 17254
rect -2946 17220 -2940 17254
rect -2986 17182 -2940 17220
rect -2986 17148 -2980 17182
rect -2946 17148 -2940 17182
rect -2986 17110 -2940 17148
rect -2986 17076 -2980 17110
rect -2946 17076 -2940 17110
rect -2986 17038 -2940 17076
rect -2986 17004 -2980 17038
rect -2946 17004 -2940 17038
rect -2986 16966 -2940 17004
rect -2986 16932 -2980 16966
rect -2946 16932 -2940 16966
rect -2986 16894 -2940 16932
rect -2986 16860 -2980 16894
rect -2946 16860 -2940 16894
rect -2986 16822 -2940 16860
rect -2986 16788 -2980 16822
rect -2946 16788 -2940 16822
rect -2986 16750 -2940 16788
rect -2986 16716 -2980 16750
rect -2946 16716 -2940 16750
rect -2986 16678 -2940 16716
rect -2986 16644 -2980 16678
rect -2946 16644 -2940 16678
rect -2986 16606 -2940 16644
rect -2986 16572 -2980 16606
rect -2946 16572 -2940 16606
rect -2986 16534 -2940 16572
rect -2986 16500 -2980 16534
rect -2946 16500 -2940 16534
rect -2986 16462 -2940 16500
rect -2986 16428 -2980 16462
rect -2946 16428 -2940 16462
rect -5898 16393 -5626 16394
rect -5898 16383 -3776 16393
rect -5938 16367 -3776 16383
rect -5938 16345 -5866 16367
rect -5938 16311 -5932 16345
rect -5898 16311 -5866 16345
rect -5938 16273 -5866 16311
rect -5938 16239 -5932 16273
rect -5898 16251 -5866 16273
rect -5686 16251 -3776 16367
rect -5898 16239 -3776 16251
rect -5938 16224 -3776 16239
rect -5927 16220 -3776 16224
rect -6456 16177 -5946 16184
rect -6456 16143 -6355 16177
rect -6321 16143 -6283 16177
rect -6249 16143 -6097 16177
rect -6063 16143 -6025 16177
rect -5991 16143 -5946 16177
rect -6456 16134 -5946 16143
rect -6436 16105 -6196 16134
rect -6436 16053 -6369 16105
rect -6317 16053 -6305 16105
rect -6253 16053 -6196 16105
rect -6436 16034 -6196 16053
rect -3949 16016 -3776 16220
rect -2986 16390 -2940 16428
rect -2986 16356 -2980 16390
rect -2946 16368 -2940 16390
rect -2728 18075 -2589 18093
rect -2728 18046 -2682 18075
rect -2728 18012 -2722 18046
rect -2688 18023 -2682 18046
rect -2630 18023 -2589 18075
rect -2688 18012 -2589 18023
rect -2728 18011 -2589 18012
rect -2728 17974 -2682 18011
rect -2728 17940 -2722 17974
rect -2688 17959 -2682 17974
rect -2630 17959 -2589 18011
rect -2688 17947 -2589 17959
rect -2688 17940 -2682 17947
rect -2728 17902 -2682 17940
rect -2728 17868 -2722 17902
rect -2688 17895 -2682 17902
rect -2630 17895 -2589 17947
rect -2688 17868 -2589 17895
rect -2728 17864 -2589 17868
rect -2470 18046 -2424 18093
rect -2470 18012 -2464 18046
rect -2430 18012 -2424 18046
rect -2470 17974 -2424 18012
rect -2470 17940 -2464 17974
rect -2430 17940 -2424 17974
rect -2470 17902 -2424 17940
rect -2470 17868 -2464 17902
rect -2430 17868 -2424 17902
rect -2728 17830 -2682 17864
rect -2728 17796 -2722 17830
rect -2688 17796 -2682 17830
rect -2728 17758 -2682 17796
rect -2728 17724 -2722 17758
rect -2688 17724 -2682 17758
rect -2728 17686 -2682 17724
rect -2728 17652 -2722 17686
rect -2688 17652 -2682 17686
rect -2728 17614 -2682 17652
rect -2728 17580 -2722 17614
rect -2688 17580 -2682 17614
rect -2728 17542 -2682 17580
rect -2728 17508 -2722 17542
rect -2688 17508 -2682 17542
rect -2728 17470 -2682 17508
rect -2728 17436 -2722 17470
rect -2688 17436 -2682 17470
rect -2728 17398 -2682 17436
rect -2728 17364 -2722 17398
rect -2688 17364 -2682 17398
rect -2728 17326 -2682 17364
rect -2728 17292 -2722 17326
rect -2688 17292 -2682 17326
rect -2728 17254 -2682 17292
rect -2728 17220 -2722 17254
rect -2688 17220 -2682 17254
rect -2728 17182 -2682 17220
rect -2728 17148 -2722 17182
rect -2688 17148 -2682 17182
rect -2728 17110 -2682 17148
rect -2728 17076 -2722 17110
rect -2688 17076 -2682 17110
rect -2728 17038 -2682 17076
rect -2728 17004 -2722 17038
rect -2688 17004 -2682 17038
rect -2728 16966 -2682 17004
rect -2728 16932 -2722 16966
rect -2688 16932 -2682 16966
rect -2728 16894 -2682 16932
rect -2728 16860 -2722 16894
rect -2688 16860 -2682 16894
rect -2728 16822 -2682 16860
rect -2728 16788 -2722 16822
rect -2688 16788 -2682 16822
rect -2728 16750 -2682 16788
rect -2728 16716 -2722 16750
rect -2688 16716 -2682 16750
rect -2728 16678 -2682 16716
rect -2728 16644 -2722 16678
rect -2688 16644 -2682 16678
rect -2728 16606 -2682 16644
rect -2728 16572 -2722 16606
rect -2688 16572 -2682 16606
rect -2728 16534 -2682 16572
rect -2728 16500 -2722 16534
rect -2688 16500 -2682 16534
rect -2728 16462 -2682 16500
rect -2728 16428 -2722 16462
rect -2688 16428 -2682 16462
rect -2728 16390 -2682 16428
rect -2946 16356 -2841 16368
rect -2986 16338 -2841 16356
rect -2986 16318 -2934 16338
rect -2986 16284 -2980 16318
rect -2946 16286 -2934 16318
rect -2882 16286 -2841 16338
rect -2946 16284 -2841 16286
rect -2986 16274 -2841 16284
rect -2986 16246 -2934 16274
rect -2986 16212 -2980 16246
rect -2946 16222 -2934 16246
rect -2882 16222 -2841 16274
rect -2946 16212 -2841 16222
rect -2986 16210 -2841 16212
rect -2986 16174 -2934 16210
rect -2986 16140 -2980 16174
rect -2946 16158 -2934 16174
rect -2882 16158 -2841 16210
rect -2946 16140 -2841 16158
rect -2986 16127 -2841 16140
rect -2728 16356 -2722 16390
rect -2688 16356 -2682 16390
rect -2470 17830 -2424 17868
rect -2470 17796 -2464 17830
rect -2430 17796 -2424 17830
rect -2470 17758 -2424 17796
rect -2470 17724 -2464 17758
rect -2430 17724 -2424 17758
rect -2470 17686 -2424 17724
rect -2470 17652 -2464 17686
rect -2430 17652 -2424 17686
rect -2470 17614 -2424 17652
rect -2470 17580 -2464 17614
rect -2430 17580 -2424 17614
rect -2470 17542 -2424 17580
rect -2470 17508 -2464 17542
rect -2430 17508 -2424 17542
rect -2470 17470 -2424 17508
rect -2470 17436 -2464 17470
rect -2430 17436 -2424 17470
rect -2470 17398 -2424 17436
rect -2470 17364 -2464 17398
rect -2430 17364 -2424 17398
rect -2470 17326 -2424 17364
rect -2470 17292 -2464 17326
rect -2430 17292 -2424 17326
rect -2470 17254 -2424 17292
rect -2470 17220 -2464 17254
rect -2430 17220 -2424 17254
rect -2470 17182 -2424 17220
rect -2470 17148 -2464 17182
rect -2430 17148 -2424 17182
rect -2470 17110 -2424 17148
rect -2470 17076 -2464 17110
rect -2430 17076 -2424 17110
rect -2470 17038 -2424 17076
rect -2470 17004 -2464 17038
rect -2430 17004 -2424 17038
rect -2470 16966 -2424 17004
rect -2470 16932 -2464 16966
rect -2430 16932 -2424 16966
rect -2470 16894 -2424 16932
rect -2470 16860 -2464 16894
rect -2430 16860 -2424 16894
rect -2470 16822 -2424 16860
rect -2470 16788 -2464 16822
rect -2430 16788 -2424 16822
rect -2470 16750 -2424 16788
rect -2470 16716 -2464 16750
rect -2430 16716 -2424 16750
rect -2470 16678 -2424 16716
rect -2470 16644 -2464 16678
rect -2430 16644 -2424 16678
rect -2470 16606 -2424 16644
rect -2470 16572 -2464 16606
rect -2430 16572 -2424 16606
rect -2470 16534 -2424 16572
rect -2470 16500 -2464 16534
rect -2430 16500 -2424 16534
rect -2470 16462 -2424 16500
rect -2470 16428 -2464 16462
rect -2430 16428 -2424 16462
rect -2470 16390 -2424 16428
rect -2470 16364 -2464 16390
rect -2728 16318 -2682 16356
rect -2728 16284 -2722 16318
rect -2688 16284 -2682 16318
rect -2728 16246 -2682 16284
rect -2728 16212 -2722 16246
rect -2688 16212 -2682 16246
rect -2728 16174 -2682 16212
rect -2728 16140 -2722 16174
rect -2688 16140 -2682 16174
rect -2986 16093 -2940 16127
rect -2728 16093 -2682 16140
rect -2471 16356 -2464 16364
rect -2430 16364 -2424 16390
rect -2212 18075 -2080 18093
rect -2212 18046 -2173 18075
rect -2212 18012 -2206 18046
rect -2121 18023 -2080 18075
rect -2172 18012 -2080 18023
rect -2212 18011 -2080 18012
rect -2212 17974 -2173 18011
rect -2212 17940 -2206 17974
rect -2121 17959 -2080 18011
rect -2172 17947 -2080 17959
rect -2212 17902 -2173 17940
rect -2212 17868 -2206 17902
rect -2121 17895 -2080 17947
rect -2172 17868 -2080 17895
rect -2212 17864 -2080 17868
rect -1954 18046 -1908 18093
rect -1954 18012 -1948 18046
rect -1914 18012 -1908 18046
rect -1954 17974 -1908 18012
rect -1954 17940 -1948 17974
rect -1914 17940 -1908 17974
rect -1954 17902 -1908 17940
rect -1954 17868 -1948 17902
rect -1914 17868 -1908 17902
rect -2212 17830 -2166 17864
rect -2212 17796 -2206 17830
rect -2172 17796 -2166 17830
rect -2212 17758 -2166 17796
rect -2212 17724 -2206 17758
rect -2172 17724 -2166 17758
rect -2212 17686 -2166 17724
rect -2212 17652 -2206 17686
rect -2172 17652 -2166 17686
rect -2212 17614 -2166 17652
rect -2212 17580 -2206 17614
rect -2172 17580 -2166 17614
rect -2212 17542 -2166 17580
rect -2212 17508 -2206 17542
rect -2172 17508 -2166 17542
rect -2212 17470 -2166 17508
rect -2212 17436 -2206 17470
rect -2172 17436 -2166 17470
rect -2212 17398 -2166 17436
rect -2212 17364 -2206 17398
rect -2172 17364 -2166 17398
rect -2212 17326 -2166 17364
rect -2212 17292 -2206 17326
rect -2172 17292 -2166 17326
rect -2212 17254 -2166 17292
rect -2212 17220 -2206 17254
rect -2172 17220 -2166 17254
rect -2212 17182 -2166 17220
rect -2212 17148 -2206 17182
rect -2172 17148 -2166 17182
rect -2212 17110 -2166 17148
rect -2212 17076 -2206 17110
rect -2172 17076 -2166 17110
rect -2212 17038 -2166 17076
rect -2212 17004 -2206 17038
rect -2172 17004 -2166 17038
rect -2212 16966 -2166 17004
rect -2212 16932 -2206 16966
rect -2172 16932 -2166 16966
rect -2212 16894 -2166 16932
rect -2212 16860 -2206 16894
rect -2172 16860 -2166 16894
rect -2212 16822 -2166 16860
rect -2212 16788 -2206 16822
rect -2172 16788 -2166 16822
rect -2212 16750 -2166 16788
rect -2212 16716 -2206 16750
rect -2172 16716 -2166 16750
rect -2212 16678 -2166 16716
rect -2212 16644 -2206 16678
rect -2172 16644 -2166 16678
rect -2212 16606 -2166 16644
rect -2212 16572 -2206 16606
rect -2172 16572 -2166 16606
rect -2212 16534 -2166 16572
rect -2212 16500 -2206 16534
rect -2172 16500 -2166 16534
rect -2212 16462 -2166 16500
rect -2212 16428 -2206 16462
rect -2172 16428 -2166 16462
rect -2212 16390 -2166 16428
rect -2430 16356 -2341 16364
rect -2471 16334 -2341 16356
rect -2471 16318 -2434 16334
rect -2471 16284 -2464 16318
rect -2471 16282 -2434 16284
rect -2382 16282 -2341 16334
rect -2471 16270 -2341 16282
rect -2471 16246 -2434 16270
rect -2471 16212 -2464 16246
rect -2382 16218 -2341 16270
rect -2430 16212 -2341 16218
rect -2471 16206 -2341 16212
rect -2471 16174 -2434 16206
rect -2471 16140 -2464 16174
rect -2382 16154 -2341 16206
rect -2430 16140 -2341 16154
rect -2471 16123 -2341 16140
rect -2212 16356 -2206 16390
rect -2172 16356 -2166 16390
rect -1954 17830 -1908 17868
rect -1954 17796 -1948 17830
rect -1914 17796 -1908 17830
rect -1954 17758 -1908 17796
rect -1954 17724 -1948 17758
rect -1914 17724 -1908 17758
rect -1954 17686 -1908 17724
rect -1954 17652 -1948 17686
rect -1914 17652 -1908 17686
rect -1954 17614 -1908 17652
rect -1954 17580 -1948 17614
rect -1914 17580 -1908 17614
rect -1954 17542 -1908 17580
rect -1954 17508 -1948 17542
rect -1914 17508 -1908 17542
rect -1954 17470 -1908 17508
rect -1954 17436 -1948 17470
rect -1914 17436 -1908 17470
rect -1954 17398 -1908 17436
rect -1954 17364 -1948 17398
rect -1914 17364 -1908 17398
rect -1954 17326 -1908 17364
rect -1954 17292 -1948 17326
rect -1914 17292 -1908 17326
rect -1954 17254 -1908 17292
rect -1954 17220 -1948 17254
rect -1914 17220 -1908 17254
rect -1954 17182 -1908 17220
rect -1954 17148 -1948 17182
rect -1914 17148 -1908 17182
rect -1954 17110 -1908 17148
rect -1954 17076 -1948 17110
rect -1914 17076 -1908 17110
rect -1954 17038 -1908 17076
rect -1954 17004 -1948 17038
rect -1914 17004 -1908 17038
rect -1954 16966 -1908 17004
rect -1954 16932 -1948 16966
rect -1914 16932 -1908 16966
rect -1954 16894 -1908 16932
rect -1954 16860 -1948 16894
rect -1914 16860 -1908 16894
rect -1954 16822 -1908 16860
rect -1954 16788 -1948 16822
rect -1914 16788 -1908 16822
rect -1954 16750 -1908 16788
rect -1954 16716 -1948 16750
rect -1914 16716 -1908 16750
rect -1954 16678 -1908 16716
rect -1954 16644 -1948 16678
rect -1914 16644 -1908 16678
rect -1954 16606 -1908 16644
rect -1954 16572 -1948 16606
rect -1914 16572 -1908 16606
rect -1954 16534 -1908 16572
rect -1954 16500 -1948 16534
rect -1914 16500 -1908 16534
rect -1954 16462 -1908 16500
rect -1954 16428 -1948 16462
rect -1914 16428 -1908 16462
rect -1954 16390 -1908 16428
rect -1954 16370 -1948 16390
rect -2212 16318 -2166 16356
rect -2212 16284 -2206 16318
rect -2172 16284 -2166 16318
rect -2212 16246 -2166 16284
rect -2212 16212 -2206 16246
rect -2172 16212 -2166 16246
rect -2212 16174 -2166 16212
rect -2212 16140 -2206 16174
rect -2172 16140 -2166 16174
rect -2470 16093 -2424 16123
rect -2212 16093 -2166 16140
rect -1957 16356 -1948 16370
rect -1914 16370 -1908 16390
rect -1696 18071 -1565 18093
rect -1696 18046 -1658 18071
rect -1696 18012 -1690 18046
rect -1606 18019 -1565 18071
rect -1656 18012 -1565 18019
rect -1696 18007 -1565 18012
rect -1696 17974 -1658 18007
rect -1696 17940 -1690 17974
rect -1606 17955 -1565 18007
rect -1656 17943 -1565 17955
rect -1696 17902 -1658 17940
rect -1696 17868 -1690 17902
rect -1606 17891 -1565 17943
rect -1656 17868 -1565 17891
rect -1696 17860 -1565 17868
rect -1438 18046 -1392 18093
rect -1438 18012 -1432 18046
rect -1398 18012 -1392 18046
rect -1438 17974 -1392 18012
rect -1438 17940 -1432 17974
rect -1398 17940 -1392 17974
rect -1438 17902 -1392 17940
rect -1438 17868 -1432 17902
rect -1398 17868 -1392 17902
rect -1696 17830 -1650 17860
rect -1696 17796 -1690 17830
rect -1656 17796 -1650 17830
rect -1696 17758 -1650 17796
rect -1696 17724 -1690 17758
rect -1656 17724 -1650 17758
rect -1696 17686 -1650 17724
rect -1696 17652 -1690 17686
rect -1656 17652 -1650 17686
rect -1696 17614 -1650 17652
rect -1696 17580 -1690 17614
rect -1656 17580 -1650 17614
rect -1696 17542 -1650 17580
rect -1696 17508 -1690 17542
rect -1656 17508 -1650 17542
rect -1696 17470 -1650 17508
rect -1696 17436 -1690 17470
rect -1656 17436 -1650 17470
rect -1696 17398 -1650 17436
rect -1696 17364 -1690 17398
rect -1656 17364 -1650 17398
rect -1696 17326 -1650 17364
rect -1696 17292 -1690 17326
rect -1656 17292 -1650 17326
rect -1696 17254 -1650 17292
rect -1696 17220 -1690 17254
rect -1656 17220 -1650 17254
rect -1696 17182 -1650 17220
rect -1696 17148 -1690 17182
rect -1656 17148 -1650 17182
rect -1696 17110 -1650 17148
rect -1696 17076 -1690 17110
rect -1656 17076 -1650 17110
rect -1696 17038 -1650 17076
rect -1696 17004 -1690 17038
rect -1656 17004 -1650 17038
rect -1696 16966 -1650 17004
rect -1696 16932 -1690 16966
rect -1656 16932 -1650 16966
rect -1696 16894 -1650 16932
rect -1696 16860 -1690 16894
rect -1656 16860 -1650 16894
rect -1696 16822 -1650 16860
rect -1696 16788 -1690 16822
rect -1656 16788 -1650 16822
rect -1696 16750 -1650 16788
rect -1696 16716 -1690 16750
rect -1656 16716 -1650 16750
rect -1696 16678 -1650 16716
rect -1696 16644 -1690 16678
rect -1656 16644 -1650 16678
rect -1696 16606 -1650 16644
rect -1696 16572 -1690 16606
rect -1656 16572 -1650 16606
rect -1696 16534 -1650 16572
rect -1696 16500 -1690 16534
rect -1656 16500 -1650 16534
rect -1696 16462 -1650 16500
rect -1696 16428 -1690 16462
rect -1656 16428 -1650 16462
rect -1696 16390 -1650 16428
rect -1914 16356 -1827 16370
rect -1957 16340 -1827 16356
rect -1957 16318 -1920 16340
rect -1957 16284 -1948 16318
rect -1868 16288 -1827 16340
rect -1914 16284 -1827 16288
rect -1957 16276 -1827 16284
rect -1957 16246 -1920 16276
rect -1957 16212 -1948 16246
rect -1868 16224 -1827 16276
rect -1914 16212 -1827 16224
rect -1957 16174 -1920 16212
rect -1957 16140 -1948 16174
rect -1868 16160 -1827 16212
rect -1914 16140 -1827 16160
rect -1957 16129 -1827 16140
rect -1696 16356 -1690 16390
rect -1656 16356 -1650 16390
rect -1438 17830 -1392 17868
rect -1438 17796 -1432 17830
rect -1398 17796 -1392 17830
rect -1438 17758 -1392 17796
rect -1438 17724 -1432 17758
rect -1398 17724 -1392 17758
rect -1438 17686 -1392 17724
rect -1438 17652 -1432 17686
rect -1398 17652 -1392 17686
rect -1438 17614 -1392 17652
rect -1438 17580 -1432 17614
rect -1398 17580 -1392 17614
rect -1438 17542 -1392 17580
rect -1438 17508 -1432 17542
rect -1398 17508 -1392 17542
rect -1438 17470 -1392 17508
rect -1438 17436 -1432 17470
rect -1398 17436 -1392 17470
rect -1438 17398 -1392 17436
rect -1438 17364 -1432 17398
rect -1398 17364 -1392 17398
rect -1438 17326 -1392 17364
rect -1438 17292 -1432 17326
rect -1398 17292 -1392 17326
rect -1438 17254 -1392 17292
rect -1438 17220 -1432 17254
rect -1398 17220 -1392 17254
rect -1438 17182 -1392 17220
rect -1438 17148 -1432 17182
rect -1398 17148 -1392 17182
rect -1438 17110 -1392 17148
rect -1438 17076 -1432 17110
rect -1398 17076 -1392 17110
rect -1438 17038 -1392 17076
rect -1438 17004 -1432 17038
rect -1398 17004 -1392 17038
rect -1438 16966 -1392 17004
rect -1438 16932 -1432 16966
rect -1398 16932 -1392 16966
rect -1438 16894 -1392 16932
rect -1438 16860 -1432 16894
rect -1398 16860 -1392 16894
rect -1438 16822 -1392 16860
rect -1438 16788 -1432 16822
rect -1398 16788 -1392 16822
rect -1438 16750 -1392 16788
rect -1438 16716 -1432 16750
rect -1398 16716 -1392 16750
rect -1438 16678 -1392 16716
rect -1438 16644 -1432 16678
rect -1398 16644 -1392 16678
rect -1438 16606 -1392 16644
rect -1438 16572 -1432 16606
rect -1398 16572 -1392 16606
rect -1438 16534 -1392 16572
rect -1438 16500 -1432 16534
rect -1398 16500 -1392 16534
rect -1438 16462 -1392 16500
rect -1438 16428 -1432 16462
rect -1398 16428 -1392 16462
rect -1438 16390 -1392 16428
rect -1438 16371 -1432 16390
rect -1696 16318 -1650 16356
rect -1696 16284 -1690 16318
rect -1656 16284 -1650 16318
rect -1696 16246 -1650 16284
rect -1696 16212 -1690 16246
rect -1656 16212 -1650 16246
rect -1696 16174 -1650 16212
rect -1696 16140 -1690 16174
rect -1656 16140 -1650 16174
rect -1954 16093 -1908 16129
rect -1696 16093 -1650 16140
rect -1441 16356 -1432 16371
rect -1398 16371 -1392 16390
rect -1180 18063 -1046 18093
rect -1180 18046 -1139 18063
rect -1180 18012 -1174 18046
rect -1140 18012 -1139 18046
rect -1180 18011 -1139 18012
rect -1087 18011 -1046 18063
rect -1180 17999 -1046 18011
rect -1180 17974 -1139 17999
rect -1180 17940 -1174 17974
rect -1140 17947 -1139 17974
rect -1087 17947 -1046 17999
rect -1140 17940 -1046 17947
rect -1180 17935 -1046 17940
rect -1180 17902 -1139 17935
rect -1180 17868 -1174 17902
rect -1140 17883 -1139 17902
rect -1087 17883 -1046 17935
rect -1140 17868 -1046 17883
rect -1180 17852 -1046 17868
rect -922 18046 -876 18093
rect -922 18012 -916 18046
rect -882 18012 -876 18046
rect -922 17974 -876 18012
rect -922 17940 -916 17974
rect -882 17940 -876 17974
rect -922 17902 -876 17940
rect -922 17868 -916 17902
rect -882 17868 -876 17902
rect -1180 17830 -1134 17852
rect -1180 17796 -1174 17830
rect -1140 17796 -1134 17830
rect -1180 17758 -1134 17796
rect -1180 17724 -1174 17758
rect -1140 17724 -1134 17758
rect -1180 17686 -1134 17724
rect -1180 17652 -1174 17686
rect -1140 17652 -1134 17686
rect -1180 17614 -1134 17652
rect -1180 17580 -1174 17614
rect -1140 17580 -1134 17614
rect -1180 17542 -1134 17580
rect -1180 17508 -1174 17542
rect -1140 17508 -1134 17542
rect -1180 17470 -1134 17508
rect -1180 17436 -1174 17470
rect -1140 17436 -1134 17470
rect -1180 17398 -1134 17436
rect -1180 17364 -1174 17398
rect -1140 17364 -1134 17398
rect -1180 17326 -1134 17364
rect -1180 17292 -1174 17326
rect -1140 17292 -1134 17326
rect -1180 17254 -1134 17292
rect -1180 17220 -1174 17254
rect -1140 17220 -1134 17254
rect -1180 17182 -1134 17220
rect -1180 17148 -1174 17182
rect -1140 17148 -1134 17182
rect -1180 17110 -1134 17148
rect -1180 17076 -1174 17110
rect -1140 17076 -1134 17110
rect -1180 17038 -1134 17076
rect -1180 17004 -1174 17038
rect -1140 17004 -1134 17038
rect -1180 16966 -1134 17004
rect -1180 16932 -1174 16966
rect -1140 16932 -1134 16966
rect -1180 16894 -1134 16932
rect -1180 16860 -1174 16894
rect -1140 16860 -1134 16894
rect -1180 16822 -1134 16860
rect -1180 16788 -1174 16822
rect -1140 16788 -1134 16822
rect -1180 16750 -1134 16788
rect -1180 16716 -1174 16750
rect -1140 16716 -1134 16750
rect -1180 16678 -1134 16716
rect -1180 16644 -1174 16678
rect -1140 16644 -1134 16678
rect -1180 16606 -1134 16644
rect -1180 16572 -1174 16606
rect -1140 16572 -1134 16606
rect -1180 16534 -1134 16572
rect -1180 16500 -1174 16534
rect -1140 16500 -1134 16534
rect -1180 16462 -1134 16500
rect -1180 16428 -1174 16462
rect -1140 16428 -1134 16462
rect -1180 16390 -1134 16428
rect -1398 16356 -1311 16371
rect -1441 16341 -1311 16356
rect -1441 16318 -1404 16341
rect -1441 16284 -1432 16318
rect -1352 16289 -1311 16341
rect -1398 16284 -1311 16289
rect -1441 16277 -1311 16284
rect -1441 16246 -1404 16277
rect -1441 16212 -1432 16246
rect -1352 16225 -1311 16277
rect -1398 16213 -1311 16225
rect -1441 16174 -1404 16212
rect -1441 16140 -1432 16174
rect -1352 16161 -1311 16213
rect -1398 16140 -1311 16161
rect -1441 16130 -1311 16140
rect -1180 16356 -1174 16390
rect -1140 16356 -1134 16390
rect -1180 16318 -1134 16356
rect -1180 16284 -1174 16318
rect -1140 16284 -1134 16318
rect -1180 16246 -1134 16284
rect -1180 16212 -1174 16246
rect -1140 16212 -1134 16246
rect -1180 16174 -1134 16212
rect -1180 16140 -1174 16174
rect -1140 16140 -1134 16174
rect -1438 16093 -1392 16130
rect -1180 16093 -1134 16140
rect -922 17830 -876 17868
rect -665 18067 -535 18097
rect -665 18046 -628 18067
rect -665 18012 -658 18046
rect -576 18015 -535 18067
rect -624 18012 -535 18015
rect -665 18003 -535 18012
rect -665 17974 -628 18003
rect -665 17940 -658 17974
rect -576 17951 -535 18003
rect -624 17940 -535 17951
rect -665 17939 -535 17940
rect -665 17902 -628 17939
rect -665 17868 -658 17902
rect -576 17887 -535 17939
rect -624 17868 -535 17887
rect -665 17856 -535 17868
rect -406 18046 -360 18093
rect -406 18012 -400 18046
rect -366 18012 -360 18046
rect -406 17974 -360 18012
rect -406 17940 -400 17974
rect -366 17940 -360 17974
rect -406 17902 -360 17940
rect -406 17868 -400 17902
rect -366 17868 -360 17902
rect -922 17796 -916 17830
rect -882 17796 -876 17830
rect -922 17758 -876 17796
rect -922 17724 -916 17758
rect -882 17724 -876 17758
rect -922 17686 -876 17724
rect -922 17652 -916 17686
rect -882 17652 -876 17686
rect -922 17614 -876 17652
rect -922 17580 -916 17614
rect -882 17580 -876 17614
rect -922 17542 -876 17580
rect -922 17508 -916 17542
rect -882 17508 -876 17542
rect -922 17470 -876 17508
rect -922 17436 -916 17470
rect -882 17436 -876 17470
rect -922 17398 -876 17436
rect -922 17364 -916 17398
rect -882 17364 -876 17398
rect -922 17326 -876 17364
rect -922 17292 -916 17326
rect -882 17292 -876 17326
rect -922 17254 -876 17292
rect -922 17220 -916 17254
rect -882 17220 -876 17254
rect -922 17182 -876 17220
rect -922 17148 -916 17182
rect -882 17148 -876 17182
rect -922 17110 -876 17148
rect -922 17076 -916 17110
rect -882 17076 -876 17110
rect -922 17038 -876 17076
rect -922 17004 -916 17038
rect -882 17004 -876 17038
rect -922 16966 -876 17004
rect -922 16932 -916 16966
rect -882 16932 -876 16966
rect -922 16894 -876 16932
rect -922 16860 -916 16894
rect -882 16860 -876 16894
rect -922 16822 -876 16860
rect -922 16788 -916 16822
rect -882 16788 -876 16822
rect -922 16750 -876 16788
rect -922 16716 -916 16750
rect -882 16716 -876 16750
rect -922 16678 -876 16716
rect -922 16644 -916 16678
rect -882 16644 -876 16678
rect -922 16606 -876 16644
rect -922 16572 -916 16606
rect -882 16572 -876 16606
rect -922 16534 -876 16572
rect -922 16500 -916 16534
rect -882 16500 -876 16534
rect -922 16462 -876 16500
rect -922 16428 -916 16462
rect -882 16428 -876 16462
rect -922 16390 -876 16428
rect -922 16356 -916 16390
rect -882 16374 -876 16390
rect -664 17830 -618 17856
rect -664 17796 -658 17830
rect -624 17796 -618 17830
rect -664 17758 -618 17796
rect -664 17724 -658 17758
rect -624 17724 -618 17758
rect -664 17686 -618 17724
rect -664 17652 -658 17686
rect -624 17652 -618 17686
rect -664 17614 -618 17652
rect -664 17580 -658 17614
rect -624 17580 -618 17614
rect -664 17542 -618 17580
rect -664 17508 -658 17542
rect -624 17508 -618 17542
rect -664 17470 -618 17508
rect -664 17436 -658 17470
rect -624 17436 -618 17470
rect -664 17398 -618 17436
rect -664 17364 -658 17398
rect -624 17364 -618 17398
rect -664 17326 -618 17364
rect -664 17292 -658 17326
rect -624 17292 -618 17326
rect -664 17254 -618 17292
rect -664 17220 -658 17254
rect -624 17220 -618 17254
rect -664 17182 -618 17220
rect -664 17148 -658 17182
rect -624 17148 -618 17182
rect -664 17110 -618 17148
rect -664 17076 -658 17110
rect -624 17076 -618 17110
rect -664 17038 -618 17076
rect -664 17004 -658 17038
rect -624 17004 -618 17038
rect -664 16966 -618 17004
rect -664 16932 -658 16966
rect -624 16932 -618 16966
rect -664 16894 -618 16932
rect -664 16860 -658 16894
rect -624 16860 -618 16894
rect -664 16822 -618 16860
rect -664 16788 -658 16822
rect -624 16788 -618 16822
rect -664 16750 -618 16788
rect -664 16716 -658 16750
rect -624 16716 -618 16750
rect -664 16678 -618 16716
rect -664 16644 -658 16678
rect -624 16644 -618 16678
rect -664 16606 -618 16644
rect -664 16572 -658 16606
rect -624 16572 -618 16606
rect -664 16534 -618 16572
rect -664 16500 -658 16534
rect -624 16500 -618 16534
rect -664 16462 -618 16500
rect -664 16428 -658 16462
rect -624 16428 -618 16462
rect -664 16390 -618 16428
rect -882 16356 -789 16374
rect -922 16344 -789 16356
rect -922 16318 -882 16344
rect -922 16284 -916 16318
rect -830 16292 -789 16344
rect -882 16284 -789 16292
rect -922 16280 -789 16284
rect -922 16246 -882 16280
rect -922 16212 -916 16246
rect -830 16228 -789 16280
rect -882 16216 -789 16228
rect -922 16174 -882 16212
rect -922 16140 -916 16174
rect -830 16164 -789 16216
rect -882 16140 -789 16164
rect -922 16133 -789 16140
rect -664 16356 -658 16390
rect -624 16356 -618 16390
rect -406 17830 -360 17868
rect -406 17796 -400 17830
rect -366 17796 -360 17830
rect -406 17758 -360 17796
rect -406 17724 -400 17758
rect -366 17724 -360 17758
rect 23170 18084 23216 18122
rect 23170 18050 23176 18084
rect 23210 18050 23216 18084
rect 23170 18012 23216 18050
rect 23170 17978 23176 18012
rect 23210 17978 23216 18012
rect 23170 17940 23216 17978
rect 23170 17906 23176 17940
rect 23210 17906 23216 17940
rect 23170 17868 23216 17906
rect 24228 18626 24234 18629
rect 24268 18629 24280 18660
rect 24680 18686 24692 18698
rect 24726 18698 24732 18720
rect 25744 18720 25790 18747
rect 24726 18686 24738 18698
rect 24680 18655 24738 18686
rect 24268 18626 24274 18629
rect 24228 18588 24274 18626
rect 24228 18554 24234 18588
rect 24268 18554 24274 18588
rect 24228 18516 24274 18554
rect 24228 18482 24234 18516
rect 24268 18482 24274 18516
rect 24228 18444 24274 18482
rect 24228 18410 24234 18444
rect 24268 18410 24274 18444
rect 24228 18372 24274 18410
rect 24228 18338 24234 18372
rect 24268 18338 24274 18372
rect 24228 18300 24274 18338
rect 24680 18603 24684 18655
rect 24736 18603 24738 18655
rect 24680 18591 24738 18603
rect 24680 18539 24684 18591
rect 24736 18539 24738 18591
rect 24680 18527 24738 18539
rect 24680 18475 24684 18527
rect 24736 18475 24738 18527
rect 24680 18470 24692 18475
rect 24726 18470 24738 18475
rect 24680 18463 24738 18470
rect 24680 18411 24684 18463
rect 24736 18411 24738 18463
rect 24680 18399 24692 18411
rect 24726 18399 24738 18411
rect 24680 18347 24684 18399
rect 24736 18347 24738 18399
rect 24680 18326 24692 18347
rect 24726 18326 24738 18347
rect 24680 18306 24738 18326
rect 25744 18686 25750 18720
rect 25784 18686 25790 18720
rect 26802 18720 26848 18747
rect 26802 18698 26808 18720
rect 25744 18648 25790 18686
rect 25744 18614 25750 18648
rect 25784 18614 25790 18648
rect 25744 18576 25790 18614
rect 25744 18542 25750 18576
rect 25784 18542 25790 18576
rect 25744 18504 25790 18542
rect 25744 18470 25750 18504
rect 25784 18470 25790 18504
rect 25744 18432 25790 18470
rect 25744 18398 25750 18432
rect 25784 18398 25790 18432
rect 25744 18360 25790 18398
rect 25744 18326 25750 18360
rect 25784 18326 25790 18360
rect 24228 18266 24234 18300
rect 24268 18266 24274 18300
rect 24228 18228 24274 18266
rect 24228 18194 24234 18228
rect 24268 18194 24274 18228
rect 24228 18156 24274 18194
rect 24228 18122 24234 18156
rect 24268 18122 24274 18156
rect 24228 18084 24274 18122
rect 24228 18050 24234 18084
rect 24268 18050 24274 18084
rect 24228 18012 24274 18050
rect 24228 17978 24234 18012
rect 24268 17978 24274 18012
rect 24228 17940 24274 17978
rect 24228 17906 24234 17940
rect 24268 17906 24274 17940
rect 24228 17899 24274 17906
rect 24686 18288 24732 18306
rect 24686 18254 24692 18288
rect 24726 18254 24732 18288
rect 24686 18216 24732 18254
rect 24686 18182 24692 18216
rect 24726 18182 24732 18216
rect 24686 18144 24732 18182
rect 24686 18110 24692 18144
rect 24726 18110 24732 18144
rect 24686 18072 24732 18110
rect 24686 18038 24692 18072
rect 24726 18038 24732 18072
rect 24686 18000 24732 18038
rect 24686 17966 24692 18000
rect 24726 17966 24732 18000
rect 24686 17928 24732 17966
rect 23170 17834 23176 17868
rect 23210 17834 23216 17868
rect 23170 17796 23216 17834
rect 23170 17762 23176 17796
rect 23210 17762 23216 17796
rect 23170 17747 23216 17762
rect 24222 17868 24280 17899
rect 24222 17834 24234 17868
rect 24268 17834 24280 17868
rect 24222 17796 24280 17834
rect 24222 17762 24234 17796
rect 24268 17762 24280 17796
rect -406 17686 -360 17724
rect 24222 17706 24280 17762
rect -406 17652 -400 17686
rect -366 17652 -360 17686
rect -406 17614 -360 17652
rect -406 17580 -400 17614
rect -366 17580 -360 17614
rect -406 17542 -360 17580
rect -406 17508 -400 17542
rect -366 17508 -360 17542
rect 23226 17700 24280 17706
rect 23226 17666 23273 17700
rect 23307 17666 23345 17700
rect 23379 17666 23417 17700
rect 23451 17666 23489 17700
rect 23523 17666 23561 17700
rect 23595 17666 23633 17700
rect 23667 17666 23705 17700
rect 23739 17666 23777 17700
rect 23811 17666 23849 17700
rect 23883 17666 23921 17700
rect 23955 17666 23993 17700
rect 24027 17666 24065 17700
rect 24099 17666 24137 17700
rect 24171 17666 24280 17700
rect 23226 17653 24280 17666
rect 24686 17894 24692 17928
rect 24726 17894 24732 17928
rect 24686 17856 24732 17894
rect 24686 17822 24692 17856
rect 24726 17822 24732 17856
rect 24686 17784 24732 17822
rect 24686 17750 24692 17784
rect 24726 17750 24732 17784
rect 24686 17712 24732 17750
rect 24686 17678 24692 17712
rect 24726 17678 24732 17712
rect 23226 17535 24541 17653
rect -406 17470 -360 17508
rect -406 17436 -400 17470
rect -366 17436 -360 17470
rect -406 17398 -360 17436
rect -406 17364 -400 17398
rect -366 17364 -360 17398
rect -406 17326 -360 17364
rect -406 17292 -400 17326
rect -366 17292 -360 17326
rect -406 17254 -360 17292
rect -406 17220 -400 17254
rect -366 17220 -360 17254
rect -406 17182 -360 17220
rect -406 17148 -400 17182
rect -366 17148 -360 17182
rect 23200 17208 24192 17214
rect 23200 17174 23247 17208
rect 23281 17174 23319 17208
rect 23353 17174 23391 17208
rect 23425 17174 23463 17208
rect 23497 17174 23535 17208
rect 23569 17174 23607 17208
rect 23641 17174 23679 17208
rect 23713 17174 23751 17208
rect 23785 17174 23823 17208
rect 23857 17174 23895 17208
rect 23929 17174 23967 17208
rect 24001 17174 24039 17208
rect 24073 17174 24111 17208
rect 24145 17174 24192 17208
rect 23200 17168 24192 17174
rect -406 17110 -360 17148
rect -406 17076 -400 17110
rect -366 17076 -360 17110
rect -406 17038 -360 17076
rect -406 17004 -400 17038
rect -366 17004 -360 17038
rect -406 16966 -360 17004
rect -406 16932 -400 16966
rect -366 16932 -360 16966
rect -406 16894 -360 16932
rect -406 16860 -400 16894
rect -366 16860 -360 16894
rect -406 16822 -360 16860
rect -406 16788 -400 16822
rect -366 16788 -360 16822
rect -406 16750 -360 16788
rect -406 16716 -400 16750
rect -366 16716 -360 16750
rect -406 16678 -360 16716
rect -406 16644 -400 16678
rect -366 16644 -360 16678
rect -406 16606 -360 16644
rect -406 16572 -400 16606
rect -366 16572 -360 16606
rect -406 16534 -360 16572
rect -406 16500 -400 16534
rect -366 16500 -360 16534
rect -406 16462 -360 16500
rect -406 16428 -400 16462
rect -366 16428 -360 16462
rect -406 16390 -360 16428
rect -406 16368 -400 16390
rect -664 16318 -618 16356
rect -664 16284 -658 16318
rect -624 16284 -618 16318
rect -664 16246 -618 16284
rect -664 16212 -658 16246
rect -624 16212 -618 16246
rect -664 16174 -618 16212
rect -664 16140 -658 16174
rect -624 16140 -618 16174
rect -922 16093 -876 16133
rect -664 16093 -618 16140
rect -413 16356 -400 16368
rect -366 16368 -360 16390
rect 10297 17061 11322 17122
rect 10297 17054 10358 17061
rect 11256 17054 11322 17061
rect -366 16356 -283 16368
rect -413 16338 -283 16356
rect -413 16318 -376 16338
rect -413 16284 -400 16318
rect -324 16286 -283 16338
rect -366 16284 -283 16286
rect -413 16274 -283 16284
rect -413 16246 -376 16274
rect -413 16212 -400 16246
rect -324 16222 -283 16274
rect -366 16212 -283 16222
rect -413 16210 -283 16212
rect -413 16174 -376 16210
rect -413 16140 -400 16174
rect -324 16158 -283 16210
rect -366 16140 -283 16158
rect -413 16127 -283 16140
rect -15 16341 241 16377
rect -15 16161 23 16341
rect 203 16161 241 16341
rect -15 16127 241 16161
rect -406 16093 -360 16127
rect -2930 16046 -2738 16052
rect -2930 16016 -2887 16046
rect -3954 16012 -2887 16016
rect -2853 16012 -2815 16046
rect -2781 16016 -2738 16046
rect -2672 16046 -2480 16052
rect -2672 16016 -2629 16046
rect -2781 16012 -2629 16016
rect -2595 16012 -2557 16046
rect -2523 16016 -2480 16046
rect -2414 16046 -2222 16052
rect -2414 16016 -2371 16046
rect -2523 16012 -2371 16016
rect -2337 16012 -2299 16046
rect -2265 16016 -2222 16046
rect -2156 16046 -1964 16052
rect -2156 16016 -2113 16046
rect -2265 16012 -2113 16016
rect -2079 16012 -2041 16046
rect -2007 16016 -1964 16046
rect -1898 16046 -1706 16052
rect -1898 16016 -1855 16046
rect -2007 16012 -1855 16016
rect -1821 16012 -1783 16046
rect -1749 16016 -1706 16046
rect -1640 16046 -1448 16052
rect -1640 16016 -1597 16046
rect -1749 16012 -1597 16016
rect -1563 16012 -1525 16046
rect -1491 16016 -1448 16046
rect -1382 16046 -1190 16052
rect -1382 16016 -1339 16046
rect -1491 16012 -1339 16016
rect -1305 16012 -1267 16046
rect -1233 16016 -1190 16046
rect -1124 16046 -932 16052
rect -1124 16016 -1081 16046
rect -1233 16012 -1081 16016
rect -1047 16012 -1009 16046
rect -975 16016 -932 16046
rect -866 16046 -674 16052
rect -866 16016 -823 16046
rect -975 16012 -823 16016
rect -789 16012 -751 16046
rect -717 16016 -674 16046
rect -608 16046 -416 16052
rect -608 16016 -565 16046
rect -717 16012 -565 16016
rect -531 16012 -493 16046
rect -459 16016 -416 16046
rect -459 16012 -404 16016
rect -3954 15936 -404 16012
rect -6095 15212 -5697 15213
rect -5120 15212 -4068 15218
rect -7593 15200 -4068 15212
rect -7593 15171 -4214 15200
rect -7593 15163 -5006 15171
rect -7593 15057 -7075 15163
rect -6825 15162 -5006 15163
rect -6825 15057 -6059 15162
rect -7593 15056 -6059 15057
rect -5737 15137 -5006 15162
rect -4972 15137 -4214 15171
rect -5737 15099 -4214 15137
rect -5737 15065 -5006 15099
rect -4972 15065 -4214 15099
rect -5737 15056 -4214 15065
rect -7593 15020 -4214 15056
rect -4098 15020 -4068 15200
rect -7593 15002 -4068 15020
rect -7593 14997 -4913 15002
rect -7138 14903 -6714 14997
rect -7138 14902 -6715 14903
rect -6095 14875 -5697 14997
rect -5466 14944 -5226 14964
rect -5466 14892 -5437 14944
rect -5385 14892 -5373 14944
rect -5321 14892 -5309 14944
rect -5257 14892 -5226 14944
rect -5061 14909 -4913 14997
rect -5466 14874 -5226 14892
rect -3949 14885 -3776 15936
rect 10297 15018 10333 17054
rect 11281 15018 11322 17054
rect 23144 17121 23190 17136
rect 23144 17087 23150 17121
rect 23184 17087 23190 17121
rect 24202 17121 24248 17136
rect 24202 17106 24208 17121
rect 23144 17049 23190 17087
rect 23144 17015 23150 17049
rect 23184 17015 23190 17049
rect 23144 16977 23190 17015
rect 23144 16943 23150 16977
rect 23184 16943 23190 16977
rect 24196 17087 24208 17106
rect 24242 17106 24248 17121
rect 24395 17106 24541 17535
rect 24686 17640 24732 17678
rect 24686 17606 24692 17640
rect 24726 17606 24732 17640
rect 24686 17568 24732 17606
rect 25744 18288 25790 18326
rect 26796 18686 26808 18698
rect 26842 18698 26848 18720
rect 27860 18720 27906 18747
rect 26842 18686 26854 18698
rect 26796 18659 26854 18686
rect 26796 18607 26798 18659
rect 26850 18607 26854 18659
rect 26796 18595 26854 18607
rect 26796 18543 26798 18595
rect 26850 18543 26854 18595
rect 26796 18542 26808 18543
rect 26842 18542 26854 18543
rect 26796 18531 26854 18542
rect 26796 18479 26798 18531
rect 26850 18479 26854 18531
rect 26796 18470 26808 18479
rect 26842 18470 26854 18479
rect 26796 18467 26854 18470
rect 26796 18415 26798 18467
rect 26850 18415 26854 18467
rect 26796 18403 26808 18415
rect 26842 18403 26854 18415
rect 26796 18351 26798 18403
rect 26850 18351 26854 18403
rect 26796 18326 26808 18351
rect 26842 18326 26854 18351
rect 26796 18306 26854 18326
rect 27860 18686 27866 18720
rect 27900 18686 27906 18720
rect 27860 18648 27906 18686
rect 27860 18614 27866 18648
rect 27900 18614 27906 18648
rect 27860 18576 27906 18614
rect 27860 18542 27866 18576
rect 27900 18542 27906 18576
rect 27860 18504 27906 18542
rect 27860 18470 27866 18504
rect 27900 18470 27906 18504
rect 27860 18432 27906 18470
rect 27860 18398 27866 18432
rect 27900 18398 27906 18432
rect 27860 18360 27906 18398
rect 27860 18326 27866 18360
rect 27900 18326 27906 18360
rect 42606 18724 42652 18762
rect 42606 18690 42612 18724
rect 42646 18690 42652 18724
rect 42606 18652 42652 18690
rect 42606 18618 42612 18652
rect 42646 18618 42652 18652
rect 42606 18580 42652 18618
rect 42606 18546 42612 18580
rect 42646 18546 42652 18580
rect 42606 18508 42652 18546
rect 42606 18474 42612 18508
rect 42646 18474 42652 18508
rect 42606 18436 42652 18474
rect 42606 18402 42612 18436
rect 42646 18402 42652 18436
rect 42606 18364 42652 18402
rect 25744 18254 25750 18288
rect 25784 18254 25790 18288
rect 25744 18216 25790 18254
rect 25744 18182 25750 18216
rect 25784 18182 25790 18216
rect 25744 18144 25790 18182
rect 25744 18110 25750 18144
rect 25784 18110 25790 18144
rect 25744 18072 25790 18110
rect 25744 18038 25750 18072
rect 25784 18038 25790 18072
rect 25744 18000 25790 18038
rect 25744 17966 25750 18000
rect 25784 17966 25790 18000
rect 25744 17928 25790 17966
rect 25744 17894 25750 17928
rect 25784 17894 25790 17928
rect 25744 17856 25790 17894
rect 25744 17822 25750 17856
rect 25784 17822 25790 17856
rect 25744 17784 25790 17822
rect 25744 17750 25750 17784
rect 25784 17750 25790 17784
rect 25744 17712 25790 17750
rect 25744 17678 25750 17712
rect 25784 17678 25790 17712
rect 25744 17640 25790 17678
rect 25744 17606 25750 17640
rect 25784 17606 25790 17640
rect 25744 17596 25790 17606
rect 26802 18288 26848 18306
rect 26802 18254 26808 18288
rect 26842 18254 26848 18288
rect 26802 18216 26848 18254
rect 26802 18182 26808 18216
rect 26842 18182 26848 18216
rect 26802 18144 26848 18182
rect 26802 18110 26808 18144
rect 26842 18110 26848 18144
rect 26802 18072 26848 18110
rect 26802 18038 26808 18072
rect 26842 18038 26848 18072
rect 26802 18000 26848 18038
rect 26802 17966 26808 18000
rect 26842 17966 26848 18000
rect 26802 17928 26848 17966
rect 26802 17894 26808 17928
rect 26842 17894 26848 17928
rect 26802 17856 26848 17894
rect 26802 17822 26808 17856
rect 26842 17822 26848 17856
rect 26802 17784 26848 17822
rect 26802 17750 26808 17784
rect 26842 17750 26848 17784
rect 26802 17712 26848 17750
rect 26802 17678 26808 17712
rect 26842 17678 26848 17712
rect 26802 17640 26848 17678
rect 26802 17606 26808 17640
rect 26842 17606 26848 17640
rect 24686 17534 24692 17568
rect 24726 17534 24732 17568
rect 24686 17496 24732 17534
rect 24686 17462 24692 17496
rect 24726 17462 24732 17496
rect 24686 17424 24732 17462
rect 24686 17390 24692 17424
rect 24726 17390 24732 17424
rect 24686 17352 24732 17390
rect 24686 17318 24692 17352
rect 24726 17318 24732 17352
rect 24686 17280 24732 17318
rect 24686 17246 24692 17280
rect 24726 17246 24732 17280
rect 24686 17208 24732 17246
rect 25738 17568 25796 17596
rect 25738 17557 25750 17568
rect 25784 17557 25796 17568
rect 25738 17505 25741 17557
rect 25793 17505 25796 17557
rect 25738 17496 25796 17505
rect 25738 17493 25750 17496
rect 25784 17493 25796 17496
rect 25738 17441 25741 17493
rect 25793 17441 25796 17493
rect 25738 17429 25796 17441
rect 25738 17377 25741 17429
rect 25793 17377 25796 17429
rect 25738 17365 25796 17377
rect 25738 17313 25741 17365
rect 25793 17313 25796 17365
rect 25738 17301 25796 17313
rect 25738 17249 25741 17301
rect 25793 17249 25796 17301
rect 25738 17246 25750 17249
rect 25784 17246 25796 17249
rect 25738 17208 25796 17246
rect 26802 17568 26848 17606
rect 27860 18288 27906 18326
rect 27860 18254 27866 18288
rect 27900 18254 27906 18288
rect 27860 18216 27906 18254
rect 27860 18182 27866 18216
rect 27900 18182 27906 18216
rect 39316 18300 39496 18344
rect 39316 18248 39348 18300
rect 39400 18248 39412 18300
rect 39464 18248 39496 18300
rect 39316 18204 39496 18248
rect 42606 18330 42612 18364
rect 42646 18330 42652 18364
rect 42606 18292 42652 18330
rect 42606 18258 42612 18292
rect 42646 18258 42652 18292
rect 42606 18220 42652 18258
rect 27860 18144 27906 18182
rect 27860 18110 27866 18144
rect 27900 18110 27906 18144
rect 27860 18072 27906 18110
rect 27860 18038 27866 18072
rect 27900 18038 27906 18072
rect 42606 18186 42612 18220
rect 42646 18186 42652 18220
rect 42606 18148 42652 18186
rect 42606 18114 42612 18148
rect 42646 18114 42652 18148
rect 42606 18076 42652 18114
rect 27860 18000 27906 18038
rect 39194 18055 39386 18061
rect 39194 18021 39237 18055
rect 39271 18021 39309 18055
rect 39343 18021 39386 18055
rect 39194 18015 39386 18021
rect 39452 18055 39644 18061
rect 39452 18021 39495 18055
rect 39529 18021 39567 18055
rect 39601 18021 39644 18055
rect 39452 18015 39644 18021
rect 42606 18042 42612 18076
rect 42646 18042 42652 18076
rect 27860 17966 27866 18000
rect 27900 17966 27906 18000
rect 42606 18004 42652 18042
rect 27860 17928 27906 17966
rect 27860 17894 27866 17928
rect 27900 17894 27906 17928
rect 27860 17856 27906 17894
rect 27860 17822 27866 17856
rect 27900 17822 27906 17856
rect 27860 17784 27906 17822
rect 27860 17750 27866 17784
rect 27900 17750 27906 17784
rect 27860 17712 27906 17750
rect 27860 17678 27866 17712
rect 27900 17678 27906 17712
rect 27860 17640 27906 17678
rect 27860 17606 27866 17640
rect 27900 17606 27906 17640
rect 27860 17596 27906 17606
rect 39138 17959 39184 17974
rect 39396 17964 39442 17974
rect 39138 17925 39144 17959
rect 39178 17925 39184 17959
rect 39138 17887 39184 17925
rect 39138 17853 39144 17887
rect 39178 17853 39184 17887
rect 39138 17815 39184 17853
rect 39346 17959 39476 17964
rect 39346 17925 39402 17959
rect 39436 17925 39476 17959
rect 39346 17873 39385 17925
rect 39437 17873 39476 17925
rect 39346 17853 39402 17873
rect 39436 17853 39476 17873
rect 39346 17834 39476 17853
rect 39654 17959 39700 17974
rect 39654 17925 39660 17959
rect 39694 17925 39700 17959
rect 39654 17887 39700 17925
rect 39654 17853 39660 17887
rect 39694 17853 39700 17887
rect 39138 17781 39144 17815
rect 39178 17781 39184 17815
rect 39138 17743 39184 17781
rect 39138 17709 39144 17743
rect 39178 17709 39184 17743
rect 39138 17671 39184 17709
rect 39138 17637 39144 17671
rect 39178 17637 39184 17671
rect 39138 17599 39184 17637
rect 26802 17534 26808 17568
rect 26842 17534 26848 17568
rect 26802 17496 26848 17534
rect 26802 17462 26808 17496
rect 26842 17462 26848 17496
rect 26802 17424 26848 17462
rect 26802 17390 26808 17424
rect 26842 17390 26848 17424
rect 26802 17352 26848 17390
rect 26802 17318 26808 17352
rect 26842 17318 26848 17352
rect 26802 17280 26848 17318
rect 26802 17246 26808 17280
rect 26842 17246 26848 17280
rect 26802 17208 26848 17246
rect 24686 17174 24692 17208
rect 24726 17174 24732 17208
rect 24686 17147 24732 17174
rect 25744 17174 25750 17208
rect 25784 17174 25790 17208
rect 25744 17147 25790 17174
rect 26802 17174 26808 17208
rect 26842 17174 26848 17208
rect 26802 17147 26848 17174
rect 27848 17568 28082 17596
rect 27848 17555 27866 17568
rect 27900 17555 28082 17568
rect 27848 17503 27855 17555
rect 27907 17503 28082 17555
rect 27848 17496 28082 17503
rect 27848 17491 27866 17496
rect 27900 17491 28082 17496
rect 27848 17439 27855 17491
rect 27907 17439 28082 17491
rect 27848 17427 28082 17439
rect 27848 17375 27855 17427
rect 27907 17375 28082 17427
rect 27848 17363 28082 17375
rect 27848 17311 27855 17363
rect 27907 17311 28082 17363
rect 27848 17299 28082 17311
rect 27848 17247 27855 17299
rect 27907 17247 28082 17299
rect 27848 17246 27866 17247
rect 27900 17246 28082 17247
rect 27848 17208 28082 17246
rect 27848 17174 27866 17208
rect 27900 17174 28082 17208
rect 27848 17147 28082 17174
rect 24242 17100 25734 17106
rect 24242 17087 24789 17100
rect 24196 17066 24789 17087
rect 24823 17066 24861 17100
rect 24895 17066 24933 17100
rect 24967 17066 25005 17100
rect 25039 17066 25077 17100
rect 25111 17066 25149 17100
rect 25183 17066 25221 17100
rect 25255 17066 25293 17100
rect 25327 17066 25365 17100
rect 25399 17066 25437 17100
rect 25471 17066 25509 17100
rect 25543 17066 25581 17100
rect 25615 17066 25653 17100
rect 25687 17066 25734 17100
rect 24196 17050 25734 17066
rect 25800 17100 26792 17106
rect 25800 17066 25847 17100
rect 25881 17066 25919 17100
rect 25953 17066 25991 17100
rect 26025 17066 26063 17100
rect 26097 17066 26135 17100
rect 26169 17066 26207 17100
rect 26241 17066 26279 17100
rect 26313 17066 26351 17100
rect 26385 17066 26423 17100
rect 26457 17066 26495 17100
rect 26529 17066 26567 17100
rect 26601 17066 26639 17100
rect 26673 17066 26711 17100
rect 26745 17066 26792 17100
rect 25800 17050 26792 17066
rect 26858 17100 27850 17106
rect 26858 17066 26905 17100
rect 26939 17066 26977 17100
rect 27011 17066 27049 17100
rect 27083 17066 27121 17100
rect 27155 17066 27193 17100
rect 27227 17066 27265 17100
rect 27299 17066 27337 17100
rect 27371 17066 27409 17100
rect 27443 17066 27481 17100
rect 27515 17066 27553 17100
rect 27587 17066 27625 17100
rect 27659 17066 27697 17100
rect 27731 17066 27769 17100
rect 27803 17066 27850 17100
rect 26858 17060 27850 17066
rect 26858 17050 27838 17060
rect 24196 17049 27838 17050
rect 24196 17015 24208 17049
rect 24242 17015 27838 17049
rect 24196 16978 27838 17015
rect 24196 16977 24832 16978
rect 24196 16948 24208 16977
rect 23144 16905 23190 16943
rect 23144 16871 23150 16905
rect 23184 16871 23190 16905
rect 23144 16833 23190 16871
rect 23144 16799 23150 16833
rect 23184 16799 23190 16833
rect 23144 16761 23190 16799
rect 23144 16727 23150 16761
rect 23184 16727 23190 16761
rect 23144 16689 23190 16727
rect 23144 16655 23150 16689
rect 23184 16655 23190 16689
rect 23144 16617 23190 16655
rect 23144 16583 23150 16617
rect 23184 16583 23190 16617
rect 23144 16545 23190 16583
rect 23144 16511 23150 16545
rect 23184 16511 23190 16545
rect 23144 16473 23190 16511
rect 23144 16439 23150 16473
rect 23184 16439 23190 16473
rect 23144 16401 23190 16439
rect 23144 16367 23150 16401
rect 23184 16367 23190 16401
rect 23144 16329 23190 16367
rect 23144 16295 23150 16329
rect 23184 16295 23190 16329
rect 23144 16257 23190 16295
rect 23144 16223 23150 16257
rect 23184 16223 23190 16257
rect 23144 16185 23190 16223
rect 22522 16117 22962 16152
rect 23144 16151 23150 16185
rect 23184 16151 23190 16185
rect 23144 16136 23190 16151
rect 24202 16943 24208 16948
rect 24242 16948 24832 16977
rect 24242 16943 24248 16948
rect 24202 16905 24248 16943
rect 24202 16871 24208 16905
rect 24242 16871 24248 16905
rect 24202 16833 24248 16871
rect 24202 16799 24208 16833
rect 24242 16799 24248 16833
rect 24202 16761 24248 16799
rect 24202 16727 24208 16761
rect 24242 16727 24248 16761
rect 24202 16689 24248 16727
rect 24202 16655 24208 16689
rect 24242 16655 24248 16689
rect 24202 16617 24248 16655
rect 24202 16583 24208 16617
rect 24242 16583 24248 16617
rect 27908 16812 28082 17147
rect 39138 17565 39144 17599
rect 39178 17565 39184 17599
rect 39138 17527 39184 17565
rect 39138 17493 39144 17527
rect 39178 17493 39184 17527
rect 39138 17455 39184 17493
rect 39138 17421 39144 17455
rect 39178 17421 39184 17455
rect 39138 17383 39184 17421
rect 39138 17349 39144 17383
rect 39178 17349 39184 17383
rect 39138 17311 39184 17349
rect 39138 17277 39144 17311
rect 39178 17277 39184 17311
rect 39138 17239 39184 17277
rect 39138 17205 39144 17239
rect 39178 17205 39184 17239
rect 39138 17167 39184 17205
rect 39138 17133 39144 17167
rect 39178 17133 39184 17167
rect 39138 17095 39184 17133
rect 39138 17061 39144 17095
rect 39178 17061 39184 17095
rect 39138 17023 39184 17061
rect 39138 17004 39144 17023
rect 39136 16989 39144 17004
rect 39178 17004 39184 17023
rect 39396 17815 39442 17834
rect 39396 17781 39402 17815
rect 39436 17781 39442 17815
rect 39396 17743 39442 17781
rect 39396 17709 39402 17743
rect 39436 17709 39442 17743
rect 39396 17671 39442 17709
rect 39396 17637 39402 17671
rect 39436 17637 39442 17671
rect 39396 17599 39442 17637
rect 39396 17565 39402 17599
rect 39436 17565 39442 17599
rect 39396 17527 39442 17565
rect 39396 17493 39402 17527
rect 39436 17493 39442 17527
rect 39396 17455 39442 17493
rect 39396 17421 39402 17455
rect 39436 17421 39442 17455
rect 39396 17383 39442 17421
rect 39396 17349 39402 17383
rect 39436 17349 39442 17383
rect 39396 17311 39442 17349
rect 39396 17277 39402 17311
rect 39436 17277 39442 17311
rect 39396 17239 39442 17277
rect 39396 17205 39402 17239
rect 39436 17205 39442 17239
rect 39396 17167 39442 17205
rect 39396 17133 39402 17167
rect 39436 17133 39442 17167
rect 39396 17095 39442 17133
rect 39396 17061 39402 17095
rect 39436 17061 39442 17095
rect 39396 17023 39442 17061
rect 39178 16989 39196 17004
rect 39136 16934 39196 16989
rect 39396 16989 39402 17023
rect 39436 16989 39442 17023
rect 39396 16974 39442 16989
rect 39654 17815 39700 17853
rect 39654 17781 39660 17815
rect 39694 17781 39700 17815
rect 39654 17743 39700 17781
rect 39654 17709 39660 17743
rect 39694 17709 39700 17743
rect 39654 17671 39700 17709
rect 39654 17637 39660 17671
rect 39694 17637 39700 17671
rect 39654 17599 39700 17637
rect 39654 17565 39660 17599
rect 39694 17565 39700 17599
rect 39654 17527 39700 17565
rect 39654 17493 39660 17527
rect 39694 17493 39700 17527
rect 39654 17455 39700 17493
rect 39654 17421 39660 17455
rect 39694 17421 39700 17455
rect 39654 17383 39700 17421
rect 39654 17349 39660 17383
rect 39694 17349 39700 17383
rect 39654 17311 39700 17349
rect 39654 17277 39660 17311
rect 39694 17277 39700 17311
rect 39654 17239 39700 17277
rect 39654 17205 39660 17239
rect 39694 17205 39700 17239
rect 39654 17167 39700 17205
rect 39654 17133 39660 17167
rect 39694 17144 39700 17167
rect 42606 17970 42612 18004
rect 42646 17970 42652 18004
rect 42606 17932 42652 17970
rect 42606 17898 42612 17932
rect 42646 17898 42652 17932
rect 42606 17860 42652 17898
rect 42606 17826 42612 17860
rect 42646 17826 42652 17860
rect 42606 17788 42652 17826
rect 42606 17754 42612 17788
rect 42646 17754 42652 17788
rect 42606 17716 42652 17754
rect 42606 17682 42612 17716
rect 42646 17682 42652 17716
rect 42606 17644 42652 17682
rect 42606 17610 42612 17644
rect 42646 17610 42652 17644
rect 42606 17572 42652 17610
rect 42606 17538 42612 17572
rect 42646 17538 42652 17572
rect 42606 17500 42652 17538
rect 42606 17466 42612 17500
rect 42646 17466 42652 17500
rect 42606 17428 42652 17466
rect 42606 17394 42612 17428
rect 42646 17394 42652 17428
rect 42606 17356 42652 17394
rect 42606 17322 42612 17356
rect 42646 17322 42652 17356
rect 42606 17284 42652 17322
rect 42606 17250 42612 17284
rect 42646 17250 42652 17284
rect 42606 17212 42652 17250
rect 42606 17178 42612 17212
rect 42646 17178 42652 17212
rect 39694 17143 39966 17144
rect 39694 17133 41816 17143
rect 39654 17117 41816 17133
rect 39654 17095 39726 17117
rect 39654 17061 39660 17095
rect 39694 17061 39726 17095
rect 39654 17023 39726 17061
rect 39654 16989 39660 17023
rect 39694 17001 39726 17023
rect 39906 17001 41816 17117
rect 39694 16989 41816 17001
rect 39654 16974 41816 16989
rect 39665 16970 41816 16974
rect 39136 16927 39646 16934
rect 39136 16893 39237 16927
rect 39271 16893 39309 16927
rect 39343 16893 39495 16927
rect 39529 16893 39567 16927
rect 39601 16893 39646 16927
rect 39136 16884 39646 16893
rect 24202 16545 24248 16583
rect 24596 16602 25017 16610
rect 24596 16568 24609 16602
rect 24643 16568 24681 16602
rect 24715 16568 24753 16602
rect 24787 16568 24825 16602
rect 24859 16568 24897 16602
rect 24931 16568 24969 16602
rect 25003 16568 25017 16602
rect 24596 16560 25017 16568
rect 27127 16602 27548 16610
rect 27127 16568 27140 16602
rect 27174 16568 27212 16602
rect 27246 16568 27284 16602
rect 27318 16568 27356 16602
rect 27390 16568 27428 16602
rect 27462 16568 27500 16602
rect 27534 16568 27548 16602
rect 27127 16560 27548 16568
rect 24202 16511 24208 16545
rect 24242 16511 24248 16545
rect 24202 16473 24248 16511
rect 24202 16439 24208 16473
rect 24242 16439 24248 16473
rect 24202 16401 24248 16439
rect 24202 16367 24208 16401
rect 24242 16367 24248 16401
rect 24202 16329 24248 16367
rect 24202 16295 24208 16329
rect 24242 16295 24248 16329
rect 27908 16315 27939 16812
rect 24202 16257 24248 16295
rect 24202 16223 24208 16257
rect 24242 16223 24248 16257
rect 24202 16185 24248 16223
rect 24202 16151 24208 16185
rect 24242 16151 24248 16185
rect 24202 16136 24248 16151
rect 24590 16284 25023 16303
rect 24590 16250 24609 16284
rect 24643 16250 24681 16284
rect 24715 16250 24753 16284
rect 24787 16250 24825 16284
rect 24859 16250 24897 16284
rect 24931 16250 24969 16284
rect 25003 16250 25023 16284
rect 22522 15745 22553 16117
rect 22925 16104 22962 16117
rect 22925 16098 24192 16104
rect 22925 16064 23247 16098
rect 23281 16064 23319 16098
rect 23353 16064 23391 16098
rect 23425 16064 23463 16098
rect 23497 16064 23535 16098
rect 23569 16064 23607 16098
rect 23641 16064 23679 16098
rect 23713 16064 23751 16098
rect 23785 16064 23823 16098
rect 23857 16064 23895 16098
rect 23929 16064 23967 16098
rect 24001 16064 24039 16098
rect 24073 16064 24111 16098
rect 24145 16064 24192 16098
rect 22925 16058 24192 16064
rect 22925 15745 22962 16058
rect 24590 15966 25023 16250
rect 27122 16284 27939 16315
rect 27122 16250 27140 16284
rect 27174 16250 27212 16284
rect 27246 16250 27284 16284
rect 27318 16250 27356 16284
rect 27390 16250 27428 16284
rect 27462 16250 27500 16284
rect 27534 16250 27939 16284
rect 27122 16248 27939 16250
rect 28055 16248 28082 16812
rect 39156 16855 39396 16884
rect 39156 16803 39223 16855
rect 39275 16803 39287 16855
rect 39339 16803 39396 16855
rect 39156 16784 39396 16803
rect 41643 16766 41816 16970
rect 42606 17140 42652 17178
rect 42606 17106 42612 17140
rect 42646 17118 42652 17140
rect 42864 18825 43003 18843
rect 42864 18796 42910 18825
rect 42864 18762 42870 18796
rect 42904 18773 42910 18796
rect 42962 18773 43003 18825
rect 42904 18762 43003 18773
rect 42864 18761 43003 18762
rect 42864 18724 42910 18761
rect 42864 18690 42870 18724
rect 42904 18709 42910 18724
rect 42962 18709 43003 18761
rect 42904 18697 43003 18709
rect 42904 18690 42910 18697
rect 42864 18652 42910 18690
rect 42864 18618 42870 18652
rect 42904 18645 42910 18652
rect 42962 18645 43003 18697
rect 42904 18618 43003 18645
rect 42864 18614 43003 18618
rect 43122 18796 43168 18843
rect 43122 18762 43128 18796
rect 43162 18762 43168 18796
rect 43122 18724 43168 18762
rect 43122 18690 43128 18724
rect 43162 18690 43168 18724
rect 43122 18652 43168 18690
rect 43122 18618 43128 18652
rect 43162 18618 43168 18652
rect 42864 18580 42910 18614
rect 42864 18546 42870 18580
rect 42904 18546 42910 18580
rect 42864 18508 42910 18546
rect 42864 18474 42870 18508
rect 42904 18474 42910 18508
rect 42864 18436 42910 18474
rect 42864 18402 42870 18436
rect 42904 18402 42910 18436
rect 42864 18364 42910 18402
rect 42864 18330 42870 18364
rect 42904 18330 42910 18364
rect 42864 18292 42910 18330
rect 42864 18258 42870 18292
rect 42904 18258 42910 18292
rect 42864 18220 42910 18258
rect 42864 18186 42870 18220
rect 42904 18186 42910 18220
rect 42864 18148 42910 18186
rect 42864 18114 42870 18148
rect 42904 18114 42910 18148
rect 42864 18076 42910 18114
rect 42864 18042 42870 18076
rect 42904 18042 42910 18076
rect 42864 18004 42910 18042
rect 42864 17970 42870 18004
rect 42904 17970 42910 18004
rect 42864 17932 42910 17970
rect 42864 17898 42870 17932
rect 42904 17898 42910 17932
rect 42864 17860 42910 17898
rect 42864 17826 42870 17860
rect 42904 17826 42910 17860
rect 42864 17788 42910 17826
rect 42864 17754 42870 17788
rect 42904 17754 42910 17788
rect 42864 17716 42910 17754
rect 42864 17682 42870 17716
rect 42904 17682 42910 17716
rect 42864 17644 42910 17682
rect 42864 17610 42870 17644
rect 42904 17610 42910 17644
rect 42864 17572 42910 17610
rect 42864 17538 42870 17572
rect 42904 17538 42910 17572
rect 42864 17500 42910 17538
rect 42864 17466 42870 17500
rect 42904 17466 42910 17500
rect 42864 17428 42910 17466
rect 42864 17394 42870 17428
rect 42904 17394 42910 17428
rect 42864 17356 42910 17394
rect 42864 17322 42870 17356
rect 42904 17322 42910 17356
rect 42864 17284 42910 17322
rect 42864 17250 42870 17284
rect 42904 17250 42910 17284
rect 42864 17212 42910 17250
rect 42864 17178 42870 17212
rect 42904 17178 42910 17212
rect 42864 17140 42910 17178
rect 42646 17106 42751 17118
rect 42606 17088 42751 17106
rect 42606 17068 42658 17088
rect 42606 17034 42612 17068
rect 42646 17036 42658 17068
rect 42710 17036 42751 17088
rect 42646 17034 42751 17036
rect 42606 17024 42751 17034
rect 42606 16996 42658 17024
rect 42606 16962 42612 16996
rect 42646 16972 42658 16996
rect 42710 16972 42751 17024
rect 42646 16962 42751 16972
rect 42606 16960 42751 16962
rect 42606 16924 42658 16960
rect 42606 16890 42612 16924
rect 42646 16908 42658 16924
rect 42710 16908 42751 16960
rect 42646 16890 42751 16908
rect 42606 16877 42751 16890
rect 42864 17106 42870 17140
rect 42904 17106 42910 17140
rect 43122 18580 43168 18618
rect 43122 18546 43128 18580
rect 43162 18546 43168 18580
rect 43122 18508 43168 18546
rect 43122 18474 43128 18508
rect 43162 18474 43168 18508
rect 43122 18436 43168 18474
rect 43122 18402 43128 18436
rect 43162 18402 43168 18436
rect 43122 18364 43168 18402
rect 43122 18330 43128 18364
rect 43162 18330 43168 18364
rect 43122 18292 43168 18330
rect 43122 18258 43128 18292
rect 43162 18258 43168 18292
rect 43122 18220 43168 18258
rect 43122 18186 43128 18220
rect 43162 18186 43168 18220
rect 43122 18148 43168 18186
rect 43122 18114 43128 18148
rect 43162 18114 43168 18148
rect 43122 18076 43168 18114
rect 43122 18042 43128 18076
rect 43162 18042 43168 18076
rect 43122 18004 43168 18042
rect 43122 17970 43128 18004
rect 43162 17970 43168 18004
rect 43122 17932 43168 17970
rect 43122 17898 43128 17932
rect 43162 17898 43168 17932
rect 43122 17860 43168 17898
rect 43122 17826 43128 17860
rect 43162 17826 43168 17860
rect 43122 17788 43168 17826
rect 43122 17754 43128 17788
rect 43162 17754 43168 17788
rect 43122 17716 43168 17754
rect 43122 17682 43128 17716
rect 43162 17682 43168 17716
rect 43122 17644 43168 17682
rect 43122 17610 43128 17644
rect 43162 17610 43168 17644
rect 43122 17572 43168 17610
rect 43122 17538 43128 17572
rect 43162 17538 43168 17572
rect 43122 17500 43168 17538
rect 43122 17466 43128 17500
rect 43162 17466 43168 17500
rect 43122 17428 43168 17466
rect 43122 17394 43128 17428
rect 43162 17394 43168 17428
rect 43122 17356 43168 17394
rect 43122 17322 43128 17356
rect 43162 17322 43168 17356
rect 43122 17284 43168 17322
rect 43122 17250 43128 17284
rect 43162 17250 43168 17284
rect 43122 17212 43168 17250
rect 43122 17178 43128 17212
rect 43162 17178 43168 17212
rect 43122 17140 43168 17178
rect 43122 17114 43128 17140
rect 42864 17068 42910 17106
rect 42864 17034 42870 17068
rect 42904 17034 42910 17068
rect 42864 16996 42910 17034
rect 42864 16962 42870 16996
rect 42904 16962 42910 16996
rect 42864 16924 42910 16962
rect 42864 16890 42870 16924
rect 42904 16890 42910 16924
rect 42606 16843 42652 16877
rect 42864 16843 42910 16890
rect 43121 17106 43128 17114
rect 43162 17114 43168 17140
rect 43380 18825 43512 18843
rect 43380 18796 43419 18825
rect 43380 18762 43386 18796
rect 43471 18773 43512 18825
rect 43420 18762 43512 18773
rect 43380 18761 43512 18762
rect 43380 18724 43419 18761
rect 43380 18690 43386 18724
rect 43471 18709 43512 18761
rect 43420 18697 43512 18709
rect 43380 18652 43419 18690
rect 43380 18618 43386 18652
rect 43471 18645 43512 18697
rect 43420 18618 43512 18645
rect 43380 18614 43512 18618
rect 43638 18796 43684 18843
rect 43638 18762 43644 18796
rect 43678 18762 43684 18796
rect 43638 18724 43684 18762
rect 43638 18690 43644 18724
rect 43678 18690 43684 18724
rect 43638 18652 43684 18690
rect 43638 18618 43644 18652
rect 43678 18618 43684 18652
rect 43380 18580 43426 18614
rect 43380 18546 43386 18580
rect 43420 18546 43426 18580
rect 43380 18508 43426 18546
rect 43380 18474 43386 18508
rect 43420 18474 43426 18508
rect 43380 18436 43426 18474
rect 43380 18402 43386 18436
rect 43420 18402 43426 18436
rect 43380 18364 43426 18402
rect 43380 18330 43386 18364
rect 43420 18330 43426 18364
rect 43380 18292 43426 18330
rect 43380 18258 43386 18292
rect 43420 18258 43426 18292
rect 43380 18220 43426 18258
rect 43380 18186 43386 18220
rect 43420 18186 43426 18220
rect 43380 18148 43426 18186
rect 43380 18114 43386 18148
rect 43420 18114 43426 18148
rect 43380 18076 43426 18114
rect 43380 18042 43386 18076
rect 43420 18042 43426 18076
rect 43380 18004 43426 18042
rect 43380 17970 43386 18004
rect 43420 17970 43426 18004
rect 43380 17932 43426 17970
rect 43380 17898 43386 17932
rect 43420 17898 43426 17932
rect 43380 17860 43426 17898
rect 43380 17826 43386 17860
rect 43420 17826 43426 17860
rect 43380 17788 43426 17826
rect 43380 17754 43386 17788
rect 43420 17754 43426 17788
rect 43380 17716 43426 17754
rect 43380 17682 43386 17716
rect 43420 17682 43426 17716
rect 43380 17644 43426 17682
rect 43380 17610 43386 17644
rect 43420 17610 43426 17644
rect 43380 17572 43426 17610
rect 43380 17538 43386 17572
rect 43420 17538 43426 17572
rect 43380 17500 43426 17538
rect 43380 17466 43386 17500
rect 43420 17466 43426 17500
rect 43380 17428 43426 17466
rect 43380 17394 43386 17428
rect 43420 17394 43426 17428
rect 43380 17356 43426 17394
rect 43380 17322 43386 17356
rect 43420 17322 43426 17356
rect 43380 17284 43426 17322
rect 43380 17250 43386 17284
rect 43420 17250 43426 17284
rect 43380 17212 43426 17250
rect 43380 17178 43386 17212
rect 43420 17178 43426 17212
rect 43380 17140 43426 17178
rect 43162 17106 43251 17114
rect 43121 17084 43251 17106
rect 43121 17068 43158 17084
rect 43121 17034 43128 17068
rect 43121 17032 43158 17034
rect 43210 17032 43251 17084
rect 43121 17020 43251 17032
rect 43121 16996 43158 17020
rect 43121 16962 43128 16996
rect 43210 16968 43251 17020
rect 43162 16962 43251 16968
rect 43121 16956 43251 16962
rect 43121 16924 43158 16956
rect 43121 16890 43128 16924
rect 43210 16904 43251 16956
rect 43162 16890 43251 16904
rect 43121 16873 43251 16890
rect 43380 17106 43386 17140
rect 43420 17106 43426 17140
rect 43638 18580 43684 18618
rect 43638 18546 43644 18580
rect 43678 18546 43684 18580
rect 43638 18508 43684 18546
rect 43638 18474 43644 18508
rect 43678 18474 43684 18508
rect 43638 18436 43684 18474
rect 43638 18402 43644 18436
rect 43678 18402 43684 18436
rect 43638 18364 43684 18402
rect 43638 18330 43644 18364
rect 43678 18330 43684 18364
rect 43638 18292 43684 18330
rect 43638 18258 43644 18292
rect 43678 18258 43684 18292
rect 43638 18220 43684 18258
rect 43638 18186 43644 18220
rect 43678 18186 43684 18220
rect 43638 18148 43684 18186
rect 43638 18114 43644 18148
rect 43678 18114 43684 18148
rect 43638 18076 43684 18114
rect 43638 18042 43644 18076
rect 43678 18042 43684 18076
rect 43638 18004 43684 18042
rect 43638 17970 43644 18004
rect 43678 17970 43684 18004
rect 43638 17932 43684 17970
rect 43638 17898 43644 17932
rect 43678 17898 43684 17932
rect 43638 17860 43684 17898
rect 43638 17826 43644 17860
rect 43678 17826 43684 17860
rect 43638 17788 43684 17826
rect 43638 17754 43644 17788
rect 43678 17754 43684 17788
rect 43638 17716 43684 17754
rect 43638 17682 43644 17716
rect 43678 17682 43684 17716
rect 43638 17644 43684 17682
rect 43638 17610 43644 17644
rect 43678 17610 43684 17644
rect 43638 17572 43684 17610
rect 43638 17538 43644 17572
rect 43678 17538 43684 17572
rect 43638 17500 43684 17538
rect 43638 17466 43644 17500
rect 43678 17466 43684 17500
rect 43638 17428 43684 17466
rect 43638 17394 43644 17428
rect 43678 17394 43684 17428
rect 43638 17356 43684 17394
rect 43638 17322 43644 17356
rect 43678 17322 43684 17356
rect 43638 17284 43684 17322
rect 43638 17250 43644 17284
rect 43678 17250 43684 17284
rect 43638 17212 43684 17250
rect 43638 17178 43644 17212
rect 43678 17178 43684 17212
rect 43638 17140 43684 17178
rect 43638 17120 43644 17140
rect 43380 17068 43426 17106
rect 43380 17034 43386 17068
rect 43420 17034 43426 17068
rect 43380 16996 43426 17034
rect 43380 16962 43386 16996
rect 43420 16962 43426 16996
rect 43380 16924 43426 16962
rect 43380 16890 43386 16924
rect 43420 16890 43426 16924
rect 43122 16843 43168 16873
rect 43380 16843 43426 16890
rect 43635 17106 43644 17120
rect 43678 17120 43684 17140
rect 43896 18821 44027 18843
rect 43896 18796 43934 18821
rect 43896 18762 43902 18796
rect 43986 18769 44027 18821
rect 43936 18762 44027 18769
rect 43896 18757 44027 18762
rect 43896 18724 43934 18757
rect 43896 18690 43902 18724
rect 43986 18705 44027 18757
rect 43936 18693 44027 18705
rect 43896 18652 43934 18690
rect 43896 18618 43902 18652
rect 43986 18641 44027 18693
rect 43936 18618 44027 18641
rect 43896 18610 44027 18618
rect 44154 18796 44200 18843
rect 44154 18762 44160 18796
rect 44194 18762 44200 18796
rect 44154 18724 44200 18762
rect 44154 18690 44160 18724
rect 44194 18690 44200 18724
rect 44154 18652 44200 18690
rect 44154 18618 44160 18652
rect 44194 18618 44200 18652
rect 43896 18580 43942 18610
rect 43896 18546 43902 18580
rect 43936 18546 43942 18580
rect 43896 18508 43942 18546
rect 43896 18474 43902 18508
rect 43936 18474 43942 18508
rect 43896 18436 43942 18474
rect 43896 18402 43902 18436
rect 43936 18402 43942 18436
rect 43896 18364 43942 18402
rect 43896 18330 43902 18364
rect 43936 18330 43942 18364
rect 43896 18292 43942 18330
rect 43896 18258 43902 18292
rect 43936 18258 43942 18292
rect 43896 18220 43942 18258
rect 43896 18186 43902 18220
rect 43936 18186 43942 18220
rect 43896 18148 43942 18186
rect 43896 18114 43902 18148
rect 43936 18114 43942 18148
rect 43896 18076 43942 18114
rect 43896 18042 43902 18076
rect 43936 18042 43942 18076
rect 43896 18004 43942 18042
rect 43896 17970 43902 18004
rect 43936 17970 43942 18004
rect 43896 17932 43942 17970
rect 43896 17898 43902 17932
rect 43936 17898 43942 17932
rect 43896 17860 43942 17898
rect 43896 17826 43902 17860
rect 43936 17826 43942 17860
rect 43896 17788 43942 17826
rect 43896 17754 43902 17788
rect 43936 17754 43942 17788
rect 43896 17716 43942 17754
rect 43896 17682 43902 17716
rect 43936 17682 43942 17716
rect 43896 17644 43942 17682
rect 43896 17610 43902 17644
rect 43936 17610 43942 17644
rect 43896 17572 43942 17610
rect 43896 17538 43902 17572
rect 43936 17538 43942 17572
rect 43896 17500 43942 17538
rect 43896 17466 43902 17500
rect 43936 17466 43942 17500
rect 43896 17428 43942 17466
rect 43896 17394 43902 17428
rect 43936 17394 43942 17428
rect 43896 17356 43942 17394
rect 43896 17322 43902 17356
rect 43936 17322 43942 17356
rect 43896 17284 43942 17322
rect 43896 17250 43902 17284
rect 43936 17250 43942 17284
rect 43896 17212 43942 17250
rect 43896 17178 43902 17212
rect 43936 17178 43942 17212
rect 43896 17140 43942 17178
rect 43678 17106 43765 17120
rect 43635 17090 43765 17106
rect 43635 17068 43672 17090
rect 43635 17034 43644 17068
rect 43724 17038 43765 17090
rect 43678 17034 43765 17038
rect 43635 17026 43765 17034
rect 43635 16996 43672 17026
rect 43635 16962 43644 16996
rect 43724 16974 43765 17026
rect 43678 16962 43765 16974
rect 43635 16924 43672 16962
rect 43635 16890 43644 16924
rect 43724 16910 43765 16962
rect 43678 16890 43765 16910
rect 43635 16879 43765 16890
rect 43896 17106 43902 17140
rect 43936 17106 43942 17140
rect 44154 18580 44200 18618
rect 44154 18546 44160 18580
rect 44194 18546 44200 18580
rect 44154 18508 44200 18546
rect 44154 18474 44160 18508
rect 44194 18474 44200 18508
rect 44154 18436 44200 18474
rect 44154 18402 44160 18436
rect 44194 18402 44200 18436
rect 44154 18364 44200 18402
rect 44154 18330 44160 18364
rect 44194 18330 44200 18364
rect 44154 18292 44200 18330
rect 44154 18258 44160 18292
rect 44194 18258 44200 18292
rect 44154 18220 44200 18258
rect 44154 18186 44160 18220
rect 44194 18186 44200 18220
rect 44154 18148 44200 18186
rect 44154 18114 44160 18148
rect 44194 18114 44200 18148
rect 44154 18076 44200 18114
rect 44154 18042 44160 18076
rect 44194 18042 44200 18076
rect 44154 18004 44200 18042
rect 44154 17970 44160 18004
rect 44194 17970 44200 18004
rect 44154 17932 44200 17970
rect 44154 17898 44160 17932
rect 44194 17898 44200 17932
rect 44154 17860 44200 17898
rect 44154 17826 44160 17860
rect 44194 17826 44200 17860
rect 44154 17788 44200 17826
rect 44154 17754 44160 17788
rect 44194 17754 44200 17788
rect 44154 17716 44200 17754
rect 44154 17682 44160 17716
rect 44194 17682 44200 17716
rect 44154 17644 44200 17682
rect 44154 17610 44160 17644
rect 44194 17610 44200 17644
rect 44154 17572 44200 17610
rect 44154 17538 44160 17572
rect 44194 17538 44200 17572
rect 44154 17500 44200 17538
rect 44154 17466 44160 17500
rect 44194 17466 44200 17500
rect 44154 17428 44200 17466
rect 44154 17394 44160 17428
rect 44194 17394 44200 17428
rect 44154 17356 44200 17394
rect 44154 17322 44160 17356
rect 44194 17322 44200 17356
rect 44154 17284 44200 17322
rect 44154 17250 44160 17284
rect 44194 17250 44200 17284
rect 44154 17212 44200 17250
rect 44154 17178 44160 17212
rect 44194 17178 44200 17212
rect 44154 17140 44200 17178
rect 44154 17121 44160 17140
rect 43896 17068 43942 17106
rect 43896 17034 43902 17068
rect 43936 17034 43942 17068
rect 43896 16996 43942 17034
rect 43896 16962 43902 16996
rect 43936 16962 43942 16996
rect 43896 16924 43942 16962
rect 43896 16890 43902 16924
rect 43936 16890 43942 16924
rect 43638 16843 43684 16879
rect 43896 16843 43942 16890
rect 44151 17106 44160 17121
rect 44194 17121 44200 17140
rect 44412 18813 44546 18843
rect 44412 18796 44453 18813
rect 44412 18762 44418 18796
rect 44452 18762 44453 18796
rect 44412 18761 44453 18762
rect 44505 18761 44546 18813
rect 44412 18749 44546 18761
rect 44412 18724 44453 18749
rect 44412 18690 44418 18724
rect 44452 18697 44453 18724
rect 44505 18697 44546 18749
rect 44452 18690 44546 18697
rect 44412 18685 44546 18690
rect 44412 18652 44453 18685
rect 44412 18618 44418 18652
rect 44452 18633 44453 18652
rect 44505 18633 44546 18685
rect 44452 18618 44546 18633
rect 44412 18602 44546 18618
rect 44670 18796 44716 18843
rect 44670 18762 44676 18796
rect 44710 18762 44716 18796
rect 44670 18724 44716 18762
rect 44670 18690 44676 18724
rect 44710 18690 44716 18724
rect 44670 18652 44716 18690
rect 44670 18618 44676 18652
rect 44710 18618 44716 18652
rect 44412 18580 44458 18602
rect 44412 18546 44418 18580
rect 44452 18546 44458 18580
rect 44412 18508 44458 18546
rect 44412 18474 44418 18508
rect 44452 18474 44458 18508
rect 44412 18436 44458 18474
rect 44412 18402 44418 18436
rect 44452 18402 44458 18436
rect 44412 18364 44458 18402
rect 44412 18330 44418 18364
rect 44452 18330 44458 18364
rect 44412 18292 44458 18330
rect 44412 18258 44418 18292
rect 44452 18258 44458 18292
rect 44412 18220 44458 18258
rect 44412 18186 44418 18220
rect 44452 18186 44458 18220
rect 44412 18148 44458 18186
rect 44412 18114 44418 18148
rect 44452 18114 44458 18148
rect 44412 18076 44458 18114
rect 44412 18042 44418 18076
rect 44452 18042 44458 18076
rect 44412 18004 44458 18042
rect 44412 17970 44418 18004
rect 44452 17970 44458 18004
rect 44412 17932 44458 17970
rect 44412 17898 44418 17932
rect 44452 17898 44458 17932
rect 44412 17860 44458 17898
rect 44412 17826 44418 17860
rect 44452 17826 44458 17860
rect 44412 17788 44458 17826
rect 44412 17754 44418 17788
rect 44452 17754 44458 17788
rect 44412 17716 44458 17754
rect 44412 17682 44418 17716
rect 44452 17682 44458 17716
rect 44412 17644 44458 17682
rect 44412 17610 44418 17644
rect 44452 17610 44458 17644
rect 44412 17572 44458 17610
rect 44412 17538 44418 17572
rect 44452 17538 44458 17572
rect 44412 17500 44458 17538
rect 44412 17466 44418 17500
rect 44452 17466 44458 17500
rect 44412 17428 44458 17466
rect 44412 17394 44418 17428
rect 44452 17394 44458 17428
rect 44412 17356 44458 17394
rect 44412 17322 44418 17356
rect 44452 17322 44458 17356
rect 44412 17284 44458 17322
rect 44412 17250 44418 17284
rect 44452 17250 44458 17284
rect 44412 17212 44458 17250
rect 44412 17178 44418 17212
rect 44452 17178 44458 17212
rect 44412 17140 44458 17178
rect 44194 17106 44281 17121
rect 44151 17091 44281 17106
rect 44151 17068 44188 17091
rect 44151 17034 44160 17068
rect 44240 17039 44281 17091
rect 44194 17034 44281 17039
rect 44151 17027 44281 17034
rect 44151 16996 44188 17027
rect 44151 16962 44160 16996
rect 44240 16975 44281 17027
rect 44194 16963 44281 16975
rect 44151 16924 44188 16962
rect 44151 16890 44160 16924
rect 44240 16911 44281 16963
rect 44194 16890 44281 16911
rect 44151 16880 44281 16890
rect 44412 17106 44418 17140
rect 44452 17106 44458 17140
rect 44412 17068 44458 17106
rect 44412 17034 44418 17068
rect 44452 17034 44458 17068
rect 44412 16996 44458 17034
rect 44412 16962 44418 16996
rect 44452 16962 44458 16996
rect 44412 16924 44458 16962
rect 44412 16890 44418 16924
rect 44452 16890 44458 16924
rect 44154 16843 44200 16880
rect 44412 16843 44458 16890
rect 44670 18580 44716 18618
rect 44927 18817 45057 18847
rect 44927 18796 44964 18817
rect 44927 18762 44934 18796
rect 45016 18765 45057 18817
rect 44968 18762 45057 18765
rect 44927 18753 45057 18762
rect 44927 18724 44964 18753
rect 44927 18690 44934 18724
rect 45016 18701 45057 18753
rect 44968 18690 45057 18701
rect 44927 18689 45057 18690
rect 44927 18652 44964 18689
rect 44927 18618 44934 18652
rect 45016 18637 45057 18689
rect 44968 18618 45057 18637
rect 44927 18606 45057 18618
rect 45186 18796 45232 18843
rect 45186 18762 45192 18796
rect 45226 18762 45232 18796
rect 45186 18724 45232 18762
rect 45186 18690 45192 18724
rect 45226 18690 45232 18724
rect 45186 18652 45232 18690
rect 45186 18618 45192 18652
rect 45226 18618 45232 18652
rect 44670 18546 44676 18580
rect 44710 18546 44716 18580
rect 44670 18508 44716 18546
rect 44670 18474 44676 18508
rect 44710 18474 44716 18508
rect 44670 18436 44716 18474
rect 44670 18402 44676 18436
rect 44710 18402 44716 18436
rect 44670 18364 44716 18402
rect 44670 18330 44676 18364
rect 44710 18330 44716 18364
rect 44670 18292 44716 18330
rect 44670 18258 44676 18292
rect 44710 18258 44716 18292
rect 44670 18220 44716 18258
rect 44670 18186 44676 18220
rect 44710 18186 44716 18220
rect 44670 18148 44716 18186
rect 44670 18114 44676 18148
rect 44710 18114 44716 18148
rect 44670 18076 44716 18114
rect 44670 18042 44676 18076
rect 44710 18042 44716 18076
rect 44670 18004 44716 18042
rect 44670 17970 44676 18004
rect 44710 17970 44716 18004
rect 44670 17932 44716 17970
rect 44670 17898 44676 17932
rect 44710 17898 44716 17932
rect 44670 17860 44716 17898
rect 44670 17826 44676 17860
rect 44710 17826 44716 17860
rect 44670 17788 44716 17826
rect 44670 17754 44676 17788
rect 44710 17754 44716 17788
rect 44670 17716 44716 17754
rect 44670 17682 44676 17716
rect 44710 17682 44716 17716
rect 44670 17644 44716 17682
rect 44670 17610 44676 17644
rect 44710 17610 44716 17644
rect 44670 17572 44716 17610
rect 44670 17538 44676 17572
rect 44710 17538 44716 17572
rect 44670 17500 44716 17538
rect 44670 17466 44676 17500
rect 44710 17466 44716 17500
rect 44670 17428 44716 17466
rect 44670 17394 44676 17428
rect 44710 17394 44716 17428
rect 44670 17356 44716 17394
rect 44670 17322 44676 17356
rect 44710 17322 44716 17356
rect 44670 17284 44716 17322
rect 44670 17250 44676 17284
rect 44710 17250 44716 17284
rect 44670 17212 44716 17250
rect 44670 17178 44676 17212
rect 44710 17178 44716 17212
rect 44670 17140 44716 17178
rect 44670 17106 44676 17140
rect 44710 17124 44716 17140
rect 44928 18580 44974 18606
rect 44928 18546 44934 18580
rect 44968 18546 44974 18580
rect 44928 18508 44974 18546
rect 44928 18474 44934 18508
rect 44968 18474 44974 18508
rect 44928 18436 44974 18474
rect 44928 18402 44934 18436
rect 44968 18402 44974 18436
rect 44928 18364 44974 18402
rect 44928 18330 44934 18364
rect 44968 18330 44974 18364
rect 44928 18292 44974 18330
rect 44928 18258 44934 18292
rect 44968 18258 44974 18292
rect 44928 18220 44974 18258
rect 44928 18186 44934 18220
rect 44968 18186 44974 18220
rect 44928 18148 44974 18186
rect 44928 18114 44934 18148
rect 44968 18114 44974 18148
rect 44928 18076 44974 18114
rect 44928 18042 44934 18076
rect 44968 18042 44974 18076
rect 44928 18004 44974 18042
rect 44928 17970 44934 18004
rect 44968 17970 44974 18004
rect 44928 17932 44974 17970
rect 44928 17898 44934 17932
rect 44968 17898 44974 17932
rect 44928 17860 44974 17898
rect 44928 17826 44934 17860
rect 44968 17826 44974 17860
rect 44928 17788 44974 17826
rect 44928 17754 44934 17788
rect 44968 17754 44974 17788
rect 44928 17716 44974 17754
rect 44928 17682 44934 17716
rect 44968 17682 44974 17716
rect 44928 17644 44974 17682
rect 44928 17610 44934 17644
rect 44968 17610 44974 17644
rect 44928 17572 44974 17610
rect 44928 17538 44934 17572
rect 44968 17538 44974 17572
rect 44928 17500 44974 17538
rect 44928 17466 44934 17500
rect 44968 17466 44974 17500
rect 44928 17428 44974 17466
rect 44928 17394 44934 17428
rect 44968 17394 44974 17428
rect 44928 17356 44974 17394
rect 44928 17322 44934 17356
rect 44968 17322 44974 17356
rect 44928 17284 44974 17322
rect 44928 17250 44934 17284
rect 44968 17250 44974 17284
rect 44928 17212 44974 17250
rect 44928 17178 44934 17212
rect 44968 17178 44974 17212
rect 44928 17140 44974 17178
rect 44710 17106 44803 17124
rect 44670 17094 44803 17106
rect 44670 17068 44710 17094
rect 44670 17034 44676 17068
rect 44762 17042 44803 17094
rect 44710 17034 44803 17042
rect 44670 17030 44803 17034
rect 44670 16996 44710 17030
rect 44670 16962 44676 16996
rect 44762 16978 44803 17030
rect 44710 16966 44803 16978
rect 44670 16924 44710 16962
rect 44670 16890 44676 16924
rect 44762 16914 44803 16966
rect 44710 16890 44803 16914
rect 44670 16883 44803 16890
rect 44928 17106 44934 17140
rect 44968 17106 44974 17140
rect 45186 18580 45232 18618
rect 45186 18546 45192 18580
rect 45226 18546 45232 18580
rect 45186 18508 45232 18546
rect 45186 18474 45192 18508
rect 45226 18474 45232 18508
rect 45186 18436 45232 18474
rect 45186 18402 45192 18436
rect 45226 18402 45232 18436
rect 45186 18364 45232 18402
rect 45186 18330 45192 18364
rect 45226 18330 45232 18364
rect 45186 18292 45232 18330
rect 45186 18258 45192 18292
rect 45226 18258 45232 18292
rect 45186 18220 45232 18258
rect 45186 18186 45192 18220
rect 45226 18186 45232 18220
rect 45186 18148 45232 18186
rect 45186 18114 45192 18148
rect 45226 18114 45232 18148
rect 45186 18076 45232 18114
rect 45186 18042 45192 18076
rect 45226 18042 45232 18076
rect 45186 18004 45232 18042
rect 45186 17970 45192 18004
rect 45226 17970 45232 18004
rect 45186 17932 45232 17970
rect 45186 17898 45192 17932
rect 45226 17898 45232 17932
rect 45186 17860 45232 17898
rect 45186 17826 45192 17860
rect 45226 17826 45232 17860
rect 45186 17788 45232 17826
rect 45186 17754 45192 17788
rect 45226 17754 45232 17788
rect 45186 17716 45232 17754
rect 45186 17682 45192 17716
rect 45226 17682 45232 17716
rect 45186 17644 45232 17682
rect 45186 17610 45192 17644
rect 45226 17610 45232 17644
rect 45186 17572 45232 17610
rect 45186 17538 45192 17572
rect 45226 17538 45232 17572
rect 45186 17500 45232 17538
rect 45186 17466 45192 17500
rect 45226 17466 45232 17500
rect 45186 17428 45232 17466
rect 45186 17394 45192 17428
rect 45226 17394 45232 17428
rect 45186 17356 45232 17394
rect 45186 17322 45192 17356
rect 45226 17322 45232 17356
rect 45186 17284 45232 17322
rect 45186 17250 45192 17284
rect 45226 17250 45232 17284
rect 45186 17212 45232 17250
rect 45186 17178 45192 17212
rect 45226 17178 45232 17212
rect 45186 17140 45232 17178
rect 45186 17118 45192 17140
rect 44928 17068 44974 17106
rect 44928 17034 44934 17068
rect 44968 17034 44974 17068
rect 44928 16996 44974 17034
rect 44928 16962 44934 16996
rect 44968 16962 44974 16996
rect 44928 16924 44974 16962
rect 44928 16890 44934 16924
rect 44968 16890 44974 16924
rect 44670 16843 44716 16883
rect 44928 16843 44974 16890
rect 45179 17106 45192 17118
rect 45226 17118 45232 17140
rect 45530 18213 46586 18320
rect 45226 17106 45309 17118
rect 45179 17088 45309 17106
rect 45179 17068 45216 17088
rect 45179 17034 45192 17068
rect 45268 17036 45309 17088
rect 45226 17034 45309 17036
rect 45179 17024 45309 17034
rect 45179 16996 45216 17024
rect 45179 16962 45192 16996
rect 45268 16972 45309 17024
rect 45226 16962 45309 16972
rect 45179 16960 45309 16962
rect 45179 16924 45216 16960
rect 45179 16890 45192 16924
rect 45268 16908 45309 16960
rect 45226 16890 45309 16908
rect 45179 16877 45309 16890
rect 45530 16881 45602 18213
rect 46486 16881 46586 18213
rect 45186 16843 45232 16877
rect 45530 16814 46586 16881
rect 42662 16796 42854 16802
rect 42662 16766 42705 16796
rect 41638 16762 42705 16766
rect 42739 16762 42777 16796
rect 42811 16766 42854 16796
rect 42920 16796 43112 16802
rect 42920 16766 42963 16796
rect 42811 16762 42963 16766
rect 42997 16762 43035 16796
rect 43069 16766 43112 16796
rect 43178 16796 43370 16802
rect 43178 16766 43221 16796
rect 43069 16762 43221 16766
rect 43255 16762 43293 16796
rect 43327 16766 43370 16796
rect 43436 16796 43628 16802
rect 43436 16766 43479 16796
rect 43327 16762 43479 16766
rect 43513 16762 43551 16796
rect 43585 16766 43628 16796
rect 43694 16796 43886 16802
rect 43694 16766 43737 16796
rect 43585 16762 43737 16766
rect 43771 16762 43809 16796
rect 43843 16766 43886 16796
rect 43952 16796 44144 16802
rect 43952 16766 43995 16796
rect 43843 16762 43995 16766
rect 44029 16762 44067 16796
rect 44101 16766 44144 16796
rect 44210 16796 44402 16802
rect 44210 16766 44253 16796
rect 44101 16762 44253 16766
rect 44287 16762 44325 16796
rect 44359 16766 44402 16796
rect 44468 16796 44660 16802
rect 44468 16766 44511 16796
rect 44359 16762 44511 16766
rect 44545 16762 44583 16796
rect 44617 16766 44660 16796
rect 44726 16796 44918 16802
rect 44726 16766 44769 16796
rect 44617 16762 44769 16766
rect 44803 16762 44841 16796
rect 44875 16766 44918 16796
rect 44984 16796 45176 16802
rect 44984 16766 45027 16796
rect 44875 16762 45027 16766
rect 45061 16762 45099 16796
rect 45133 16766 45176 16796
rect 45133 16762 45188 16766
rect 41638 16686 45188 16762
rect 27122 16222 28082 16248
rect 24590 15932 24609 15966
rect 24643 15932 24681 15966
rect 24715 15932 24753 15966
rect 24787 15932 24825 15966
rect 24859 15932 24897 15966
rect 24931 15932 24969 15966
rect 25003 15932 25023 15966
rect 24590 15912 25023 15932
rect 27121 15966 27554 15985
rect 27121 15932 27140 15966
rect 27174 15932 27212 15966
rect 27246 15932 27284 15966
rect 27318 15932 27356 15966
rect 27390 15932 27428 15966
rect 27462 15932 27500 15966
rect 27534 15932 27554 15966
rect 39497 15962 39895 15963
rect 37999 15961 40679 15962
rect 22522 15712 22962 15745
rect 23819 15648 25022 15672
rect 23819 15614 24609 15648
rect 24643 15614 24681 15648
rect 24715 15614 24753 15648
rect 24787 15614 24825 15648
rect 24859 15614 24897 15648
rect 24931 15614 24969 15648
rect 25003 15614 25022 15648
rect 23819 15584 25022 15614
rect 27121 15648 27554 15932
rect 27121 15614 27140 15648
rect 27174 15614 27212 15648
rect 27246 15614 27284 15648
rect 27318 15614 27356 15648
rect 27390 15614 27428 15648
rect 27462 15614 27500 15648
rect 27534 15614 27554 15648
rect 27121 15594 27554 15614
rect 36395 15921 40679 15961
rect 36395 15913 40586 15921
rect 36395 15807 38517 15913
rect 38767 15912 40586 15913
rect 38767 15807 39533 15912
rect 36395 15806 39533 15807
rect 39855 15887 40586 15912
rect 40620 15887 40679 15921
rect 39855 15849 40679 15887
rect 39855 15815 40586 15849
rect 40620 15815 40679 15849
rect 39855 15806 40679 15815
rect 36395 15747 40679 15806
rect 36395 15695 38413 15747
rect 10297 15011 10358 15018
rect 11256 15011 11322 15018
rect 10297 14952 11322 15011
rect -3949 14851 -3862 14885
rect -3828 14851 -3776 14885
rect 16552 14864 17162 14890
rect 16552 14858 18116 14864
rect 16552 14854 17171 14858
rect -7465 14788 -7419 14835
rect -7465 14754 -7459 14788
rect -7425 14754 -7419 14788
rect -7465 14716 -7419 14754
rect -7465 14682 -7459 14716
rect -7425 14682 -7419 14716
rect -7465 14644 -7419 14682
rect -7465 14610 -7459 14644
rect -7425 14610 -7419 14644
rect -7465 14572 -7419 14610
rect -7465 14538 -7459 14572
rect -7425 14538 -7419 14572
rect -7465 14500 -7419 14538
rect -7465 14466 -7459 14500
rect -7425 14466 -7419 14500
rect -7465 14428 -7419 14466
rect -7465 14394 -7459 14428
rect -7425 14394 -7419 14428
rect -7465 14356 -7419 14394
rect -7465 14322 -7459 14356
rect -7425 14322 -7419 14356
rect -7465 14284 -7419 14322
rect -7465 14250 -7459 14284
rect -7425 14250 -7419 14284
rect -7465 14212 -7419 14250
rect -7465 14178 -7459 14212
rect -7425 14178 -7419 14212
rect -7465 14140 -7419 14178
rect -7465 14106 -7459 14140
rect -7425 14106 -7419 14140
rect -7465 14068 -7419 14106
rect -7465 14034 -7459 14068
rect -7425 14034 -7419 14068
rect -7465 13996 -7419 14034
rect -7465 13962 -7459 13996
rect -7425 13962 -7419 13996
rect -7465 13924 -7419 13962
rect -7465 13890 -7459 13924
rect -7425 13890 -7419 13924
rect -7465 13852 -7419 13890
rect -7465 13818 -7459 13852
rect -7425 13818 -7419 13852
rect -7465 13780 -7419 13818
rect -7465 13746 -7459 13780
rect -7425 13746 -7419 13780
rect -7465 13708 -7419 13746
rect -7465 13674 -7459 13708
rect -7425 13674 -7419 13708
rect -7465 13636 -7419 13674
rect -7465 13602 -7459 13636
rect -7425 13602 -7419 13636
rect -7465 13564 -7419 13602
rect -7465 13530 -7459 13564
rect -7425 13530 -7419 13564
rect -7465 13492 -7419 13530
rect -7465 13458 -7459 13492
rect -7425 13458 -7419 13492
rect -7465 13420 -7419 13458
rect -7465 13386 -7459 13420
rect -7425 13386 -7419 13420
rect -7465 13348 -7419 13386
rect -7465 13314 -7459 13348
rect -7425 13314 -7419 13348
rect -7465 13276 -7419 13314
rect -7465 13242 -7459 13276
rect -7425 13242 -7419 13276
rect -7465 13204 -7419 13242
rect -7465 13170 -7459 13204
rect -7425 13170 -7419 13204
rect -7465 13132 -7419 13170
rect -7465 13119 -7459 13132
rect -7500 13098 -7459 13119
rect -7425 13119 -7419 13132
rect -7207 14788 -7161 14835
rect -6949 14822 -6903 14835
rect -7207 14754 -7201 14788
rect -7167 14754 -7161 14788
rect -7207 14716 -7161 14754
rect -7207 14682 -7201 14716
rect -7167 14682 -7161 14716
rect -7207 14644 -7161 14682
rect -7207 14610 -7201 14644
rect -7167 14610 -7161 14644
rect -7207 14572 -7161 14610
rect -7207 14538 -7201 14572
rect -7167 14538 -7161 14572
rect -7207 14500 -7161 14538
rect -6994 14788 -6844 14822
rect -6994 14768 -6943 14788
rect -6909 14768 -6844 14788
rect -6994 14716 -6947 14768
rect -6895 14716 -6844 14768
rect -6994 14704 -6943 14716
rect -6909 14704 -6844 14716
rect -6994 14652 -6947 14704
rect -6895 14652 -6844 14704
rect -6994 14644 -6844 14652
rect -6994 14640 -6943 14644
rect -6909 14640 -6844 14644
rect -6994 14588 -6947 14640
rect -6895 14588 -6844 14640
rect -6994 14572 -6844 14588
rect -6994 14538 -6943 14572
rect -6909 14538 -6844 14572
rect -6994 14536 -6844 14538
rect -6691 14788 -6645 14835
rect -6691 14754 -6685 14788
rect -6651 14754 -6645 14788
rect -6691 14716 -6645 14754
rect -6691 14682 -6685 14716
rect -6651 14682 -6645 14716
rect -6691 14644 -6645 14682
rect -6691 14610 -6685 14644
rect -6651 14610 -6645 14644
rect -6691 14572 -6645 14610
rect -6691 14538 -6685 14572
rect -6651 14538 -6645 14572
rect -7207 14466 -7201 14500
rect -7167 14466 -7161 14500
rect -7207 14428 -7161 14466
rect -7207 14394 -7201 14428
rect -7167 14394 -7161 14428
rect -7207 14356 -7161 14394
rect -7207 14322 -7201 14356
rect -7167 14322 -7161 14356
rect -7207 14284 -7161 14322
rect -7207 14250 -7201 14284
rect -7167 14250 -7161 14284
rect -7207 14212 -7161 14250
rect -7207 14178 -7201 14212
rect -7167 14178 -7161 14212
rect -7207 14140 -7161 14178
rect -7207 14106 -7201 14140
rect -7167 14106 -7161 14140
rect -7207 14068 -7161 14106
rect -7207 14034 -7201 14068
rect -7167 14034 -7161 14068
rect -7207 13996 -7161 14034
rect -7207 13962 -7201 13996
rect -7167 13962 -7161 13996
rect -7207 13924 -7161 13962
rect -7207 13890 -7201 13924
rect -7167 13890 -7161 13924
rect -7207 13852 -7161 13890
rect -7207 13818 -7201 13852
rect -7167 13818 -7161 13852
rect -7207 13780 -7161 13818
rect -7207 13746 -7201 13780
rect -7167 13746 -7161 13780
rect -7207 13708 -7161 13746
rect -7207 13674 -7201 13708
rect -7167 13674 -7161 13708
rect -7207 13636 -7161 13674
rect -7207 13602 -7201 13636
rect -7167 13602 -7161 13636
rect -7207 13564 -7161 13602
rect -7207 13530 -7201 13564
rect -7167 13530 -7161 13564
rect -7207 13492 -7161 13530
rect -7207 13458 -7201 13492
rect -7167 13458 -7161 13492
rect -7207 13420 -7161 13458
rect -7207 13386 -7201 13420
rect -7167 13386 -7161 13420
rect -7207 13348 -7161 13386
rect -7207 13314 -7201 13348
rect -7167 13314 -7161 13348
rect -7207 13276 -7161 13314
rect -7207 13242 -7201 13276
rect -7167 13242 -7161 13276
rect -7207 13204 -7161 13242
rect -7207 13170 -7201 13204
rect -7167 13170 -7161 13204
rect -7207 13132 -7161 13170
rect -7425 13098 -7350 13119
rect -7500 13065 -7350 13098
rect -7500 13060 -7453 13065
rect -7500 13026 -7459 13060
rect -7500 13013 -7453 13026
rect -7401 13013 -7350 13065
rect -7500 13001 -7350 13013
rect -7500 12988 -7453 13001
rect -7500 12954 -7459 12988
rect -7500 12949 -7453 12954
rect -7401 12949 -7350 13001
rect -7500 12937 -7350 12949
rect -7500 12916 -7453 12937
rect -7500 12882 -7459 12916
rect -7401 12885 -7350 12937
rect -7425 12882 -7350 12885
rect -7500 12833 -7350 12882
rect -7207 13098 -7201 13132
rect -7167 13098 -7161 13132
rect -7207 13060 -7161 13098
rect -7207 13026 -7201 13060
rect -7167 13026 -7161 13060
rect -7207 12988 -7161 13026
rect -7207 12954 -7201 12988
rect -7167 12954 -7161 12988
rect -7207 12916 -7161 12954
rect -7207 12882 -7201 12916
rect -7167 12882 -7161 12916
rect -7207 12835 -7161 12882
rect -6949 14500 -6903 14536
rect -6949 14466 -6943 14500
rect -6909 14466 -6903 14500
rect -6949 14428 -6903 14466
rect -6949 14394 -6943 14428
rect -6909 14394 -6903 14428
rect -6949 14356 -6903 14394
rect -6949 14322 -6943 14356
rect -6909 14322 -6903 14356
rect -6949 14284 -6903 14322
rect -6949 14250 -6943 14284
rect -6909 14250 -6903 14284
rect -6949 14212 -6903 14250
rect -6949 14178 -6943 14212
rect -6909 14178 -6903 14212
rect -6949 14140 -6903 14178
rect -6949 14106 -6943 14140
rect -6909 14106 -6903 14140
rect -6949 14068 -6903 14106
rect -6949 14034 -6943 14068
rect -6909 14034 -6903 14068
rect -6949 13996 -6903 14034
rect -6949 13962 -6943 13996
rect -6909 13962 -6903 13996
rect -6949 13924 -6903 13962
rect -6949 13890 -6943 13924
rect -6909 13890 -6903 13924
rect -6949 13852 -6903 13890
rect -6949 13818 -6943 13852
rect -6909 13818 -6903 13852
rect -6949 13780 -6903 13818
rect -6949 13746 -6943 13780
rect -6909 13746 -6903 13780
rect -6949 13708 -6903 13746
rect -6949 13674 -6943 13708
rect -6909 13674 -6903 13708
rect -6949 13636 -6903 13674
rect -6949 13602 -6943 13636
rect -6909 13602 -6903 13636
rect -6949 13564 -6903 13602
rect -6949 13530 -6943 13564
rect -6909 13530 -6903 13564
rect -6949 13492 -6903 13530
rect -6949 13458 -6943 13492
rect -6909 13458 -6903 13492
rect -6949 13420 -6903 13458
rect -6949 13386 -6943 13420
rect -6909 13386 -6903 13420
rect -6949 13348 -6903 13386
rect -6949 13314 -6943 13348
rect -6909 13314 -6903 13348
rect -6949 13276 -6903 13314
rect -6949 13242 -6943 13276
rect -6909 13242 -6903 13276
rect -6949 13204 -6903 13242
rect -6949 13170 -6943 13204
rect -6909 13170 -6903 13204
rect -6949 13132 -6903 13170
rect -6949 13098 -6943 13132
rect -6909 13098 -6903 13132
rect -6949 13060 -6903 13098
rect -6949 13026 -6943 13060
rect -6909 13026 -6903 13060
rect -6949 12988 -6903 13026
rect -6949 12954 -6943 12988
rect -6909 12954 -6903 12988
rect -6949 12916 -6903 12954
rect -6949 12882 -6943 12916
rect -6909 12882 -6903 12916
rect -6949 12835 -6903 12882
rect -6691 14500 -6645 14538
rect -6691 14466 -6685 14500
rect -6651 14466 -6645 14500
rect -6691 14428 -6645 14466
rect -6691 14394 -6685 14428
rect -6651 14394 -6645 14428
rect -6691 14356 -6645 14394
rect -6691 14322 -6685 14356
rect -6651 14322 -6645 14356
rect -6691 14284 -6645 14322
rect -6691 14250 -6685 14284
rect -6651 14250 -6645 14284
rect -6691 14212 -6645 14250
rect -6691 14178 -6685 14212
rect -6651 14178 -6645 14212
rect -6691 14140 -6645 14178
rect -6691 14106 -6685 14140
rect -6651 14106 -6645 14140
rect -6691 14068 -6645 14106
rect -6691 14034 -6685 14068
rect -6651 14034 -6645 14068
rect -6691 13996 -6645 14034
rect -6691 13962 -6685 13996
rect -6651 13962 -6645 13996
rect -6691 13924 -6645 13962
rect -6691 13890 -6685 13924
rect -6651 13890 -6645 13924
rect -6691 13852 -6645 13890
rect -6691 13818 -6685 13852
rect -6651 13818 -6645 13852
rect -6691 13780 -6645 13818
rect -6691 13746 -6685 13780
rect -6651 13746 -6645 13780
rect -6691 13708 -6645 13746
rect -6691 13674 -6685 13708
rect -6651 13674 -6645 13708
rect -6691 13636 -6645 13674
rect -6691 13602 -6685 13636
rect -6651 13602 -6645 13636
rect -6691 13564 -6645 13602
rect -6691 13530 -6685 13564
rect -6651 13530 -6645 13564
rect -6691 13492 -6645 13530
rect -6691 13458 -6685 13492
rect -6651 13458 -6645 13492
rect -6691 13420 -6645 13458
rect -6691 13386 -6685 13420
rect -6651 13386 -6645 13420
rect -6691 13348 -6645 13386
rect -6691 13314 -6685 13348
rect -6651 13314 -6645 13348
rect -6691 13276 -6645 13314
rect -6691 13242 -6685 13276
rect -6651 13242 -6645 13276
rect -6691 13204 -6645 13242
rect -6691 13170 -6685 13204
rect -6651 13170 -6645 13204
rect -6691 13132 -6645 13170
rect -6691 13098 -6685 13132
rect -6651 13098 -6645 13132
rect -6433 14788 -6387 14835
rect -6433 14754 -6427 14788
rect -6393 14754 -6387 14788
rect -6433 14716 -6387 14754
rect -6433 14682 -6427 14716
rect -6393 14682 -6387 14716
rect -6433 14644 -6387 14682
rect -6433 14610 -6427 14644
rect -6393 14610 -6387 14644
rect -6433 14572 -6387 14610
rect -6433 14538 -6427 14572
rect -6393 14538 -6387 14572
rect -6433 14500 -6387 14538
rect -6433 14466 -6427 14500
rect -6393 14466 -6387 14500
rect -6433 14428 -6387 14466
rect -6433 14394 -6427 14428
rect -6393 14394 -6387 14428
rect -6433 14356 -6387 14394
rect -6433 14322 -6427 14356
rect -6393 14322 -6387 14356
rect -6433 14284 -6387 14322
rect -6433 14250 -6427 14284
rect -6393 14250 -6387 14284
rect -6433 14212 -6387 14250
rect -6433 14178 -6427 14212
rect -6393 14178 -6387 14212
rect -6433 14140 -6387 14178
rect -6433 14106 -6427 14140
rect -6393 14106 -6387 14140
rect -6433 14068 -6387 14106
rect -6433 14034 -6427 14068
rect -6393 14034 -6387 14068
rect -6433 13996 -6387 14034
rect -6433 13962 -6427 13996
rect -6393 13962 -6387 13996
rect -6433 13924 -6387 13962
rect -6433 13890 -6427 13924
rect -6393 13890 -6387 13924
rect -6433 13852 -6387 13890
rect -6433 13818 -6427 13852
rect -6393 13818 -6387 13852
rect -6433 13780 -6387 13818
rect -6433 13746 -6427 13780
rect -6393 13746 -6387 13780
rect -6433 13708 -6387 13746
rect -6433 13674 -6427 13708
rect -6393 13674 -6387 13708
rect -6433 13636 -6387 13674
rect -6433 13602 -6427 13636
rect -6393 13602 -6387 13636
rect -6433 13564 -6387 13602
rect -6433 13530 -6427 13564
rect -6393 13530 -6387 13564
rect -6433 13492 -6387 13530
rect -6433 13458 -6427 13492
rect -6393 13458 -6387 13492
rect -6433 13420 -6387 13458
rect -6433 13386 -6427 13420
rect -6393 13386 -6387 13420
rect -6433 13348 -6387 13386
rect -6433 13314 -6427 13348
rect -6393 13314 -6387 13348
rect -6433 13276 -6387 13314
rect -6433 13242 -6427 13276
rect -6393 13242 -6387 13276
rect -6433 13204 -6387 13242
rect -6433 13170 -6427 13204
rect -6393 13170 -6387 13204
rect -6433 13132 -6387 13170
rect -6433 13130 -6427 13132
rect -6691 13060 -6645 13098
rect -6691 13026 -6685 13060
rect -6651 13026 -6645 13060
rect -6691 12988 -6645 13026
rect -6691 12954 -6685 12988
rect -6651 12954 -6645 12988
rect -6691 12916 -6645 12954
rect -6691 12882 -6685 12916
rect -6651 12882 -6645 12916
rect -6691 12835 -6645 12882
rect -6481 13098 -6427 13130
rect -6393 13130 -6387 13132
rect -6175 14788 -6129 14835
rect -5917 14809 -5871 14835
rect -6175 14754 -6169 14788
rect -6135 14754 -6129 14788
rect -6175 14716 -6129 14754
rect -6175 14682 -6169 14716
rect -6135 14682 -6129 14716
rect -6175 14644 -6129 14682
rect -6175 14610 -6169 14644
rect -6135 14610 -6129 14644
rect -6175 14572 -6129 14610
rect -6175 14538 -6169 14572
rect -6135 14538 -6129 14572
rect -6175 14500 -6129 14538
rect -5983 14788 -5833 14809
rect -5983 14755 -5911 14788
rect -5983 14703 -5936 14755
rect -5877 14754 -5833 14788
rect -5884 14716 -5833 14754
rect -5983 14691 -5911 14703
rect -5983 14639 -5936 14691
rect -5877 14682 -5833 14716
rect -5884 14644 -5833 14682
rect -5983 14627 -5911 14639
rect -5983 14575 -5936 14627
rect -5877 14610 -5833 14644
rect -5884 14575 -5833 14610
rect -5983 14572 -5833 14575
rect -5983 14538 -5911 14572
rect -5877 14538 -5833 14572
rect -5983 14523 -5833 14538
rect -5659 14788 -5613 14835
rect -5659 14754 -5653 14788
rect -5619 14754 -5613 14788
rect -5659 14716 -5613 14754
rect -5659 14682 -5653 14716
rect -5619 14682 -5613 14716
rect -5659 14644 -5613 14682
rect -5659 14610 -5653 14644
rect -5619 14610 -5613 14644
rect -5659 14572 -5613 14610
rect -5659 14538 -5653 14572
rect -5619 14538 -5613 14572
rect -6175 14466 -6169 14500
rect -6135 14466 -6129 14500
rect -6175 14428 -6129 14466
rect -6175 14394 -6169 14428
rect -6135 14394 -6129 14428
rect -6175 14356 -6129 14394
rect -6175 14322 -6169 14356
rect -6135 14322 -6129 14356
rect -6175 14284 -6129 14322
rect -6175 14250 -6169 14284
rect -6135 14250 -6129 14284
rect -6175 14212 -6129 14250
rect -6175 14178 -6169 14212
rect -6135 14178 -6129 14212
rect -6175 14140 -6129 14178
rect -6175 14106 -6169 14140
rect -6135 14106 -6129 14140
rect -6175 14068 -6129 14106
rect -6175 14034 -6169 14068
rect -6135 14034 -6129 14068
rect -6175 13996 -6129 14034
rect -6175 13962 -6169 13996
rect -6135 13962 -6129 13996
rect -6175 13924 -6129 13962
rect -6175 13890 -6169 13924
rect -6135 13890 -6129 13924
rect -6175 13852 -6129 13890
rect -6175 13818 -6169 13852
rect -6135 13818 -6129 13852
rect -6175 13780 -6129 13818
rect -6175 13746 -6169 13780
rect -6135 13746 -6129 13780
rect -6175 13708 -6129 13746
rect -6175 13674 -6169 13708
rect -6135 13674 -6129 13708
rect -6175 13636 -6129 13674
rect -6175 13602 -6169 13636
rect -6135 13602 -6129 13636
rect -6175 13564 -6129 13602
rect -6175 13530 -6169 13564
rect -6135 13530 -6129 13564
rect -6175 13492 -6129 13530
rect -6175 13458 -6169 13492
rect -6135 13458 -6129 13492
rect -6175 13420 -6129 13458
rect -6175 13386 -6169 13420
rect -6135 13386 -6129 13420
rect -6175 13348 -6129 13386
rect -6175 13314 -6169 13348
rect -6135 13314 -6129 13348
rect -6175 13276 -6129 13314
rect -6175 13242 -6169 13276
rect -6135 13242 -6129 13276
rect -6175 13204 -6129 13242
rect -6175 13170 -6169 13204
rect -6135 13170 -6129 13204
rect -6175 13132 -6129 13170
rect -6393 13098 -6331 13130
rect -6481 13076 -6331 13098
rect -6481 13024 -6434 13076
rect -6382 13024 -6331 13076
rect -6481 13012 -6331 13024
rect -6481 12960 -6434 13012
rect -6382 12960 -6331 13012
rect -6481 12954 -6427 12960
rect -6393 12954 -6331 12960
rect -6481 12948 -6331 12954
rect -6481 12896 -6434 12948
rect -6382 12896 -6331 12948
rect -6481 12882 -6427 12896
rect -6393 12882 -6331 12896
rect -6481 12844 -6331 12882
rect -6175 13098 -6169 13132
rect -6135 13098 -6129 13132
rect -6175 13060 -6129 13098
rect -6175 13026 -6169 13060
rect -6135 13026 -6129 13060
rect -6175 12988 -6129 13026
rect -6175 12954 -6169 12988
rect -6135 12954 -6129 12988
rect -6175 12916 -6129 12954
rect -6175 12882 -6169 12916
rect -6135 12882 -6129 12916
rect -6433 12835 -6387 12844
rect -6175 12835 -6129 12882
rect -5917 14500 -5871 14523
rect -5917 14466 -5911 14500
rect -5877 14466 -5871 14500
rect -5917 14428 -5871 14466
rect -5917 14394 -5911 14428
rect -5877 14394 -5871 14428
rect -5917 14356 -5871 14394
rect -5917 14322 -5911 14356
rect -5877 14322 -5871 14356
rect -5917 14284 -5871 14322
rect -5917 14250 -5911 14284
rect -5877 14250 -5871 14284
rect -5917 14212 -5871 14250
rect -5917 14178 -5911 14212
rect -5877 14178 -5871 14212
rect -5917 14140 -5871 14178
rect -5917 14106 -5911 14140
rect -5877 14106 -5871 14140
rect -5917 14068 -5871 14106
rect -5917 14034 -5911 14068
rect -5877 14034 -5871 14068
rect -5917 13996 -5871 14034
rect -5917 13962 -5911 13996
rect -5877 13962 -5871 13996
rect -5917 13924 -5871 13962
rect -5917 13890 -5911 13924
rect -5877 13890 -5871 13924
rect -5917 13852 -5871 13890
rect -5917 13818 -5911 13852
rect -5877 13818 -5871 13852
rect -5917 13780 -5871 13818
rect -5917 13746 -5911 13780
rect -5877 13746 -5871 13780
rect -5917 13708 -5871 13746
rect -5917 13674 -5911 13708
rect -5877 13674 -5871 13708
rect -5917 13636 -5871 13674
rect -5917 13602 -5911 13636
rect -5877 13602 -5871 13636
rect -5917 13564 -5871 13602
rect -5917 13530 -5911 13564
rect -5877 13530 -5871 13564
rect -5917 13492 -5871 13530
rect -5917 13458 -5911 13492
rect -5877 13458 -5871 13492
rect -5917 13420 -5871 13458
rect -5917 13386 -5911 13420
rect -5877 13386 -5871 13420
rect -5917 13348 -5871 13386
rect -5917 13314 -5911 13348
rect -5877 13314 -5871 13348
rect -5917 13276 -5871 13314
rect -5917 13242 -5911 13276
rect -5877 13242 -5871 13276
rect -5917 13204 -5871 13242
rect -5917 13170 -5911 13204
rect -5877 13170 -5871 13204
rect -5917 13132 -5871 13170
rect -5917 13098 -5911 13132
rect -5877 13098 -5871 13132
rect -5917 13060 -5871 13098
rect -5917 13026 -5911 13060
rect -5877 13026 -5871 13060
rect -5917 12988 -5871 13026
rect -5917 12954 -5911 12988
rect -5877 12954 -5871 12988
rect -5917 12916 -5871 12954
rect -5917 12882 -5911 12916
rect -5877 12882 -5871 12916
rect -5917 12835 -5871 12882
rect -5659 14500 -5613 14538
rect -5659 14466 -5653 14500
rect -5619 14466 -5613 14500
rect -5659 14428 -5613 14466
rect -5659 14394 -5653 14428
rect -5619 14394 -5613 14428
rect -5659 14356 -5613 14394
rect -5659 14322 -5653 14356
rect -5619 14322 -5613 14356
rect -5659 14284 -5613 14322
rect -5659 14250 -5653 14284
rect -5619 14250 -5613 14284
rect -5659 14212 -5613 14250
rect -5659 14178 -5653 14212
rect -5619 14178 -5613 14212
rect -5659 14140 -5613 14178
rect -5659 14106 -5653 14140
rect -5619 14106 -5613 14140
rect -5659 14068 -5613 14106
rect -5659 14034 -5653 14068
rect -5619 14034 -5613 14068
rect -5659 13996 -5613 14034
rect -5659 13962 -5653 13996
rect -5619 13962 -5613 13996
rect -5659 13924 -5613 13962
rect -5659 13890 -5653 13924
rect -5619 13890 -5613 13924
rect -5659 13852 -5613 13890
rect -5659 13818 -5653 13852
rect -5619 13818 -5613 13852
rect -5659 13780 -5613 13818
rect -5659 13746 -5653 13780
rect -5619 13746 -5613 13780
rect -5659 13708 -5613 13746
rect -5659 13674 -5653 13708
rect -5619 13674 -5613 13708
rect -5659 13636 -5613 13674
rect -5659 13602 -5653 13636
rect -5619 13602 -5613 13636
rect -5659 13564 -5613 13602
rect -5659 13530 -5653 13564
rect -5619 13530 -5613 13564
rect -5659 13492 -5613 13530
rect -5659 13458 -5653 13492
rect -5619 13458 -5613 13492
rect -5659 13420 -5613 13458
rect -5659 13386 -5653 13420
rect -5619 13386 -5613 13420
rect -5659 13348 -5613 13386
rect -5659 13314 -5653 13348
rect -5619 13314 -5613 13348
rect -5659 13276 -5613 13314
rect -5659 13242 -5653 13276
rect -5619 13242 -5613 13276
rect -5659 13204 -5613 13242
rect -5659 13170 -5653 13204
rect -5619 13170 -5613 13204
rect -5659 13132 -5613 13170
rect -5401 14788 -5355 14835
rect -5401 14754 -5395 14788
rect -5361 14754 -5355 14788
rect -5401 14716 -5355 14754
rect -5401 14682 -5395 14716
rect -5361 14682 -5355 14716
rect -5401 14644 -5355 14682
rect -5401 14610 -5395 14644
rect -5361 14610 -5355 14644
rect -5401 14572 -5355 14610
rect -5401 14538 -5395 14572
rect -5361 14538 -5355 14572
rect -5401 14500 -5355 14538
rect -5401 14466 -5395 14500
rect -5361 14466 -5355 14500
rect -5401 14428 -5355 14466
rect -5401 14394 -5395 14428
rect -5361 14394 -5355 14428
rect -5401 14356 -5355 14394
rect -5401 14322 -5395 14356
rect -5361 14322 -5355 14356
rect -5401 14284 -5355 14322
rect -5401 14250 -5395 14284
rect -5361 14250 -5355 14284
rect -5401 14212 -5355 14250
rect -5401 14178 -5395 14212
rect -5361 14178 -5355 14212
rect -5401 14140 -5355 14178
rect -5401 14106 -5395 14140
rect -5361 14106 -5355 14140
rect -5401 14068 -5355 14106
rect -5401 14034 -5395 14068
rect -5361 14034 -5355 14068
rect -5401 13996 -5355 14034
rect -5401 13962 -5395 13996
rect -5361 13962 -5355 13996
rect -5401 13924 -5355 13962
rect -5401 13890 -5395 13924
rect -5361 13890 -5355 13924
rect -5401 13852 -5355 13890
rect -5401 13818 -5395 13852
rect -5361 13818 -5355 13852
rect -5401 13780 -5355 13818
rect -5401 13746 -5395 13780
rect -5361 13746 -5355 13780
rect -5401 13708 -5355 13746
rect -5401 13674 -5395 13708
rect -5361 13674 -5355 13708
rect -5401 13636 -5355 13674
rect -5401 13602 -5395 13636
rect -5361 13602 -5355 13636
rect -5401 13564 -5355 13602
rect -5401 13530 -5395 13564
rect -5361 13530 -5355 13564
rect -5401 13492 -5355 13530
rect -5401 13458 -5395 13492
rect -5361 13458 -5355 13492
rect -5401 13420 -5355 13458
rect -5401 13386 -5395 13420
rect -5361 13386 -5355 13420
rect -5401 13348 -5355 13386
rect -5401 13314 -5395 13348
rect -5361 13314 -5355 13348
rect -5401 13276 -5355 13314
rect -5401 13242 -5395 13276
rect -5361 13242 -5355 13276
rect -5401 13204 -5355 13242
rect -5401 13170 -5395 13204
rect -5361 13170 -5355 13204
rect -5401 13140 -5355 13170
rect -5143 14788 -5097 14835
rect -4885 14809 -4839 14835
rect -3949 14813 -3776 14851
rect -5143 14754 -5137 14788
rect -5103 14754 -5097 14788
rect -5143 14716 -5097 14754
rect -5143 14682 -5137 14716
rect -5103 14682 -5097 14716
rect -5143 14644 -5097 14682
rect -5143 14610 -5137 14644
rect -5103 14610 -5097 14644
rect -5143 14572 -5097 14610
rect -5143 14538 -5137 14572
rect -5103 14538 -5097 14572
rect -5143 14500 -5097 14538
rect -4946 14788 -4796 14809
rect -4946 14755 -4879 14788
rect -4946 14703 -4899 14755
rect -4845 14754 -4796 14788
rect -4847 14716 -4796 14754
rect -4946 14691 -4879 14703
rect -4946 14639 -4899 14691
rect -4845 14682 -4796 14716
rect -4847 14644 -4796 14682
rect -4946 14627 -4879 14639
rect -4946 14575 -4899 14627
rect -4845 14610 -4796 14644
rect -4847 14575 -4796 14610
rect -4946 14572 -4796 14575
rect -4946 14538 -4879 14572
rect -4845 14538 -4796 14572
rect -4946 14523 -4796 14538
rect -3949 14779 -3862 14813
rect -3828 14779 -3776 14813
rect 13044 14848 14036 14854
rect 13044 14814 13091 14848
rect 13125 14814 13163 14848
rect 13197 14814 13235 14848
rect 13269 14814 13307 14848
rect 13341 14814 13379 14848
rect 13413 14814 13451 14848
rect 13485 14814 13523 14848
rect 13557 14814 13595 14848
rect 13629 14814 13667 14848
rect 13701 14814 13739 14848
rect 13773 14814 13811 14848
rect 13845 14814 13883 14848
rect 13917 14814 13955 14848
rect 13989 14814 14036 14848
rect 13044 14808 14036 14814
rect 14102 14848 15094 14854
rect 14102 14814 14149 14848
rect 14183 14814 14221 14848
rect 14255 14814 14293 14848
rect 14327 14814 14365 14848
rect 14399 14814 14437 14848
rect 14471 14814 14509 14848
rect 14543 14814 14581 14848
rect 14615 14814 14653 14848
rect 14687 14814 14725 14848
rect 14759 14814 14797 14848
rect 14831 14814 14869 14848
rect 14903 14814 14941 14848
rect 14975 14814 15013 14848
rect 15047 14814 15094 14848
rect 14102 14808 15094 14814
rect 15614 14848 17171 14854
rect 15614 14814 15661 14848
rect 15695 14814 15733 14848
rect 15767 14814 15805 14848
rect 15839 14814 15877 14848
rect 15911 14814 15949 14848
rect 15983 14814 16021 14848
rect 16055 14814 16093 14848
rect 16127 14814 16165 14848
rect 16199 14814 16237 14848
rect 16271 14814 16309 14848
rect 16343 14814 16381 14848
rect 16415 14814 16453 14848
rect 16487 14814 16525 14848
rect 16559 14824 17171 14848
rect 17205 14824 17243 14858
rect 17277 14824 17315 14858
rect 17349 14824 17387 14858
rect 17421 14824 17459 14858
rect 17493 14824 17531 14858
rect 17565 14824 17603 14858
rect 17637 14824 17675 14858
rect 17709 14824 17747 14858
rect 17781 14824 17819 14858
rect 17853 14824 17891 14858
rect 17925 14824 17963 14858
rect 17997 14824 18035 14858
rect 18069 14824 18116 14858
rect 16559 14820 18116 14824
rect 16559 14814 16606 14820
rect 17124 14818 18116 14820
rect 18588 14842 19580 14848
rect 15614 14808 16606 14814
rect 18588 14808 18635 14842
rect 18669 14808 18707 14842
rect 18741 14808 18779 14842
rect 18813 14808 18851 14842
rect 18885 14808 18923 14842
rect 18957 14808 18995 14842
rect 19029 14808 19067 14842
rect 19101 14808 19139 14842
rect 19173 14808 19211 14842
rect 19245 14808 19283 14842
rect 19317 14808 19355 14842
rect 19389 14808 19427 14842
rect 19461 14808 19499 14842
rect 19533 14808 19580 14842
rect 18588 14802 19580 14808
rect -3949 14741 -3776 14779
rect -3949 14707 -3862 14741
rect -3828 14707 -3776 14741
rect -3949 14669 -3776 14707
rect -3949 14635 -3862 14669
rect -3828 14635 -3776 14669
rect -3949 14597 -3776 14635
rect -3949 14563 -3862 14597
rect -3828 14563 -3776 14597
rect -3949 14525 -3776 14563
rect -5143 14466 -5137 14500
rect -5103 14466 -5097 14500
rect -5143 14428 -5097 14466
rect -5143 14394 -5137 14428
rect -5103 14394 -5097 14428
rect -5143 14356 -5097 14394
rect -5143 14322 -5137 14356
rect -5103 14322 -5097 14356
rect -5143 14284 -5097 14322
rect -5143 14250 -5137 14284
rect -5103 14250 -5097 14284
rect -5143 14212 -5097 14250
rect -5143 14178 -5137 14212
rect -5103 14178 -5097 14212
rect -5143 14140 -5097 14178
rect -5143 14106 -5137 14140
rect -5103 14106 -5097 14140
rect -5143 14068 -5097 14106
rect -5143 14034 -5137 14068
rect -5103 14034 -5097 14068
rect -5143 13996 -5097 14034
rect -5143 13962 -5137 13996
rect -5103 13962 -5097 13996
rect -5143 13924 -5097 13962
rect -5143 13890 -5137 13924
rect -5103 13890 -5097 13924
rect -5143 13852 -5097 13890
rect -5143 13818 -5137 13852
rect -5103 13818 -5097 13852
rect -5143 13780 -5097 13818
rect -5143 13746 -5137 13780
rect -5103 13746 -5097 13780
rect -5143 13708 -5097 13746
rect -5143 13674 -5137 13708
rect -5103 13674 -5097 13708
rect -5143 13636 -5097 13674
rect -5143 13602 -5137 13636
rect -5103 13602 -5097 13636
rect -5143 13564 -5097 13602
rect -5143 13530 -5137 13564
rect -5103 13530 -5097 13564
rect -5143 13492 -5097 13530
rect -5143 13458 -5137 13492
rect -5103 13458 -5097 13492
rect -5143 13420 -5097 13458
rect -5143 13386 -5137 13420
rect -5103 13386 -5097 13420
rect -5143 13348 -5097 13386
rect -5143 13314 -5137 13348
rect -5103 13314 -5097 13348
rect -5143 13276 -5097 13314
rect -5143 13242 -5137 13276
rect -5103 13242 -5097 13276
rect -5143 13204 -5097 13242
rect -5143 13170 -5137 13204
rect -5103 13170 -5097 13204
rect -5659 13098 -5653 13132
rect -5619 13098 -5613 13132
rect -5659 13060 -5613 13098
rect -5659 13026 -5653 13060
rect -5619 13026 -5613 13060
rect -5659 12988 -5613 13026
rect -5659 12954 -5653 12988
rect -5619 12954 -5613 12988
rect -5659 12916 -5613 12954
rect -5659 12882 -5653 12916
rect -5619 12882 -5613 12916
rect -5659 12835 -5613 12882
rect -5451 13132 -5301 13140
rect -5451 13098 -5395 13132
rect -5361 13098 -5301 13132
rect -5451 13086 -5301 13098
rect -5451 13034 -5404 13086
rect -5352 13034 -5301 13086
rect -5451 13026 -5395 13034
rect -5361 13026 -5301 13034
rect -5451 13022 -5301 13026
rect -5451 12970 -5404 13022
rect -5352 12970 -5301 13022
rect -5451 12958 -5395 12970
rect -5361 12958 -5301 12970
rect -5451 12906 -5404 12958
rect -5352 12906 -5301 12958
rect -5451 12882 -5395 12906
rect -5361 12882 -5301 12906
rect -5451 12854 -5301 12882
rect -5143 13132 -5097 13170
rect -5143 13098 -5137 13132
rect -5103 13098 -5097 13132
rect -5143 13060 -5097 13098
rect -5143 13026 -5137 13060
rect -5103 13026 -5097 13060
rect -5143 12988 -5097 13026
rect -5143 12954 -5137 12988
rect -5103 12954 -5097 12988
rect -5143 12916 -5097 12954
rect -5143 12882 -5137 12916
rect -5103 12882 -5097 12916
rect -5401 12835 -5355 12854
rect -5143 12835 -5097 12882
rect -4885 14500 -4839 14523
rect -4885 14466 -4879 14500
rect -4845 14466 -4839 14500
rect -4885 14428 -4839 14466
rect -3949 14491 -3862 14525
rect -3828 14491 -3776 14525
rect -3949 14459 -3776 14491
rect 12988 14724 13034 14767
rect 12988 14690 12994 14724
rect 13028 14690 13034 14724
rect 12988 14652 13034 14690
rect 12988 14618 12994 14652
rect 13028 14618 13034 14652
rect 12988 14580 13034 14618
rect 12988 14546 12994 14580
rect 13028 14546 13034 14580
rect 12988 14508 13034 14546
rect 14046 14724 14092 14767
rect 14046 14690 14052 14724
rect 14086 14690 14092 14724
rect 14046 14652 14092 14690
rect 14046 14618 14052 14652
rect 14086 14618 14092 14652
rect 14046 14580 14092 14618
rect 14046 14546 14052 14580
rect 14086 14546 14092 14580
rect 14046 14530 14092 14546
rect 15104 14724 15150 14767
rect 15104 14690 15110 14724
rect 15144 14690 15150 14724
rect 15104 14652 15150 14690
rect 15104 14618 15110 14652
rect 15144 14618 15150 14652
rect 15104 14580 15150 14618
rect 15104 14546 15110 14580
rect 15144 14546 15150 14580
rect 12988 14474 12994 14508
rect 13028 14474 13034 14508
rect -4885 14394 -4879 14428
rect -4845 14394 -4839 14428
rect -4885 14356 -4839 14394
rect -4885 14322 -4879 14356
rect -4845 14322 -4839 14356
rect -4885 14284 -4839 14322
rect -4885 14250 -4879 14284
rect -4845 14250 -4839 14284
rect -4885 14212 -4839 14250
rect -4885 14178 -4879 14212
rect -4845 14178 -4839 14212
rect -4885 14140 -4839 14178
rect -4885 14106 -4879 14140
rect -4845 14106 -4839 14140
rect -4885 14068 -4839 14106
rect -4885 14034 -4879 14068
rect -4845 14034 -4839 14068
rect -4885 13996 -4839 14034
rect -4885 13962 -4879 13996
rect -4845 13962 -4839 13996
rect -4885 13924 -4839 13962
rect -4885 13890 -4879 13924
rect -4845 13890 -4839 13924
rect -4885 13852 -4839 13890
rect -4885 13818 -4879 13852
rect -4845 13818 -4839 13852
rect -4885 13780 -4839 13818
rect -4885 13746 -4879 13780
rect -4845 13746 -4839 13780
rect -4885 13708 -4839 13746
rect -4885 13674 -4879 13708
rect -4845 13674 -4839 13708
rect -4885 13636 -4839 13674
rect -4885 13602 -4879 13636
rect -4845 13602 -4839 13636
rect -4885 13564 -4839 13602
rect -4885 13530 -4879 13564
rect -4845 13530 -4839 13564
rect -4885 13492 -4839 13530
rect -4885 13458 -4879 13492
rect -4845 13458 -4839 13492
rect -4885 13420 -4839 13458
rect -4885 13386 -4879 13420
rect -4845 13386 -4839 13420
rect -4885 13348 -4839 13386
rect -4885 13314 -4879 13348
rect -4845 13314 -4839 13348
rect -4885 13276 -4839 13314
rect -4885 13242 -4879 13276
rect -4845 13242 -4839 13276
rect -4885 13204 -4839 13242
rect -4885 13170 -4879 13204
rect -4845 13170 -4839 13204
rect -4885 13132 -4839 13170
rect -4885 13098 -4879 13132
rect -4845 13098 -4839 13132
rect -4885 13060 -4839 13098
rect -4885 13026 -4879 13060
rect -4845 13026 -4839 13060
rect -4885 12988 -4839 13026
rect -4885 12954 -4879 12988
rect -4845 12954 -4839 12988
rect -4885 12916 -4839 12954
rect -4885 12882 -4879 12916
rect -4845 12882 -4839 12916
rect -4885 12835 -4839 12882
rect 12988 14436 13034 14474
rect 12988 14402 12994 14436
rect 13028 14402 13034 14436
rect 12988 14364 13034 14402
rect 12988 14330 12994 14364
rect 13028 14330 13034 14364
rect 12988 14292 13034 14330
rect 12988 14258 12994 14292
rect 13028 14258 13034 14292
rect 12988 14220 13034 14258
rect 12988 14186 12994 14220
rect 13028 14186 13034 14220
rect 12988 14148 13034 14186
rect 13932 14509 14212 14530
rect 13932 14201 13982 14509
rect 14162 14201 14212 14509
rect 13932 14186 14052 14201
rect 14086 14186 14212 14201
rect 13932 14180 14212 14186
rect 15104 14508 15150 14546
rect 15104 14474 15110 14508
rect 15144 14474 15150 14508
rect 15104 14436 15150 14474
rect 15104 14402 15110 14436
rect 15144 14402 15150 14436
rect 15104 14364 15150 14402
rect 15104 14330 15110 14364
rect 15144 14330 15150 14364
rect 15104 14292 15150 14330
rect 15104 14258 15110 14292
rect 15144 14258 15150 14292
rect 15104 14220 15150 14258
rect 15104 14186 15110 14220
rect 15144 14186 15150 14220
rect 12988 14114 12994 14148
rect 13028 14114 13034 14148
rect 12988 14076 13034 14114
rect 12988 14042 12994 14076
rect 13028 14042 13034 14076
rect 12988 14004 13034 14042
rect 12988 13970 12994 14004
rect 13028 13970 13034 14004
rect 12988 13932 13034 13970
rect 12988 13898 12994 13932
rect 13028 13898 13034 13932
rect 12988 13860 13034 13898
rect 12988 13826 12994 13860
rect 13028 13826 13034 13860
rect 12988 13788 13034 13826
rect 12988 13754 12994 13788
rect 13028 13754 13034 13788
rect 12988 13716 13034 13754
rect 12988 13682 12994 13716
rect 13028 13682 13034 13716
rect 12988 13644 13034 13682
rect 12988 13610 12994 13644
rect 13028 13610 13034 13644
rect 12988 13572 13034 13610
rect 12988 13538 12994 13572
rect 13028 13538 13034 13572
rect 12988 13500 13034 13538
rect 12988 13466 12994 13500
rect 13028 13466 13034 13500
rect 12988 13428 13034 13466
rect 12988 13394 12994 13428
rect 13028 13394 13034 13428
rect 12988 13356 13034 13394
rect 12988 13322 12994 13356
rect 13028 13322 13034 13356
rect 12988 13284 13034 13322
rect 12988 13250 12994 13284
rect 13028 13250 13034 13284
rect 12988 13212 13034 13250
rect 12988 13178 12994 13212
rect 13028 13178 13034 13212
rect 12988 13140 13034 13178
rect 12988 13106 12994 13140
rect 13028 13106 13034 13140
rect 12988 13068 13034 13106
rect 12988 13034 12994 13068
rect 13028 13034 13034 13068
rect 12988 12996 13034 13034
rect 12988 12962 12994 12996
rect 13028 12962 13034 12996
rect 12988 12924 13034 12962
rect 12988 12890 12994 12924
rect 13028 12890 13034 12924
rect -3939 12854 -3774 12875
rect -3939 12821 -3862 12854
rect -3828 12821 -3774 12854
rect -6872 12767 -6698 12787
rect -6872 12715 -6845 12767
rect -6793 12715 -6781 12767
rect -6729 12715 -6698 12767
rect -6872 12701 -6698 12715
rect -5382 12672 -4756 12676
rect -7671 12626 -4756 12672
rect -7671 12562 -5315 12626
rect -7671 12560 -6310 12562
rect -7671 12552 -6550 12560
rect -7671 12518 -7339 12552
rect -7305 12526 -6550 12552
rect -6516 12528 -6310 12560
rect -6276 12557 -5315 12562
rect -6276 12528 -5531 12557
rect -6516 12526 -5531 12528
rect -7305 12523 -5531 12526
rect -5497 12523 -5315 12557
rect -7305 12518 -5315 12523
rect -7671 12490 -5315 12518
rect -7671 12488 -6310 12490
rect -7671 12480 -6550 12488
rect -7671 12446 -7339 12480
rect -7305 12454 -6550 12480
rect -6516 12456 -6310 12488
rect -6276 12485 -5315 12490
rect -6276 12456 -5531 12485
rect -6516 12454 -5531 12456
rect -7305 12451 -5531 12454
rect -5497 12451 -5315 12485
rect -7305 12446 -5315 12451
rect -4815 12446 -4756 12626
rect -7671 12402 -4756 12446
rect -3939 12449 -3918 12821
rect -3802 12449 -3774 12821
rect -3939 12404 -3774 12449
rect 12988 12852 13034 12890
rect 12988 12818 12994 12852
rect 13028 12818 13034 12852
rect 12988 12780 13034 12818
rect 12988 12746 12994 12780
rect 13028 12746 13034 12780
rect 12988 12708 13034 12746
rect 12988 12674 12994 12708
rect 13028 12674 13034 12708
rect 12988 12636 13034 12674
rect 12988 12602 12994 12636
rect 13028 12602 13034 12636
rect 12988 12564 13034 12602
rect 12988 12530 12994 12564
rect 13028 12530 13034 12564
rect 12988 12492 13034 12530
rect 12988 12458 12994 12492
rect 13028 12458 13034 12492
rect 12988 12420 13034 12458
rect -5382 12400 -4756 12402
rect 12988 12386 12994 12420
rect 13028 12386 13034 12420
rect 12988 12348 13034 12386
rect 12988 12314 12994 12348
rect 13028 12314 13034 12348
rect 12988 12276 13034 12314
rect 12988 12242 12994 12276
rect 13028 12242 13034 12276
rect 12988 12204 13034 12242
rect 12988 12170 12994 12204
rect 13028 12170 13034 12204
rect 12988 12132 13034 12170
rect 12988 12100 12994 12132
rect 12982 12098 12994 12100
rect 13028 12100 13034 12132
rect 14046 14148 14092 14180
rect 14046 14114 14052 14148
rect 14086 14114 14092 14148
rect 14046 14076 14092 14114
rect 14046 14042 14052 14076
rect 14086 14042 14092 14076
rect 14046 14004 14092 14042
rect 14046 13970 14052 14004
rect 14086 13970 14092 14004
rect 14046 13932 14092 13970
rect 14046 13898 14052 13932
rect 14086 13898 14092 13932
rect 14046 13860 14092 13898
rect 14046 13826 14052 13860
rect 14086 13826 14092 13860
rect 14046 13788 14092 13826
rect 14046 13754 14052 13788
rect 14086 13754 14092 13788
rect 14046 13716 14092 13754
rect 14046 13682 14052 13716
rect 14086 13682 14092 13716
rect 14046 13644 14092 13682
rect 14046 13610 14052 13644
rect 14086 13610 14092 13644
rect 14046 13572 14092 13610
rect 14046 13538 14052 13572
rect 14086 13538 14092 13572
rect 14046 13500 14092 13538
rect 14046 13466 14052 13500
rect 14086 13466 14092 13500
rect 14046 13428 14092 13466
rect 14046 13394 14052 13428
rect 14086 13394 14092 13428
rect 14046 13356 14092 13394
rect 14046 13322 14052 13356
rect 14086 13322 14092 13356
rect 14046 13284 14092 13322
rect 14046 13250 14052 13284
rect 14086 13250 14092 13284
rect 14046 13212 14092 13250
rect 14046 13178 14052 13212
rect 14086 13178 14092 13212
rect 14046 13140 14092 13178
rect 14046 13106 14052 13140
rect 14086 13106 14092 13140
rect 14046 13068 14092 13106
rect 14046 13034 14052 13068
rect 14086 13034 14092 13068
rect 14046 12996 14092 13034
rect 14046 12962 14052 12996
rect 14086 12962 14092 12996
rect 14046 12924 14092 12962
rect 14046 12890 14052 12924
rect 14086 12890 14092 12924
rect 14046 12852 14092 12890
rect 14046 12818 14052 12852
rect 14086 12818 14092 12852
rect 14046 12780 14092 12818
rect 14046 12746 14052 12780
rect 14086 12746 14092 12780
rect 14046 12708 14092 12746
rect 14046 12674 14052 12708
rect 14086 12674 14092 12708
rect 14046 12636 14092 12674
rect 14046 12602 14052 12636
rect 14086 12602 14092 12636
rect 14046 12564 14092 12602
rect 14046 12530 14052 12564
rect 14086 12530 14092 12564
rect 14046 12492 14092 12530
rect 14046 12458 14052 12492
rect 14086 12458 14092 12492
rect 14046 12420 14092 12458
rect 14046 12386 14052 12420
rect 14086 12386 14092 12420
rect 14046 12348 14092 12386
rect 14046 12314 14052 12348
rect 14086 12314 14092 12348
rect 14046 12276 14092 12314
rect 14046 12242 14052 12276
rect 14086 12242 14092 12276
rect 14046 12204 14092 12242
rect 14046 12170 14052 12204
rect 14086 12170 14092 12204
rect 14046 12132 14092 12170
rect 13028 12098 13162 12100
rect 12982 12060 13162 12098
rect 12982 12026 12994 12060
rect 13028 12052 13162 12060
rect 12982 11988 13014 12026
rect 12982 11954 12994 11988
rect 12982 11916 13014 11954
rect 12982 11882 12994 11916
rect 12982 11844 13014 11882
rect 12982 11810 12994 11844
rect 12982 11808 13014 11810
rect 13130 11808 13162 12052
rect 12982 11770 13162 11808
rect 14046 12098 14052 12132
rect 14086 12098 14092 12132
rect 15104 14148 15150 14186
rect 15104 14114 15110 14148
rect 15144 14114 15150 14148
rect 15104 14076 15150 14114
rect 15104 14042 15110 14076
rect 15144 14042 15150 14076
rect 15104 14004 15150 14042
rect 15104 13970 15110 14004
rect 15144 13970 15150 14004
rect 15104 13932 15150 13970
rect 15104 13898 15110 13932
rect 15144 13898 15150 13932
rect 15104 13860 15150 13898
rect 15104 13826 15110 13860
rect 15144 13826 15150 13860
rect 15104 13788 15150 13826
rect 15104 13754 15110 13788
rect 15144 13754 15150 13788
rect 15104 13716 15150 13754
rect 15104 13682 15110 13716
rect 15144 13682 15150 13716
rect 15104 13644 15150 13682
rect 15104 13610 15110 13644
rect 15144 13610 15150 13644
rect 15104 13572 15150 13610
rect 15104 13538 15110 13572
rect 15144 13538 15150 13572
rect 15104 13500 15150 13538
rect 15104 13466 15110 13500
rect 15144 13466 15150 13500
rect 15104 13428 15150 13466
rect 15104 13394 15110 13428
rect 15144 13394 15150 13428
rect 15104 13356 15150 13394
rect 15104 13322 15110 13356
rect 15144 13322 15150 13356
rect 15104 13284 15150 13322
rect 15104 13250 15110 13284
rect 15144 13250 15150 13284
rect 15104 13212 15150 13250
rect 15104 13178 15110 13212
rect 15144 13178 15150 13212
rect 15104 13140 15150 13178
rect 15104 13106 15110 13140
rect 15144 13106 15150 13140
rect 15104 13068 15150 13106
rect 15104 13034 15110 13068
rect 15144 13034 15150 13068
rect 15104 12996 15150 13034
rect 15104 12962 15110 12996
rect 15144 12962 15150 12996
rect 15104 12924 15150 12962
rect 15104 12890 15110 12924
rect 15144 12890 15150 12924
rect 15104 12852 15150 12890
rect 15104 12818 15110 12852
rect 15144 12818 15150 12852
rect 15104 12780 15150 12818
rect 15104 12746 15110 12780
rect 15144 12746 15150 12780
rect 15104 12708 15150 12746
rect 15104 12674 15110 12708
rect 15144 12674 15150 12708
rect 15104 12636 15150 12674
rect 15104 12602 15110 12636
rect 15144 12602 15150 12636
rect 15104 12564 15150 12602
rect 15104 12530 15110 12564
rect 15144 12530 15150 12564
rect 15104 12492 15150 12530
rect 15104 12458 15110 12492
rect 15144 12458 15150 12492
rect 15104 12420 15150 12458
rect 15104 12386 15110 12420
rect 15144 12386 15150 12420
rect 15104 12348 15150 12386
rect 15104 12314 15110 12348
rect 15144 12314 15150 12348
rect 15104 12276 15150 12314
rect 15104 12242 15110 12276
rect 15144 12242 15150 12276
rect 15104 12204 15150 12242
rect 15104 12170 15110 12204
rect 15144 12170 15150 12204
rect 15104 12132 15150 12170
rect 15104 12100 15110 12132
rect 14046 12060 14092 12098
rect 14046 12026 14052 12060
rect 14086 12026 14092 12060
rect 14046 11988 14092 12026
rect 14046 11954 14052 11988
rect 14086 11954 14092 11988
rect 14046 11916 14092 11954
rect 14046 11882 14052 11916
rect 14086 11882 14092 11916
rect 14046 11844 14092 11882
rect 14046 11810 14052 11844
rect 14086 11810 14092 11844
rect 12988 11767 13034 11770
rect 14046 11767 14092 11810
rect 14972 12098 15110 12100
rect 15144 12098 15150 12132
rect 14972 12060 15150 12098
rect 14972 12052 15110 12060
rect 14972 11808 14999 12052
rect 15144 12026 15150 12060
rect 15115 11988 15150 12026
rect 15144 11954 15150 11988
rect 15115 11916 15150 11954
rect 15144 11882 15150 11916
rect 15115 11844 15150 11882
rect 15144 11810 15150 11844
rect 15115 11808 15150 11810
rect 14972 11770 15150 11808
rect 15104 11767 15150 11770
rect 15558 14724 15604 14767
rect 15558 14690 15564 14724
rect 15598 14690 15604 14724
rect 15558 14652 15604 14690
rect 15558 14618 15564 14652
rect 15598 14618 15604 14652
rect 15558 14580 15604 14618
rect 15558 14546 15564 14580
rect 15598 14546 15604 14580
rect 15558 14530 15604 14546
rect 16616 14724 16662 14767
rect 16616 14690 16622 14724
rect 16656 14690 16662 14724
rect 16616 14652 16662 14690
rect 16616 14618 16622 14652
rect 16656 14618 16662 14652
rect 16616 14580 16662 14618
rect 16616 14546 16622 14580
rect 16656 14546 16662 14580
rect 15558 14509 15772 14530
rect 15558 14508 15609 14509
rect 15558 14474 15564 14508
rect 15598 14474 15609 14508
rect 15558 14436 15609 14474
rect 15558 14402 15564 14436
rect 15598 14402 15609 14436
rect 15558 14364 15609 14402
rect 15558 14330 15564 14364
rect 15598 14330 15609 14364
rect 15558 14292 15609 14330
rect 15558 14258 15564 14292
rect 15598 14258 15609 14292
rect 15558 14220 15609 14258
rect 15558 14186 15564 14220
rect 15598 14201 15609 14220
rect 15725 14201 15772 14509
rect 15598 14186 15772 14201
rect 15558 14180 15772 14186
rect 16616 14508 16662 14546
rect 16616 14474 16622 14508
rect 16656 14474 16662 14508
rect 16616 14436 16662 14474
rect 16616 14402 16622 14436
rect 16656 14402 16662 14436
rect 16616 14364 16662 14402
rect 16616 14330 16622 14364
rect 16656 14330 16662 14364
rect 16616 14292 16662 14330
rect 16616 14258 16622 14292
rect 16656 14258 16662 14292
rect 16616 14220 16662 14258
rect 16616 14186 16622 14220
rect 16656 14186 16662 14220
rect 15558 14148 15604 14180
rect 15558 14114 15564 14148
rect 15598 14114 15604 14148
rect 15558 14076 15604 14114
rect 15558 14042 15564 14076
rect 15598 14042 15604 14076
rect 15558 14004 15604 14042
rect 15558 13970 15564 14004
rect 15598 13970 15604 14004
rect 15558 13932 15604 13970
rect 15558 13898 15564 13932
rect 15598 13898 15604 13932
rect 15558 13860 15604 13898
rect 15558 13826 15564 13860
rect 15598 13826 15604 13860
rect 15558 13788 15604 13826
rect 15558 13754 15564 13788
rect 15598 13754 15604 13788
rect 15558 13716 15604 13754
rect 15558 13682 15564 13716
rect 15598 13682 15604 13716
rect 15558 13644 15604 13682
rect 15558 13610 15564 13644
rect 15598 13610 15604 13644
rect 15558 13572 15604 13610
rect 15558 13538 15564 13572
rect 15598 13538 15604 13572
rect 15558 13500 15604 13538
rect 15558 13466 15564 13500
rect 15598 13466 15604 13500
rect 15558 13428 15604 13466
rect 15558 13394 15564 13428
rect 15598 13394 15604 13428
rect 15558 13356 15604 13394
rect 15558 13322 15564 13356
rect 15598 13322 15604 13356
rect 15558 13284 15604 13322
rect 15558 13250 15564 13284
rect 15598 13250 15604 13284
rect 15558 13212 15604 13250
rect 15558 13178 15564 13212
rect 15598 13178 15604 13212
rect 15558 13140 15604 13178
rect 15558 13106 15564 13140
rect 15598 13106 15604 13140
rect 15558 13068 15604 13106
rect 15558 13034 15564 13068
rect 15598 13034 15604 13068
rect 15558 12996 15604 13034
rect 15558 12962 15564 12996
rect 15598 12962 15604 12996
rect 15558 12924 15604 12962
rect 15558 12890 15564 12924
rect 15598 12890 15604 12924
rect 15558 12852 15604 12890
rect 15558 12818 15564 12852
rect 15598 12818 15604 12852
rect 15558 12780 15604 12818
rect 15558 12746 15564 12780
rect 15598 12746 15604 12780
rect 15558 12708 15604 12746
rect 15558 12674 15564 12708
rect 15598 12674 15604 12708
rect 15558 12636 15604 12674
rect 15558 12602 15564 12636
rect 15598 12602 15604 12636
rect 15558 12564 15604 12602
rect 15558 12530 15564 12564
rect 15598 12530 15604 12564
rect 15558 12492 15604 12530
rect 15558 12458 15564 12492
rect 15598 12458 15604 12492
rect 15558 12420 15604 12458
rect 15558 12386 15564 12420
rect 15598 12386 15604 12420
rect 15558 12348 15604 12386
rect 15558 12314 15564 12348
rect 15598 12314 15604 12348
rect 15558 12276 15604 12314
rect 15558 12242 15564 12276
rect 15598 12242 15604 12276
rect 15558 12204 15604 12242
rect 15558 12170 15564 12204
rect 15598 12170 15604 12204
rect 15558 12132 15604 12170
rect 15558 12098 15564 12132
rect 15598 12098 15604 12132
rect 15558 12060 15604 12098
rect 15558 12026 15564 12060
rect 15598 12026 15604 12060
rect 15558 11988 15604 12026
rect 15558 11954 15564 11988
rect 15598 11954 15604 11988
rect 15558 11916 15604 11954
rect 15558 11882 15564 11916
rect 15598 11882 15604 11916
rect 15558 11844 15604 11882
rect 15558 11810 15564 11844
rect 15598 11810 15604 11844
rect 15558 11767 15604 11810
rect 16616 14148 16662 14186
rect 16616 14114 16622 14148
rect 16656 14114 16662 14148
rect 16616 14076 16662 14114
rect 16616 14042 16622 14076
rect 16656 14042 16662 14076
rect 16616 14004 16662 14042
rect 16616 13970 16622 14004
rect 16656 13970 16662 14004
rect 16616 13932 16662 13970
rect 16616 13898 16622 13932
rect 16656 13898 16662 13932
rect 16616 13860 16662 13898
rect 16616 13826 16622 13860
rect 16656 13826 16662 13860
rect 16616 13788 16662 13826
rect 16616 13754 16622 13788
rect 16656 13754 16662 13788
rect 16616 13716 16662 13754
rect 16616 13682 16622 13716
rect 16656 13682 16662 13716
rect 16616 13644 16662 13682
rect 16616 13610 16622 13644
rect 16656 13610 16662 13644
rect 16616 13572 16662 13610
rect 16616 13538 16622 13572
rect 16656 13538 16662 13572
rect 16616 13500 16662 13538
rect 16616 13466 16622 13500
rect 16656 13466 16662 13500
rect 16616 13428 16662 13466
rect 16616 13394 16622 13428
rect 16656 13394 16662 13428
rect 16616 13356 16662 13394
rect 16616 13322 16622 13356
rect 16656 13322 16662 13356
rect 16616 13284 16662 13322
rect 16616 13250 16622 13284
rect 16656 13250 16662 13284
rect 16616 13212 16662 13250
rect 16616 13178 16622 13212
rect 16656 13178 16662 13212
rect 16616 13140 16662 13178
rect 16616 13106 16622 13140
rect 16656 13106 16662 13140
rect 16616 13068 16662 13106
rect 16616 13034 16622 13068
rect 16656 13034 16662 13068
rect 16616 12996 16662 13034
rect 16616 12962 16622 12996
rect 16656 12962 16662 12996
rect 16616 12924 16662 12962
rect 16616 12890 16622 12924
rect 16656 12890 16662 12924
rect 16616 12852 16662 12890
rect 16616 12818 16622 12852
rect 16656 12818 16662 12852
rect 16616 12780 16662 12818
rect 16616 12746 16622 12780
rect 16656 12746 16662 12780
rect 16616 12708 16662 12746
rect 16616 12674 16622 12708
rect 16656 12674 16662 12708
rect 16616 12636 16662 12674
rect 16616 12602 16622 12636
rect 16656 12602 16662 12636
rect 16616 12564 16662 12602
rect 16616 12530 16622 12564
rect 16656 12530 16662 12564
rect 16616 12492 16662 12530
rect 16616 12458 16622 12492
rect 16656 12458 16662 12492
rect 16616 12420 16662 12458
rect 16616 12386 16622 12420
rect 16656 12386 16662 12420
rect 17068 14734 17114 14777
rect 17068 14700 17074 14734
rect 17108 14700 17114 14734
rect 17068 14662 17114 14700
rect 17068 14628 17074 14662
rect 17108 14628 17114 14662
rect 17068 14590 17114 14628
rect 17068 14556 17074 14590
rect 17108 14556 17114 14590
rect 17068 14518 17114 14556
rect 17068 14484 17074 14518
rect 17108 14484 17114 14518
rect 17068 14446 17114 14484
rect 17068 14412 17074 14446
rect 17108 14412 17114 14446
rect 17068 14374 17114 14412
rect 17068 14340 17074 14374
rect 17108 14340 17114 14374
rect 17068 14302 17114 14340
rect 17068 14268 17074 14302
rect 17108 14268 17114 14302
rect 17068 14230 17114 14268
rect 17068 14196 17074 14230
rect 17108 14196 17114 14230
rect 17068 14158 17114 14196
rect 17068 14124 17074 14158
rect 17108 14124 17114 14158
rect 17068 14086 17114 14124
rect 17068 14052 17074 14086
rect 17108 14052 17114 14086
rect 17068 14014 17114 14052
rect 17068 13980 17074 14014
rect 17108 13980 17114 14014
rect 17068 13942 17114 13980
rect 17068 13908 17074 13942
rect 17108 13908 17114 13942
rect 17068 13870 17114 13908
rect 17068 13836 17074 13870
rect 17108 13836 17114 13870
rect 17068 13798 17114 13836
rect 17068 13764 17074 13798
rect 17108 13764 17114 13798
rect 17068 13726 17114 13764
rect 17068 13692 17074 13726
rect 17108 13692 17114 13726
rect 17068 13654 17114 13692
rect 17068 13620 17074 13654
rect 17108 13620 17114 13654
rect 17068 13582 17114 13620
rect 17068 13548 17074 13582
rect 17108 13548 17114 13582
rect 17068 13510 17114 13548
rect 17068 13476 17074 13510
rect 17108 13476 17114 13510
rect 17068 13438 17114 13476
rect 17068 13404 17074 13438
rect 17108 13404 17114 13438
rect 17068 13366 17114 13404
rect 17068 13332 17074 13366
rect 17108 13332 17114 13366
rect 17068 13294 17114 13332
rect 17068 13260 17074 13294
rect 17108 13260 17114 13294
rect 17068 13222 17114 13260
rect 17068 13188 17074 13222
rect 17108 13188 17114 13222
rect 17068 13150 17114 13188
rect 17068 13116 17074 13150
rect 17108 13116 17114 13150
rect 17068 13078 17114 13116
rect 17068 13044 17074 13078
rect 17108 13044 17114 13078
rect 17068 13006 17114 13044
rect 17068 12972 17074 13006
rect 17108 12972 17114 13006
rect 17068 12934 17114 12972
rect 17068 12900 17074 12934
rect 17108 12900 17114 12934
rect 17068 12862 17114 12900
rect 17068 12828 17074 12862
rect 17108 12828 17114 12862
rect 17068 12790 17114 12828
rect 17068 12756 17074 12790
rect 17108 12756 17114 12790
rect 17068 12718 17114 12756
rect 17068 12684 17074 12718
rect 17108 12684 17114 12718
rect 17068 12646 17114 12684
rect 17068 12612 17074 12646
rect 17108 12612 17114 12646
rect 17068 12574 17114 12612
rect 17068 12540 17074 12574
rect 17108 12540 17114 12574
rect 17068 12502 17114 12540
rect 17068 12468 17074 12502
rect 17108 12468 17114 12502
rect 17068 12430 17114 12468
rect 17068 12400 17074 12430
rect 16616 12348 16662 12386
rect 16616 12314 16622 12348
rect 16656 12314 16662 12348
rect 16616 12276 16662 12314
rect 16616 12242 16622 12276
rect 16656 12242 16662 12276
rect 16616 12204 16662 12242
rect 16616 12170 16622 12204
rect 16656 12170 16662 12204
rect 16616 12132 16662 12170
rect 16616 12098 16622 12132
rect 16656 12098 16662 12132
rect 16616 12060 16662 12098
rect 16616 12026 16622 12060
rect 16656 12026 16662 12060
rect 16616 11988 16662 12026
rect 16616 11954 16622 11988
rect 16656 11954 16662 11988
rect 16616 11916 16662 11954
rect 17062 12396 17074 12400
rect 17108 12400 17114 12430
rect 18126 14734 18172 14777
rect 18126 14700 18132 14734
rect 18166 14700 18172 14734
rect 18126 14662 18172 14700
rect 18126 14628 18132 14662
rect 18166 14628 18172 14662
rect 18126 14590 18172 14628
rect 18126 14556 18132 14590
rect 18166 14556 18172 14590
rect 18126 14518 18172 14556
rect 18126 14484 18132 14518
rect 18166 14484 18172 14518
rect 18126 14446 18172 14484
rect 18126 14412 18132 14446
rect 18166 14412 18172 14446
rect 18126 14374 18172 14412
rect 18126 14340 18132 14374
rect 18166 14340 18172 14374
rect 18126 14302 18172 14340
rect 18126 14268 18132 14302
rect 18166 14268 18172 14302
rect 18126 14230 18172 14268
rect 18126 14196 18132 14230
rect 18166 14196 18172 14230
rect 18126 14158 18172 14196
rect 18126 14124 18132 14158
rect 18166 14124 18172 14158
rect 18126 14086 18172 14124
rect 18126 14052 18132 14086
rect 18166 14052 18172 14086
rect 18126 14014 18172 14052
rect 18126 13980 18132 14014
rect 18166 13980 18172 14014
rect 18126 13942 18172 13980
rect 18126 13908 18132 13942
rect 18166 13908 18172 13942
rect 18126 13870 18172 13908
rect 18126 13836 18132 13870
rect 18166 13836 18172 13870
rect 18126 13798 18172 13836
rect 18126 13764 18132 13798
rect 18166 13764 18172 13798
rect 18126 13726 18172 13764
rect 18126 13692 18132 13726
rect 18166 13692 18172 13726
rect 18126 13654 18172 13692
rect 18126 13620 18132 13654
rect 18166 13620 18172 13654
rect 18126 13582 18172 13620
rect 18126 13548 18132 13582
rect 18166 13548 18172 13582
rect 18126 13510 18172 13548
rect 18126 13476 18132 13510
rect 18166 13476 18172 13510
rect 18126 13438 18172 13476
rect 18126 13404 18132 13438
rect 18166 13404 18172 13438
rect 18126 13366 18172 13404
rect 18126 13332 18132 13366
rect 18166 13332 18172 13366
rect 18126 13294 18172 13332
rect 18126 13260 18132 13294
rect 18166 13260 18172 13294
rect 18126 13222 18172 13260
rect 18126 13188 18132 13222
rect 18166 13188 18172 13222
rect 18126 13150 18172 13188
rect 18126 13116 18132 13150
rect 18166 13116 18172 13150
rect 18126 13078 18172 13116
rect 18126 13044 18132 13078
rect 18166 13044 18172 13078
rect 18126 13006 18172 13044
rect 18126 12972 18132 13006
rect 18166 12972 18172 13006
rect 18126 12934 18172 12972
rect 18126 12900 18132 12934
rect 18166 12900 18172 12934
rect 18126 12862 18172 12900
rect 18126 12828 18132 12862
rect 18166 12828 18172 12862
rect 18126 12790 18172 12828
rect 18126 12756 18132 12790
rect 18166 12756 18172 12790
rect 18126 12718 18172 12756
rect 18126 12684 18132 12718
rect 18166 12684 18172 12718
rect 18126 12646 18172 12684
rect 18126 12612 18132 12646
rect 18166 12612 18172 12646
rect 18126 12574 18172 12612
rect 18126 12540 18132 12574
rect 18166 12540 18172 12574
rect 18126 12502 18172 12540
rect 18126 12468 18132 12502
rect 18166 12468 18172 12502
rect 18126 12430 18172 12468
rect 17108 12396 17262 12400
rect 17062 12358 17262 12396
rect 17062 12324 17074 12358
rect 17108 12351 17262 12358
rect 17062 12286 17104 12324
rect 17062 12252 17074 12286
rect 17062 12214 17104 12252
rect 17062 12180 17074 12214
rect 17062 12142 17104 12180
rect 17062 12108 17074 12142
rect 17062 12070 17104 12108
rect 17062 12036 17074 12070
rect 17062 11998 17104 12036
rect 17062 11964 17074 11998
rect 17220 11979 17262 12351
rect 17108 11964 17262 11979
rect 17062 11930 17262 11964
rect 18126 12396 18132 12430
rect 18166 12396 18172 12430
rect 18126 12358 18172 12396
rect 18126 12324 18132 12358
rect 18166 12324 18172 12358
rect 18126 12286 18172 12324
rect 18126 12252 18132 12286
rect 18166 12252 18172 12286
rect 18126 12214 18172 12252
rect 18126 12180 18132 12214
rect 18166 12180 18172 12214
rect 18126 12142 18172 12180
rect 18532 14718 18578 14761
rect 18532 14684 18538 14718
rect 18572 14684 18578 14718
rect 18532 14646 18578 14684
rect 18532 14612 18538 14646
rect 18572 14612 18578 14646
rect 18532 14574 18578 14612
rect 18532 14540 18538 14574
rect 18572 14540 18578 14574
rect 18532 14502 18578 14540
rect 18532 14468 18538 14502
rect 18572 14468 18578 14502
rect 18532 14430 18578 14468
rect 18532 14396 18538 14430
rect 18572 14396 18578 14430
rect 18532 14358 18578 14396
rect 18532 14324 18538 14358
rect 18572 14324 18578 14358
rect 18532 14286 18578 14324
rect 18532 14252 18538 14286
rect 18572 14252 18578 14286
rect 18532 14214 18578 14252
rect 18532 14180 18538 14214
rect 18572 14180 18578 14214
rect 18532 14142 18578 14180
rect 18532 14108 18538 14142
rect 18572 14108 18578 14142
rect 18532 14070 18578 14108
rect 18532 14036 18538 14070
rect 18572 14036 18578 14070
rect 18532 13998 18578 14036
rect 18532 13964 18538 13998
rect 18572 13964 18578 13998
rect 18532 13926 18578 13964
rect 18532 13892 18538 13926
rect 18572 13892 18578 13926
rect 18532 13854 18578 13892
rect 18532 13820 18538 13854
rect 18572 13820 18578 13854
rect 18532 13782 18578 13820
rect 18532 13748 18538 13782
rect 18572 13748 18578 13782
rect 18532 13710 18578 13748
rect 18532 13676 18538 13710
rect 18572 13676 18578 13710
rect 18532 13638 18578 13676
rect 18532 13604 18538 13638
rect 18572 13604 18578 13638
rect 18532 13566 18578 13604
rect 18532 13532 18538 13566
rect 18572 13532 18578 13566
rect 18532 13494 18578 13532
rect 18532 13460 18538 13494
rect 18572 13460 18578 13494
rect 18532 13422 18578 13460
rect 18532 13388 18538 13422
rect 18572 13388 18578 13422
rect 18532 13350 18578 13388
rect 18532 13316 18538 13350
rect 18572 13316 18578 13350
rect 18532 13278 18578 13316
rect 18532 13244 18538 13278
rect 18572 13244 18578 13278
rect 18532 13206 18578 13244
rect 18532 13172 18538 13206
rect 18572 13172 18578 13206
rect 18532 13134 18578 13172
rect 18532 13100 18538 13134
rect 18572 13100 18578 13134
rect 18532 13062 18578 13100
rect 18532 13028 18538 13062
rect 18572 13028 18578 13062
rect 18532 12990 18578 13028
rect 18532 12956 18538 12990
rect 18572 12956 18578 12990
rect 18532 12918 18578 12956
rect 18532 12884 18538 12918
rect 18572 12884 18578 12918
rect 18532 12846 18578 12884
rect 18532 12812 18538 12846
rect 18572 12812 18578 12846
rect 18532 12774 18578 12812
rect 18532 12740 18538 12774
rect 18572 12740 18578 12774
rect 18532 12702 18578 12740
rect 18532 12668 18538 12702
rect 18572 12668 18578 12702
rect 18532 12630 18578 12668
rect 18532 12596 18538 12630
rect 18572 12596 18578 12630
rect 18532 12558 18578 12596
rect 18532 12524 18538 12558
rect 18572 12524 18578 12558
rect 18532 12486 18578 12524
rect 18532 12452 18538 12486
rect 18572 12452 18578 12486
rect 18532 12414 18578 12452
rect 18532 12380 18538 12414
rect 18572 12380 18578 12414
rect 18532 12342 18578 12380
rect 18532 12308 18538 12342
rect 18572 12308 18578 12342
rect 18532 12270 18578 12308
rect 18532 12236 18538 12270
rect 18572 12236 18578 12270
rect 18532 12198 18578 12236
rect 18532 12164 18538 12198
rect 18572 12164 18578 12198
rect 18532 12154 18578 12164
rect 19590 14718 19636 14761
rect 19590 14684 19596 14718
rect 19630 14684 19636 14718
rect 19590 14646 19636 14684
rect 19590 14612 19596 14646
rect 19630 14612 19636 14646
rect 19590 14574 19636 14612
rect 19590 14540 19596 14574
rect 19630 14540 19636 14574
rect 19590 14502 19636 14540
rect 19590 14468 19596 14502
rect 19630 14468 19636 14502
rect 19590 14430 19636 14468
rect 19590 14396 19596 14430
rect 19630 14396 19636 14430
rect 19590 14358 19636 14396
rect 19590 14324 19596 14358
rect 19630 14324 19636 14358
rect 19590 14286 19636 14324
rect 19590 14252 19596 14286
rect 19630 14252 19636 14286
rect 19590 14214 19636 14252
rect 19590 14180 19596 14214
rect 19630 14180 19636 14214
rect 19590 14142 19636 14180
rect 19590 14108 19596 14142
rect 19630 14108 19636 14142
rect 19590 14070 19636 14108
rect 19590 14036 19596 14070
rect 19630 14036 19636 14070
rect 20522 14450 20572 14464
rect 20522 14416 20530 14450
rect 20564 14416 20572 14450
rect 20522 14378 20572 14416
rect 20522 14344 20530 14378
rect 20564 14344 20572 14378
rect 20522 14306 20572 14344
rect 20522 14272 20530 14306
rect 20564 14272 20572 14306
rect 20522 14234 20572 14272
rect 20522 14200 20530 14234
rect 20564 14200 20572 14234
rect 20522 14162 20572 14200
rect 20522 14128 20530 14162
rect 20564 14128 20572 14162
rect 20522 14090 20572 14128
rect 20522 14056 20530 14090
rect 20564 14056 20572 14090
rect 20522 14043 20572 14056
rect 20832 14450 20900 14468
rect 20832 14416 20848 14450
rect 20882 14416 20900 14450
rect 20832 14378 20900 14416
rect 20832 14344 20848 14378
rect 20882 14344 20900 14378
rect 20832 14306 20900 14344
rect 20832 14272 20848 14306
rect 20882 14272 20900 14306
rect 20832 14234 20900 14272
rect 20832 14200 20848 14234
rect 20882 14200 20900 14234
rect 20832 14162 20900 14200
rect 20832 14128 20848 14162
rect 20882 14128 20900 14162
rect 20832 14090 20900 14128
rect 20832 14056 20848 14090
rect 20882 14056 20900 14090
rect 19590 13998 19636 14036
rect 19590 13964 19596 13998
rect 19630 13964 19636 13998
rect 19590 13926 19636 13964
rect 19590 13892 19596 13926
rect 19630 13892 19636 13926
rect 19590 13854 19636 13892
rect 19590 13820 19596 13854
rect 19630 13820 19636 13854
rect 19590 13782 19636 13820
rect 19590 13748 19596 13782
rect 19630 13748 19636 13782
rect 19590 13710 19636 13748
rect 19590 13676 19596 13710
rect 19630 13676 19636 13710
rect 19590 13638 19636 13676
rect 19590 13604 19596 13638
rect 19630 13604 19636 13638
rect 19590 13566 19636 13604
rect 19590 13532 19596 13566
rect 19630 13532 19636 13566
rect 19590 13494 19636 13532
rect 19590 13460 19596 13494
rect 19630 13460 19636 13494
rect 19590 13422 19636 13460
rect 19890 13906 20338 13910
rect 20832 13906 20900 14056
rect 21086 14450 21300 15550
rect 23819 15513 24059 15584
rect 23449 15468 24059 15513
rect 23449 15434 23480 15468
rect 23514 15434 23580 15468
rect 23614 15434 23680 15468
rect 23714 15434 23780 15468
rect 23814 15434 23880 15468
rect 23914 15434 23980 15468
rect 24014 15434 24059 15468
rect 23449 15368 24059 15434
rect 23449 15334 23480 15368
rect 23514 15334 23580 15368
rect 23614 15334 23680 15368
rect 23714 15334 23780 15368
rect 23814 15334 23880 15368
rect 23914 15334 23980 15368
rect 24014 15334 24059 15368
rect 23449 15268 24059 15334
rect 24596 15330 25017 15338
rect 24596 15296 24609 15330
rect 24643 15296 24681 15330
rect 24715 15296 24753 15330
rect 24787 15296 24825 15330
rect 24859 15296 24897 15330
rect 24931 15296 24969 15330
rect 25003 15296 25017 15330
rect 24596 15288 25017 15296
rect 27127 15330 27548 15338
rect 27127 15296 27140 15330
rect 27174 15296 27212 15330
rect 27246 15296 27284 15330
rect 27318 15296 27356 15330
rect 27390 15296 27428 15330
rect 27462 15296 27500 15330
rect 27534 15296 27548 15330
rect 27127 15288 27548 15296
rect 23449 15234 23480 15268
rect 23514 15234 23580 15268
rect 23614 15234 23680 15268
rect 23714 15234 23780 15268
rect 23814 15234 23880 15268
rect 23914 15234 23980 15268
rect 24014 15234 24059 15268
rect 23449 15168 24059 15234
rect 23449 15134 23480 15168
rect 23514 15134 23580 15168
rect 23614 15134 23680 15168
rect 23714 15134 23780 15168
rect 23814 15134 23880 15168
rect 23914 15134 23980 15168
rect 24014 15134 24059 15168
rect 23449 15068 24059 15134
rect 23449 15034 23480 15068
rect 23514 15034 23580 15068
rect 23614 15034 23680 15068
rect 23714 15034 23780 15068
rect 23814 15034 23880 15068
rect 23914 15034 23980 15068
rect 24014 15034 24059 15068
rect 23449 14968 24059 15034
rect 23449 14934 23480 14968
rect 23514 14934 23580 14968
rect 23614 14934 23680 14968
rect 23714 14934 23780 14968
rect 23814 14934 23880 14968
rect 23914 14934 23980 14968
rect 24014 14934 24059 14968
rect 23449 14903 24059 14934
rect 28974 15242 29024 15256
rect 28974 15208 28982 15242
rect 29016 15208 29024 15242
rect 28974 15170 29024 15208
rect 28974 15136 28982 15170
rect 29016 15136 29024 15170
rect 28974 15098 29024 15136
rect 28974 15064 28982 15098
rect 29016 15064 29024 15098
rect 28974 15026 29024 15064
rect 28974 14992 28982 15026
rect 29016 14992 29024 15026
rect 28974 14954 29024 14992
rect 28974 14920 28982 14954
rect 29016 14920 29024 14954
rect 28974 14882 29024 14920
rect 28974 14848 28982 14882
rect 29016 14848 29024 14882
rect 28974 14835 29024 14848
rect 29188 15242 29438 15286
rect 29188 15215 29300 15242
rect 29334 15215 29438 15242
rect 29188 14843 29253 15215
rect 29369 14843 29438 15215
rect 29188 14748 29438 14843
rect 29610 15242 29660 15256
rect 29610 15208 29618 15242
rect 29652 15208 29660 15242
rect 29610 15170 29660 15208
rect 29610 15136 29618 15170
rect 29652 15136 29660 15170
rect 29610 15098 29660 15136
rect 29610 15064 29618 15098
rect 29652 15064 29660 15098
rect 29610 15026 29660 15064
rect 29610 14992 29618 15026
rect 29652 14992 29660 15026
rect 29610 14954 29660 14992
rect 29610 14920 29618 14954
rect 29652 14920 29660 14954
rect 29610 14882 29660 14920
rect 29610 14848 29618 14882
rect 29652 14848 29660 14882
rect 29610 14835 29660 14848
rect 21086 14416 21166 14450
rect 21200 14416 21300 14450
rect 21086 14378 21300 14416
rect 21086 14344 21166 14378
rect 21200 14344 21300 14378
rect 21086 14306 21300 14344
rect 21086 14272 21166 14306
rect 21200 14272 21300 14306
rect 21086 14234 21300 14272
rect 21086 14200 21166 14234
rect 21200 14200 21300 14234
rect 21086 14162 21300 14200
rect 21086 14128 21166 14162
rect 21200 14128 21300 14162
rect 21086 14090 21300 14128
rect 21086 14056 21166 14090
rect 21200 14056 21300 14090
rect 19890 13871 20904 13906
rect 19890 13499 19933 13871
rect 20305 13499 20904 13871
rect 19890 13428 20904 13499
rect 19590 13388 19596 13422
rect 19630 13388 19636 13422
rect 19590 13350 19636 13388
rect 19590 13316 19596 13350
rect 19630 13316 19636 13350
rect 19590 13278 19636 13316
rect 19590 13244 19596 13278
rect 19630 13244 19636 13278
rect 19590 13206 19636 13244
rect 19590 13172 19596 13206
rect 19630 13172 19636 13206
rect 19590 13134 19636 13172
rect 19590 13100 19596 13134
rect 19630 13100 19636 13134
rect 19590 13062 19636 13100
rect 19590 13028 19596 13062
rect 19630 13028 19636 13062
rect 19590 12990 19636 13028
rect 19590 12956 19596 12990
rect 19630 12956 19636 12990
rect 19590 12918 19636 12956
rect 19590 12884 19596 12918
rect 19630 12884 19636 12918
rect 19590 12846 19636 12884
rect 19590 12812 19596 12846
rect 19630 12812 19636 12846
rect 19590 12774 19636 12812
rect 19590 12740 19596 12774
rect 19630 12740 19636 12774
rect 19590 12702 19636 12740
rect 19590 12668 19596 12702
rect 19630 12668 19636 12702
rect 19590 12630 19636 12668
rect 19590 12596 19596 12630
rect 19630 12596 19636 12630
rect 19590 12558 19636 12596
rect 19590 12524 19596 12558
rect 19630 12524 19636 12558
rect 19590 12486 19636 12524
rect 19590 12452 19596 12486
rect 19630 12452 19636 12486
rect 19590 12414 19636 12452
rect 19590 12380 19596 12414
rect 19630 12380 19636 12414
rect 19590 12342 19636 12380
rect 19590 12308 19596 12342
rect 19630 12308 19636 12342
rect 19590 12270 19636 12308
rect 19590 12236 19596 12270
rect 19630 12236 19636 12270
rect 19590 12198 19636 12236
rect 19590 12164 19596 12198
rect 19630 12164 19636 12198
rect 18126 12108 18132 12142
rect 18166 12108 18172 12142
rect 18126 12070 18172 12108
rect 18126 12036 18132 12070
rect 18166 12036 18172 12070
rect 18126 11998 18172 12036
rect 18126 11964 18132 11998
rect 18166 11964 18172 11998
rect 16616 11882 16622 11916
rect 16656 11882 16662 11916
rect 16616 11844 16662 11882
rect 16616 11810 16622 11844
rect 16656 11810 16662 11844
rect 16616 11767 16662 11810
rect 17068 11926 17114 11930
rect 17068 11892 17074 11926
rect 17108 11892 17114 11926
rect 17068 11854 17114 11892
rect 17068 11820 17074 11854
rect 17108 11820 17114 11854
rect 17068 11777 17114 11820
rect 18126 11926 18172 11964
rect 18126 11892 18132 11926
rect 18166 11892 18172 11926
rect 18126 11854 18172 11892
rect 18466 12126 18646 12154
rect 18466 12119 18538 12126
rect 18572 12119 18646 12126
rect 18466 11939 18498 12119
rect 18614 11939 18646 12119
rect 18466 11910 18646 11939
rect 18466 11884 18538 11910
rect 18126 11820 18132 11854
rect 18166 11820 18172 11854
rect 18126 11777 18172 11820
rect 18532 11876 18538 11884
rect 18572 11884 18646 11910
rect 19590 12126 19636 12164
rect 19590 12092 19596 12126
rect 19630 12092 19636 12126
rect 19590 12054 19636 12092
rect 19590 12020 19596 12054
rect 19630 12020 19636 12054
rect 19590 11982 19636 12020
rect 19590 11948 19596 11982
rect 19630 11948 19636 11982
rect 19590 11910 19636 11948
rect 18572 11876 18578 11884
rect 18532 11838 18578 11876
rect 18532 11804 18538 11838
rect 18572 11804 18578 11838
rect 18532 11761 18578 11804
rect 19590 11876 19596 11910
rect 19630 11876 19636 11910
rect 19590 11838 19636 11876
rect 19590 11804 19596 11838
rect 19630 11804 19636 11838
rect 19590 11761 19636 11804
rect 17124 11730 18116 11736
rect 13044 11720 14036 11726
rect 13044 11686 13091 11720
rect 13125 11686 13163 11720
rect 13197 11686 13235 11720
rect 13269 11686 13307 11720
rect 13341 11686 13379 11720
rect 13413 11686 13451 11720
rect 13485 11686 13523 11720
rect 13557 11686 13595 11720
rect 13629 11686 13667 11720
rect 13701 11686 13739 11720
rect 13773 11686 13811 11720
rect 13845 11686 13883 11720
rect 13917 11686 13955 11720
rect 13989 11686 14036 11720
rect 13044 11680 14036 11686
rect 14102 11720 15094 11726
rect 14102 11686 14149 11720
rect 14183 11686 14221 11720
rect 14255 11686 14293 11720
rect 14327 11686 14365 11720
rect 14399 11686 14437 11720
rect 14471 11686 14509 11720
rect 14543 11686 14581 11720
rect 14615 11686 14653 11720
rect 14687 11686 14725 11720
rect 14759 11686 14797 11720
rect 14831 11686 14869 11720
rect 14903 11686 14941 11720
rect 14975 11686 15013 11720
rect 15047 11686 15094 11720
rect 14102 11680 15094 11686
rect 15614 11720 16606 11726
rect 15614 11686 15661 11720
rect 15695 11686 15733 11720
rect 15767 11686 15805 11720
rect 15839 11686 15877 11720
rect 15911 11686 15949 11720
rect 15983 11686 16021 11720
rect 16055 11686 16093 11720
rect 16127 11686 16165 11720
rect 16199 11686 16237 11720
rect 16271 11686 16309 11720
rect 16343 11686 16381 11720
rect 16415 11686 16453 11720
rect 16487 11686 16525 11720
rect 16559 11686 16606 11720
rect 17124 11696 17171 11730
rect 17205 11696 17243 11730
rect 17277 11696 17315 11730
rect 17349 11696 17387 11730
rect 17421 11696 17459 11730
rect 17493 11696 17531 11730
rect 17565 11696 17603 11730
rect 17637 11696 17675 11730
rect 17709 11696 17747 11730
rect 17781 11696 17819 11730
rect 17853 11696 17891 11730
rect 17925 11696 17963 11730
rect 17997 11696 18035 11730
rect 18069 11714 18342 11730
rect 18588 11714 19580 11720
rect 18069 11696 18635 11714
rect 17124 11690 18635 11696
rect 15614 11680 16606 11686
rect -8765 11242 -3667 11302
rect -8765 11236 -8573 11242
rect -8765 11202 -8722 11236
rect -8688 11202 -8650 11236
rect -8616 11202 -8573 11236
rect -8765 11196 -8573 11202
rect -8507 11236 -8315 11242
rect -8507 11202 -8464 11236
rect -8430 11202 -8392 11236
rect -8358 11202 -8315 11236
rect -8507 11196 -8315 11202
rect -8249 11236 -8057 11242
rect -8249 11202 -8206 11236
rect -8172 11202 -8134 11236
rect -8100 11202 -8057 11236
rect -8249 11196 -8057 11202
rect -7991 11236 -7799 11242
rect -7991 11202 -7948 11236
rect -7914 11202 -7876 11236
rect -7842 11202 -7799 11236
rect -7991 11196 -7799 11202
rect -7733 11236 -7541 11242
rect -7733 11202 -7690 11236
rect -7656 11202 -7618 11236
rect -7584 11202 -7541 11236
rect -7733 11196 -7541 11202
rect -7475 11236 -7283 11242
rect -7475 11202 -7432 11236
rect -7398 11202 -7360 11236
rect -7326 11202 -7283 11236
rect -7475 11196 -7283 11202
rect -7217 11236 -7025 11242
rect -7217 11202 -7174 11236
rect -7140 11202 -7102 11236
rect -7068 11202 -7025 11236
rect -7217 11196 -7025 11202
rect -6959 11236 -6767 11242
rect -6959 11202 -6916 11236
rect -6882 11202 -6844 11236
rect -6810 11202 -6767 11236
rect -6959 11196 -6767 11202
rect -6701 11236 -6509 11242
rect -6701 11202 -6658 11236
rect -6624 11202 -6586 11236
rect -6552 11202 -6509 11236
rect -6701 11196 -6509 11202
rect -6443 11236 -6251 11242
rect -6443 11202 -6400 11236
rect -6366 11202 -6328 11236
rect -6294 11202 -6251 11236
rect -6443 11196 -6251 11202
rect -6185 11236 -5993 11242
rect -6185 11202 -6142 11236
rect -6108 11202 -6070 11236
rect -6036 11202 -5993 11236
rect -6185 11196 -5993 11202
rect -5927 11236 -5735 11242
rect -5927 11202 -5884 11236
rect -5850 11202 -5812 11236
rect -5778 11202 -5735 11236
rect -5927 11196 -5735 11202
rect -5669 11236 -5477 11242
rect -5669 11202 -5626 11236
rect -5592 11202 -5554 11236
rect -5520 11202 -5477 11236
rect -5669 11196 -5477 11202
rect -5411 11236 -5219 11242
rect -5411 11202 -5368 11236
rect -5334 11202 -5296 11236
rect -5262 11202 -5219 11236
rect -5411 11196 -5219 11202
rect -5153 11236 -4961 11242
rect -5153 11202 -5110 11236
rect -5076 11202 -5038 11236
rect -5004 11202 -4961 11236
rect -5153 11196 -4961 11202
rect -4895 11236 -4703 11242
rect -4895 11202 -4852 11236
rect -4818 11202 -4780 11236
rect -4746 11202 -4703 11236
rect -4895 11196 -4703 11202
rect -4637 11236 -4445 11242
rect -4637 11202 -4594 11236
rect -4560 11202 -4522 11236
rect -4488 11202 -4445 11236
rect -4637 11196 -4445 11202
rect -4379 11236 -4187 11242
rect -4379 11202 -4336 11236
rect -4302 11202 -4264 11236
rect -4230 11202 -4187 11236
rect -4379 11196 -4187 11202
rect -4121 11236 -3929 11242
rect -4121 11202 -4078 11236
rect -4044 11202 -4006 11236
rect -3972 11202 -3929 11236
rect -4121 11196 -3929 11202
rect -3863 11236 -3671 11242
rect -3863 11202 -3820 11236
rect -3786 11202 -3748 11236
rect -3714 11202 -3671 11236
rect -3863 11196 -3671 11202
rect -8821 11149 -8775 11164
rect -8821 11115 -8815 11149
rect -8781 11115 -8775 11149
rect -8821 11077 -8775 11115
rect -8821 11043 -8815 11077
rect -8781 11043 -8775 11077
rect -8821 11005 -8775 11043
rect -8821 10971 -8815 11005
rect -8781 10971 -8775 11005
rect -8821 10933 -8775 10971
rect -8821 10899 -8815 10933
rect -8781 10899 -8775 10933
rect -8821 10861 -8775 10899
rect -8821 10827 -8815 10861
rect -8781 10827 -8775 10861
rect -8821 10789 -8775 10827
rect -8821 10755 -8815 10789
rect -8781 10755 -8775 10789
rect -8563 11149 -8517 11164
rect -8563 11115 -8557 11149
rect -8523 11115 -8517 11149
rect -8563 11077 -8517 11115
rect -8563 11043 -8557 11077
rect -8523 11043 -8517 11077
rect -8563 11005 -8517 11043
rect -8563 10971 -8557 11005
rect -8523 10971 -8517 11005
rect -8563 10933 -8517 10971
rect -8563 10899 -8557 10933
rect -8523 10899 -8517 10933
rect -8563 10861 -8517 10899
rect -8563 10827 -8557 10861
rect -8523 10827 -8517 10861
rect -8563 10789 -8517 10827
rect -8563 10773 -8557 10789
rect -8821 10717 -8775 10755
rect -8821 10683 -8815 10717
rect -8781 10683 -8775 10717
rect -8821 10645 -8775 10683
rect -8821 10611 -8815 10645
rect -8781 10611 -8775 10645
rect -8585 10766 -8557 10773
rect -8523 10773 -8517 10789
rect -8305 11149 -8259 11164
rect -8305 11115 -8299 11149
rect -8265 11115 -8259 11149
rect -8305 11077 -8259 11115
rect -8305 11043 -8299 11077
rect -8265 11043 -8259 11077
rect -8305 11005 -8259 11043
rect -8305 10971 -8299 11005
rect -8265 10971 -8259 11005
rect -8305 10933 -8259 10971
rect -8305 10899 -8299 10933
rect -8265 10899 -8259 10933
rect -8305 10861 -8259 10899
rect -8305 10827 -8299 10861
rect -8265 10827 -8259 10861
rect -8305 10789 -8259 10827
rect -8523 10766 -8496 10773
rect -8585 10714 -8566 10766
rect -8514 10714 -8496 10766
rect -8585 10702 -8557 10714
rect -8523 10702 -8496 10714
rect -8585 10650 -8566 10702
rect -8514 10650 -8496 10702
rect -8585 10645 -8496 10650
rect -8585 10640 -8557 10645
rect -8821 10573 -8775 10611
rect -10054 10492 -9276 10556
rect -8821 10539 -8815 10573
rect -8781 10539 -8775 10573
rect -8821 10501 -8775 10539
rect -8563 10611 -8557 10640
rect -8523 10640 -8496 10645
rect -8305 10755 -8299 10789
rect -8265 10755 -8259 10789
rect -8047 11149 -8001 11164
rect -8047 11115 -8041 11149
rect -8007 11115 -8001 11149
rect -8047 11077 -8001 11115
rect -8047 11043 -8041 11077
rect -8007 11043 -8001 11077
rect -8047 11005 -8001 11043
rect -8047 10971 -8041 11005
rect -8007 10971 -8001 11005
rect -8047 10933 -8001 10971
rect -8047 10899 -8041 10933
rect -8007 10899 -8001 10933
rect -8047 10861 -8001 10899
rect -8047 10827 -8041 10861
rect -8007 10827 -8001 10861
rect -8047 10789 -8001 10827
rect -8047 10773 -8041 10789
rect -8305 10717 -8259 10755
rect -8305 10683 -8299 10717
rect -8265 10683 -8259 10717
rect -8305 10645 -8259 10683
rect -8523 10611 -8517 10640
rect -8563 10573 -8517 10611
rect -8563 10539 -8557 10573
rect -8523 10539 -8517 10573
rect -8563 10501 -8517 10539
rect -8305 10611 -8299 10645
rect -8265 10611 -8259 10645
rect -8067 10755 -8041 10773
rect -8007 10773 -8001 10789
rect -7789 11149 -7743 11164
rect -7789 11115 -7783 11149
rect -7749 11115 -7743 11149
rect -7789 11077 -7743 11115
rect -7789 11043 -7783 11077
rect -7749 11043 -7743 11077
rect -7789 11005 -7743 11043
rect -7789 10971 -7783 11005
rect -7749 10971 -7743 11005
rect -7789 10933 -7743 10971
rect -7789 10899 -7783 10933
rect -7749 10899 -7743 10933
rect -7789 10861 -7743 10899
rect -7789 10827 -7783 10861
rect -7749 10827 -7743 10861
rect -7789 10789 -7743 10827
rect -8007 10755 -7981 10773
rect -8067 10733 -7981 10755
rect -8067 10681 -8051 10733
rect -7999 10681 -7981 10733
rect -8067 10645 -7981 10681
rect -8067 10640 -8041 10645
rect -8305 10573 -8259 10611
rect -8305 10539 -8299 10573
rect -8265 10539 -8259 10573
rect -8305 10501 -8259 10539
rect -8047 10611 -8041 10640
rect -8007 10640 -7981 10645
rect -7789 10755 -7783 10789
rect -7749 10755 -7743 10789
rect -7531 11149 -7485 11164
rect -7531 11115 -7525 11149
rect -7491 11115 -7485 11149
rect -7531 11077 -7485 11115
rect -7531 11043 -7525 11077
rect -7491 11043 -7485 11077
rect -7531 11005 -7485 11043
rect -7531 10971 -7525 11005
rect -7491 10971 -7485 11005
rect -7531 10933 -7485 10971
rect -7531 10899 -7525 10933
rect -7491 10899 -7485 10933
rect -7531 10861 -7485 10899
rect -7531 10827 -7525 10861
rect -7491 10827 -7485 10861
rect -7531 10789 -7485 10827
rect -7531 10773 -7525 10789
rect -7789 10717 -7743 10755
rect -7789 10683 -7783 10717
rect -7749 10683 -7743 10717
rect -7789 10645 -7743 10683
rect -8007 10611 -8001 10640
rect -8047 10573 -8001 10611
rect -8047 10539 -8041 10573
rect -8007 10539 -8001 10573
rect -8047 10501 -8001 10539
rect -7789 10611 -7783 10645
rect -7749 10611 -7743 10645
rect -7549 10755 -7525 10773
rect -7491 10773 -7485 10789
rect -7273 11149 -7227 11164
rect -7273 11115 -7267 11149
rect -7233 11115 -7227 11149
rect -7273 11077 -7227 11115
rect -7273 11043 -7267 11077
rect -7233 11043 -7227 11077
rect -7273 11005 -7227 11043
rect -7273 10971 -7267 11005
rect -7233 10971 -7227 11005
rect -7273 10933 -7227 10971
rect -7273 10899 -7267 10933
rect -7233 10899 -7227 10933
rect -7273 10861 -7227 10899
rect -7273 10827 -7267 10861
rect -7233 10827 -7227 10861
rect -7273 10789 -7227 10827
rect -7491 10755 -7466 10773
rect -7549 10732 -7466 10755
rect -7549 10680 -7534 10732
rect -7482 10680 -7466 10732
rect -7549 10645 -7466 10680
rect -7549 10640 -7525 10645
rect -7789 10573 -7743 10611
rect -7789 10539 -7783 10573
rect -7749 10539 -7743 10573
rect -7789 10501 -7743 10539
rect -7531 10611 -7525 10640
rect -7491 10640 -7466 10645
rect -7273 10755 -7267 10789
rect -7233 10755 -7227 10789
rect -7015 11149 -6969 11164
rect -7015 11115 -7009 11149
rect -6975 11115 -6969 11149
rect -7015 11077 -6969 11115
rect -7015 11043 -7009 11077
rect -6975 11043 -6969 11077
rect -7015 11005 -6969 11043
rect -7015 10971 -7009 11005
rect -6975 10971 -6969 11005
rect -7015 10933 -6969 10971
rect -7015 10899 -7009 10933
rect -6975 10899 -6969 10933
rect -7015 10861 -6969 10899
rect -7015 10827 -7009 10861
rect -6975 10827 -6969 10861
rect -7015 10789 -6969 10827
rect -7015 10773 -7009 10789
rect -7273 10717 -7227 10755
rect -7273 10683 -7267 10717
rect -7233 10683 -7227 10717
rect -7273 10645 -7227 10683
rect -7491 10611 -7485 10640
rect -7531 10573 -7485 10611
rect -7531 10539 -7525 10573
rect -7491 10539 -7485 10573
rect -7531 10501 -7485 10539
rect -7273 10611 -7267 10645
rect -7233 10611 -7227 10645
rect -7034 10755 -7009 10773
rect -6975 10773 -6969 10789
rect -6757 11149 -6711 11164
rect -6757 11115 -6751 11149
rect -6717 11115 -6711 11149
rect -6757 11077 -6711 11115
rect -6757 11043 -6751 11077
rect -6717 11043 -6711 11077
rect -6757 11005 -6711 11043
rect -6757 10971 -6751 11005
rect -6717 10971 -6711 11005
rect -6757 10933 -6711 10971
rect -6757 10899 -6751 10933
rect -6717 10899 -6711 10933
rect -6757 10861 -6711 10899
rect -6757 10827 -6751 10861
rect -6717 10827 -6711 10861
rect -6757 10789 -6711 10827
rect -6975 10755 -6949 10773
rect -7034 10733 -6949 10755
rect -7034 10681 -7018 10733
rect -6966 10681 -6949 10733
rect -7034 10645 -6949 10681
rect -7034 10640 -7009 10645
rect -7273 10573 -7227 10611
rect -7273 10539 -7267 10573
rect -7233 10539 -7227 10573
rect -7273 10501 -7227 10539
rect -7015 10611 -7009 10640
rect -6975 10640 -6949 10645
rect -6757 10755 -6751 10789
rect -6717 10755 -6711 10789
rect -6499 11149 -6453 11164
rect -6499 11115 -6493 11149
rect -6459 11115 -6453 11149
rect -6499 11077 -6453 11115
rect -6499 11043 -6493 11077
rect -6459 11043 -6453 11077
rect -6499 11005 -6453 11043
rect -6499 10971 -6493 11005
rect -6459 10971 -6453 11005
rect -6499 10933 -6453 10971
rect -6499 10899 -6493 10933
rect -6459 10899 -6453 10933
rect -6499 10861 -6453 10899
rect -6499 10827 -6493 10861
rect -6459 10827 -6453 10861
rect -6499 10789 -6453 10827
rect -6499 10773 -6493 10789
rect -6757 10717 -6711 10755
rect -6757 10683 -6751 10717
rect -6717 10683 -6711 10717
rect -6757 10645 -6711 10683
rect -6975 10611 -6969 10640
rect -7015 10573 -6969 10611
rect -7015 10539 -7009 10573
rect -6975 10539 -6969 10573
rect -7015 10501 -6969 10539
rect -6757 10611 -6751 10645
rect -6717 10611 -6711 10645
rect -6518 10755 -6493 10773
rect -6459 10773 -6453 10789
rect -6241 11149 -6195 11164
rect -6241 11115 -6235 11149
rect -6201 11115 -6195 11149
rect -6241 11077 -6195 11115
rect -6241 11043 -6235 11077
rect -6201 11043 -6195 11077
rect -6241 11005 -6195 11043
rect -6241 10971 -6235 11005
rect -6201 10971 -6195 11005
rect -6241 10933 -6195 10971
rect -6241 10899 -6235 10933
rect -6201 10899 -6195 10933
rect -6241 10861 -6195 10899
rect -6241 10827 -6235 10861
rect -6201 10827 -6195 10861
rect -6241 10789 -6195 10827
rect -6459 10755 -6432 10773
rect -6518 10731 -6432 10755
rect -6518 10679 -6502 10731
rect -6450 10679 -6432 10731
rect -6518 10645 -6432 10679
rect -6518 10640 -6493 10645
rect -6757 10573 -6711 10611
rect -6757 10539 -6751 10573
rect -6717 10539 -6711 10573
rect -6757 10501 -6711 10539
rect -6499 10611 -6493 10640
rect -6459 10640 -6432 10645
rect -6241 10755 -6235 10789
rect -6201 10755 -6195 10789
rect -5983 11149 -5937 11164
rect -5983 11115 -5977 11149
rect -5943 11115 -5937 11149
rect -5983 11077 -5937 11115
rect -5983 11043 -5977 11077
rect -5943 11043 -5937 11077
rect -5983 11005 -5937 11043
rect -5983 10971 -5977 11005
rect -5943 10971 -5937 11005
rect -5983 10933 -5937 10971
rect -5983 10899 -5977 10933
rect -5943 10899 -5937 10933
rect -5983 10861 -5937 10899
rect -5983 10827 -5977 10861
rect -5943 10827 -5937 10861
rect -5983 10789 -5937 10827
rect -5983 10773 -5977 10789
rect -6241 10717 -6195 10755
rect -6241 10683 -6235 10717
rect -6201 10683 -6195 10717
rect -6241 10645 -6195 10683
rect -6459 10611 -6453 10640
rect -6499 10573 -6453 10611
rect -6499 10539 -6493 10573
rect -6459 10539 -6453 10573
rect -6499 10501 -6453 10539
rect -6241 10611 -6235 10645
rect -6201 10611 -6195 10645
rect -6000 10755 -5977 10773
rect -5943 10773 -5937 10789
rect -5725 11149 -5679 11164
rect -5725 11115 -5719 11149
rect -5685 11115 -5679 11149
rect -5725 11077 -5679 11115
rect -5725 11043 -5719 11077
rect -5685 11043 -5679 11077
rect -5725 11005 -5679 11043
rect -5725 10971 -5719 11005
rect -5685 10971 -5679 11005
rect -5725 10933 -5679 10971
rect -5725 10899 -5719 10933
rect -5685 10899 -5679 10933
rect -5725 10861 -5679 10899
rect -5725 10827 -5719 10861
rect -5685 10827 -5679 10861
rect -5725 10789 -5679 10827
rect -5943 10755 -5920 10773
rect -6000 10732 -5920 10755
rect -6000 10680 -5986 10732
rect -5934 10680 -5920 10732
rect -6000 10645 -5920 10680
rect -6000 10640 -5977 10645
rect -6241 10573 -6195 10611
rect -6241 10539 -6235 10573
rect -6201 10539 -6195 10573
rect -6241 10501 -6195 10539
rect -5983 10611 -5977 10640
rect -5943 10640 -5920 10645
rect -5725 10755 -5719 10789
rect -5685 10755 -5679 10789
rect -5467 11149 -5421 11164
rect -5467 11115 -5461 11149
rect -5427 11115 -5421 11149
rect -5467 11077 -5421 11115
rect -5467 11043 -5461 11077
rect -5427 11043 -5421 11077
rect -5467 11005 -5421 11043
rect -5467 10971 -5461 11005
rect -5427 10971 -5421 11005
rect -5467 10933 -5421 10971
rect -5467 10899 -5461 10933
rect -5427 10899 -5421 10933
rect -5467 10861 -5421 10899
rect -5467 10827 -5461 10861
rect -5427 10827 -5421 10861
rect -5467 10789 -5421 10827
rect -5467 10773 -5461 10789
rect -5725 10717 -5679 10755
rect -5725 10683 -5719 10717
rect -5685 10683 -5679 10717
rect -5725 10645 -5679 10683
rect -5943 10611 -5937 10640
rect -5983 10573 -5937 10611
rect -5983 10539 -5977 10573
rect -5943 10539 -5937 10573
rect -5983 10501 -5937 10539
rect -5725 10611 -5719 10645
rect -5685 10611 -5679 10645
rect -5484 10755 -5461 10773
rect -5427 10773 -5421 10789
rect -5209 11149 -5163 11164
rect -5209 11115 -5203 11149
rect -5169 11115 -5163 11149
rect -5209 11077 -5163 11115
rect -5209 11043 -5203 11077
rect -5169 11043 -5163 11077
rect -5209 11005 -5163 11043
rect -5209 10971 -5203 11005
rect -5169 10971 -5163 11005
rect -5209 10933 -5163 10971
rect -5209 10899 -5203 10933
rect -5169 10899 -5163 10933
rect -5209 10861 -5163 10899
rect -5209 10827 -5203 10861
rect -5169 10827 -5163 10861
rect -5209 10789 -5163 10827
rect -5427 10755 -5404 10773
rect -5484 10731 -5404 10755
rect -5484 10679 -5470 10731
rect -5418 10679 -5404 10731
rect -5484 10645 -5404 10679
rect -5484 10640 -5461 10645
rect -5725 10573 -5679 10611
rect -5725 10539 -5719 10573
rect -5685 10539 -5679 10573
rect -5725 10501 -5679 10539
rect -5467 10611 -5461 10640
rect -5427 10640 -5404 10645
rect -5209 10755 -5203 10789
rect -5169 10755 -5163 10789
rect -4951 11149 -4905 11164
rect -4951 11115 -4945 11149
rect -4911 11115 -4905 11149
rect -4951 11077 -4905 11115
rect -4951 11043 -4945 11077
rect -4911 11043 -4905 11077
rect -4951 11005 -4905 11043
rect -4951 10971 -4945 11005
rect -4911 10971 -4905 11005
rect -4951 10933 -4905 10971
rect -4951 10899 -4945 10933
rect -4911 10899 -4905 10933
rect -4951 10861 -4905 10899
rect -4951 10827 -4945 10861
rect -4911 10827 -4905 10861
rect -4951 10789 -4905 10827
rect -4951 10773 -4945 10789
rect -5209 10717 -5163 10755
rect -5209 10683 -5203 10717
rect -5169 10683 -5163 10717
rect -5209 10645 -5163 10683
rect -5427 10611 -5421 10640
rect -5467 10573 -5421 10611
rect -5467 10539 -5461 10573
rect -5427 10539 -5421 10573
rect -5467 10501 -5421 10539
rect -5209 10611 -5203 10645
rect -5169 10611 -5163 10645
rect -4969 10755 -4945 10773
rect -4911 10773 -4905 10789
rect -4693 11149 -4647 11164
rect -4693 11115 -4687 11149
rect -4653 11115 -4647 11149
rect -4693 11077 -4647 11115
rect -4693 11043 -4687 11077
rect -4653 11043 -4647 11077
rect -4693 11005 -4647 11043
rect -4693 10971 -4687 11005
rect -4653 10971 -4647 11005
rect -4693 10933 -4647 10971
rect -4693 10899 -4687 10933
rect -4653 10899 -4647 10933
rect -4693 10861 -4647 10899
rect -4693 10827 -4687 10861
rect -4653 10827 -4647 10861
rect -4693 10789 -4647 10827
rect -4911 10755 -4887 10773
rect -4969 10732 -4887 10755
rect -4969 10680 -4954 10732
rect -4902 10680 -4887 10732
rect -4969 10645 -4887 10680
rect -4969 10640 -4945 10645
rect -5209 10573 -5163 10611
rect -5209 10539 -5203 10573
rect -5169 10539 -5163 10573
rect -5209 10501 -5163 10539
rect -4951 10611 -4945 10640
rect -4911 10640 -4887 10645
rect -4693 10755 -4687 10789
rect -4653 10755 -4647 10789
rect -4435 11149 -4389 11164
rect -4435 11115 -4429 11149
rect -4395 11115 -4389 11149
rect -4435 11077 -4389 11115
rect -4435 11043 -4429 11077
rect -4395 11043 -4389 11077
rect -4435 11005 -4389 11043
rect -4435 10971 -4429 11005
rect -4395 10971 -4389 11005
rect -4435 10933 -4389 10971
rect -4435 10899 -4429 10933
rect -4395 10899 -4389 10933
rect -4435 10861 -4389 10899
rect -4435 10827 -4429 10861
rect -4395 10827 -4389 10861
rect -4435 10789 -4389 10827
rect -4435 10773 -4429 10789
rect -4693 10717 -4647 10755
rect -4693 10683 -4687 10717
rect -4653 10683 -4647 10717
rect -4693 10645 -4647 10683
rect -4911 10611 -4905 10640
rect -4951 10573 -4905 10611
rect -4951 10539 -4945 10573
rect -4911 10539 -4905 10573
rect -4951 10501 -4905 10539
rect -4693 10611 -4687 10645
rect -4653 10611 -4647 10645
rect -4451 10755 -4429 10773
rect -4395 10773 -4389 10789
rect -4177 11149 -4131 11164
rect -4177 11115 -4171 11149
rect -4137 11115 -4131 11149
rect -4177 11077 -4131 11115
rect -4177 11043 -4171 11077
rect -4137 11043 -4131 11077
rect -4177 11005 -4131 11043
rect -4177 10971 -4171 11005
rect -4137 10971 -4131 11005
rect -4177 10933 -4131 10971
rect -4177 10899 -4171 10933
rect -4137 10899 -4131 10933
rect -4177 10861 -4131 10899
rect -4177 10827 -4171 10861
rect -4137 10827 -4131 10861
rect -4177 10789 -4131 10827
rect -4395 10755 -4372 10773
rect -4451 10732 -4372 10755
rect -4451 10680 -4438 10732
rect -4386 10680 -4372 10732
rect -4451 10645 -4372 10680
rect -4451 10640 -4429 10645
rect -4693 10573 -4647 10611
rect -4693 10539 -4687 10573
rect -4653 10539 -4647 10573
rect -4693 10501 -4647 10539
rect -4435 10611 -4429 10640
rect -4395 10640 -4372 10645
rect -4177 10755 -4171 10789
rect -4137 10755 -4131 10789
rect -3919 11149 -3873 11164
rect -3919 11115 -3913 11149
rect -3879 11115 -3873 11149
rect -3919 11077 -3873 11115
rect -3919 11043 -3913 11077
rect -3879 11043 -3873 11077
rect -3919 11005 -3873 11043
rect -3919 10971 -3913 11005
rect -3879 10971 -3873 11005
rect -3919 10933 -3873 10971
rect -3919 10899 -3913 10933
rect -3879 10899 -3873 10933
rect -3919 10861 -3873 10899
rect -3919 10827 -3913 10861
rect -3879 10827 -3873 10861
rect -3919 10789 -3873 10827
rect -3919 10773 -3913 10789
rect -4177 10717 -4131 10755
rect -4177 10683 -4171 10717
rect -4137 10683 -4131 10717
rect -4177 10645 -4131 10683
rect -4395 10611 -4389 10640
rect -4435 10573 -4389 10611
rect -4435 10539 -4429 10573
rect -4395 10539 -4389 10573
rect -4435 10501 -4389 10539
rect -4177 10611 -4171 10645
rect -4137 10611 -4131 10645
rect -3936 10755 -3913 10773
rect -3879 10773 -3873 10789
rect -3661 11149 -3615 11164
rect -3661 11115 -3655 11149
rect -3621 11115 -3615 11149
rect -3661 11077 -3615 11115
rect -3661 11043 -3655 11077
rect -3621 11043 -3615 11077
rect -3661 11005 -3615 11043
rect -3661 10971 -3655 11005
rect -3621 10971 -3615 11005
rect -3661 10933 -3615 10971
rect -3661 10899 -3655 10933
rect -3621 10899 -3615 10933
rect -3661 10861 -3615 10899
rect -3661 10827 -3655 10861
rect -3621 10827 -3615 10861
rect -3661 10789 -3615 10827
rect -3879 10755 -3855 10773
rect -3936 10732 -3855 10755
rect -3936 10680 -3922 10732
rect -3870 10680 -3855 10732
rect -3936 10645 -3855 10680
rect -3936 10640 -3913 10645
rect -4177 10573 -4131 10611
rect -4177 10539 -4171 10573
rect -4137 10539 -4131 10573
rect -4177 10501 -4131 10539
rect -3919 10611 -3913 10640
rect -3879 10640 -3855 10645
rect -3661 10755 -3655 10789
rect -3621 10755 -3615 10789
rect -3661 10717 -3615 10755
rect -3661 10683 -3655 10717
rect -3621 10683 -3615 10717
rect -3661 10645 -3615 10683
rect -3879 10611 -3873 10640
rect -3919 10573 -3873 10611
rect -3919 10539 -3913 10573
rect -3879 10539 -3873 10573
rect -3919 10501 -3873 10539
rect -3661 10611 -3655 10645
rect -3621 10611 -3615 10645
rect -3661 10573 -3615 10611
rect -3661 10539 -3655 10573
rect -3621 10539 -3615 10573
rect -3661 10501 -3615 10539
rect 13086 10950 13746 11030
rect 13086 10916 13152 10950
rect 13186 10916 13252 10950
rect 13286 10916 13352 10950
rect 13386 10916 13452 10950
rect 13486 10916 13552 10950
rect 13586 10916 13652 10950
rect 13686 10916 13746 10950
rect 13086 10863 13746 10916
rect 13086 10850 13276 10863
rect 13584 10850 13746 10863
rect 13086 10816 13152 10850
rect 13186 10816 13252 10850
rect 13586 10816 13652 10850
rect 13686 10816 13746 10850
rect 13086 10750 13276 10816
rect 13584 10750 13746 10816
rect 13086 10716 13152 10750
rect 13186 10716 13252 10750
rect 13586 10716 13652 10750
rect 13686 10716 13746 10750
rect 13086 10650 13276 10716
rect 13584 10650 13746 10716
rect 13086 10616 13152 10650
rect 13186 10616 13252 10650
rect 13586 10616 13652 10650
rect 13686 10616 13746 10650
rect 13086 10555 13276 10616
rect 13584 10555 13746 10616
rect 13086 10550 13746 10555
rect 13086 10516 13152 10550
rect 13186 10516 13252 10550
rect 13286 10516 13352 10550
rect 13386 10516 13452 10550
rect 13486 10516 13552 10550
rect 13586 10516 13652 10550
rect 13686 10516 13746 10550
rect -10054 9928 -9976 10492
rect -9412 10086 -9276 10492
rect -8856 10486 -8815 10501
rect -8781 10486 -8754 10501
rect -8856 10434 -8824 10486
rect -8772 10434 -8754 10486
rect -8856 10429 -8754 10434
rect -8856 10422 -8815 10429
rect -8781 10422 -8754 10429
rect -8856 10370 -8824 10422
rect -8772 10370 -8754 10422
rect -8856 10359 -8754 10370
rect -8563 10467 -8557 10501
rect -8523 10467 -8517 10501
rect -8563 10429 -8517 10467
rect -8563 10395 -8557 10429
rect -8523 10395 -8517 10429
rect -8821 10357 -8775 10359
rect -8821 10323 -8815 10357
rect -8781 10323 -8775 10357
rect -8821 10285 -8775 10323
rect -8821 10251 -8815 10285
rect -8781 10251 -8775 10285
rect -8821 10213 -8775 10251
rect -8821 10179 -8815 10213
rect -8781 10179 -8775 10213
rect -8821 10164 -8775 10179
rect -8563 10357 -8517 10395
rect -8324 10488 -8299 10501
rect -8265 10488 -8239 10501
rect -8324 10436 -8308 10488
rect -8256 10436 -8239 10488
rect -8324 10429 -8239 10436
rect -8324 10424 -8299 10429
rect -8265 10424 -8239 10429
rect -8324 10372 -8308 10424
rect -8256 10372 -8239 10424
rect -8324 10359 -8239 10372
rect -8047 10467 -8041 10501
rect -8007 10467 -8001 10501
rect -8047 10429 -8001 10467
rect -8047 10395 -8041 10429
rect -8007 10395 -8001 10429
rect -8563 10323 -8557 10357
rect -8523 10323 -8517 10357
rect -8563 10285 -8517 10323
rect -8563 10251 -8557 10285
rect -8523 10251 -8517 10285
rect -8563 10213 -8517 10251
rect -8563 10179 -8557 10213
rect -8523 10179 -8517 10213
rect -8563 10164 -8517 10179
rect -8305 10357 -8259 10359
rect -8305 10323 -8299 10357
rect -8265 10323 -8259 10357
rect -8305 10285 -8259 10323
rect -8305 10251 -8299 10285
rect -8265 10251 -8259 10285
rect -8305 10213 -8259 10251
rect -8305 10179 -8299 10213
rect -8265 10179 -8259 10213
rect -8305 10164 -8259 10179
rect -8047 10357 -8001 10395
rect -7808 10488 -7783 10501
rect -7749 10488 -7723 10501
rect -7808 10436 -7792 10488
rect -7740 10436 -7723 10488
rect -7808 10429 -7723 10436
rect -7808 10424 -7783 10429
rect -7749 10424 -7723 10429
rect -7808 10372 -7792 10424
rect -7740 10372 -7723 10424
rect -7808 10359 -7723 10372
rect -7531 10467 -7525 10501
rect -7491 10467 -7485 10501
rect -7531 10429 -7485 10467
rect -7531 10395 -7525 10429
rect -7491 10395 -7485 10429
rect -8047 10323 -8041 10357
rect -8007 10323 -8001 10357
rect -8047 10285 -8001 10323
rect -8047 10251 -8041 10285
rect -8007 10251 -8001 10285
rect -8047 10213 -8001 10251
rect -8047 10179 -8041 10213
rect -8007 10179 -8001 10213
rect -8047 10164 -8001 10179
rect -7789 10357 -7743 10359
rect -7789 10323 -7783 10357
rect -7749 10323 -7743 10357
rect -7789 10285 -7743 10323
rect -7789 10251 -7783 10285
rect -7749 10251 -7743 10285
rect -7789 10213 -7743 10251
rect -7789 10179 -7783 10213
rect -7749 10179 -7743 10213
rect -7789 10164 -7743 10179
rect -7531 10357 -7485 10395
rect -7290 10487 -7267 10501
rect -7233 10487 -7209 10501
rect -7290 10435 -7276 10487
rect -7224 10435 -7209 10487
rect -7290 10429 -7209 10435
rect -7290 10423 -7267 10429
rect -7233 10423 -7209 10429
rect -7290 10371 -7276 10423
rect -7224 10371 -7209 10423
rect -7290 10359 -7209 10371
rect -7015 10467 -7009 10501
rect -6975 10467 -6969 10501
rect -7015 10429 -6969 10467
rect -7015 10395 -7009 10429
rect -6975 10395 -6969 10429
rect -7531 10323 -7525 10357
rect -7491 10323 -7485 10357
rect -7531 10285 -7485 10323
rect -7531 10251 -7525 10285
rect -7491 10251 -7485 10285
rect -7531 10213 -7485 10251
rect -7531 10179 -7525 10213
rect -7491 10179 -7485 10213
rect -7531 10164 -7485 10179
rect -7273 10357 -7227 10359
rect -7273 10323 -7267 10357
rect -7233 10323 -7227 10357
rect -7273 10285 -7227 10323
rect -7273 10251 -7267 10285
rect -7233 10251 -7227 10285
rect -7273 10213 -7227 10251
rect -7273 10179 -7267 10213
rect -7233 10179 -7227 10213
rect -7273 10164 -7227 10179
rect -7015 10357 -6969 10395
rect -6776 10488 -6751 10501
rect -6717 10488 -6692 10501
rect -6776 10436 -6760 10488
rect -6708 10436 -6692 10488
rect -6776 10429 -6692 10436
rect -6776 10424 -6751 10429
rect -6717 10424 -6692 10429
rect -6776 10372 -6760 10424
rect -6708 10372 -6692 10424
rect -6776 10359 -6692 10372
rect -6499 10467 -6493 10501
rect -6459 10467 -6453 10501
rect -6499 10429 -6453 10467
rect -6499 10395 -6493 10429
rect -6459 10395 -6453 10429
rect -7015 10323 -7009 10357
rect -6975 10323 -6969 10357
rect -7015 10285 -6969 10323
rect -7015 10251 -7009 10285
rect -6975 10251 -6969 10285
rect -7015 10213 -6969 10251
rect -7015 10179 -7009 10213
rect -6975 10179 -6969 10213
rect -7015 10164 -6969 10179
rect -6757 10357 -6711 10359
rect -6757 10323 -6751 10357
rect -6717 10323 -6711 10357
rect -6757 10285 -6711 10323
rect -6757 10251 -6751 10285
rect -6717 10251 -6711 10285
rect -6757 10213 -6711 10251
rect -6757 10179 -6751 10213
rect -6717 10179 -6711 10213
rect -6757 10164 -6711 10179
rect -6499 10357 -6453 10395
rect -6260 10489 -6235 10501
rect -6201 10489 -6176 10501
rect -6260 10437 -6243 10489
rect -6191 10437 -6176 10489
rect -6260 10429 -6176 10437
rect -6260 10425 -6235 10429
rect -6201 10425 -6176 10429
rect -6260 10373 -6243 10425
rect -6191 10373 -6176 10425
rect -6260 10359 -6176 10373
rect -5983 10467 -5977 10501
rect -5943 10467 -5937 10501
rect -5983 10429 -5937 10467
rect -5983 10395 -5977 10429
rect -5943 10395 -5937 10429
rect -6499 10323 -6493 10357
rect -6459 10323 -6453 10357
rect -6499 10285 -6453 10323
rect -6499 10251 -6493 10285
rect -6459 10251 -6453 10285
rect -6499 10213 -6453 10251
rect -6499 10179 -6493 10213
rect -6459 10179 -6453 10213
rect -6499 10164 -6453 10179
rect -6241 10357 -6195 10359
rect -6241 10323 -6235 10357
rect -6201 10323 -6195 10357
rect -6241 10285 -6195 10323
rect -6241 10251 -6235 10285
rect -6201 10251 -6195 10285
rect -6241 10213 -6195 10251
rect -6241 10179 -6235 10213
rect -6201 10179 -6195 10213
rect -6241 10164 -6195 10179
rect -5983 10357 -5937 10395
rect -5742 10486 -5719 10501
rect -5685 10486 -5657 10501
rect -5742 10434 -5728 10486
rect -5676 10434 -5657 10486
rect -5742 10429 -5657 10434
rect -5742 10422 -5719 10429
rect -5685 10422 -5657 10429
rect -5742 10370 -5728 10422
rect -5676 10370 -5657 10422
rect -5742 10359 -5657 10370
rect -5467 10467 -5461 10501
rect -5427 10467 -5421 10501
rect -5467 10429 -5421 10467
rect -5467 10395 -5461 10429
rect -5427 10395 -5421 10429
rect -5983 10323 -5977 10357
rect -5943 10323 -5937 10357
rect -5983 10285 -5937 10323
rect -5983 10251 -5977 10285
rect -5943 10251 -5937 10285
rect -5983 10213 -5937 10251
rect -5983 10179 -5977 10213
rect -5943 10179 -5937 10213
rect -5983 10164 -5937 10179
rect -5725 10357 -5679 10359
rect -5725 10323 -5719 10357
rect -5685 10323 -5679 10357
rect -5725 10285 -5679 10323
rect -5725 10251 -5719 10285
rect -5685 10251 -5679 10285
rect -5725 10213 -5679 10251
rect -5725 10179 -5719 10213
rect -5685 10179 -5679 10213
rect -5725 10164 -5679 10179
rect -5467 10357 -5421 10395
rect -5227 10487 -5203 10501
rect -5169 10487 -5145 10501
rect -5227 10435 -5213 10487
rect -5161 10435 -5145 10487
rect -5227 10429 -5145 10435
rect -5227 10423 -5203 10429
rect -5169 10423 -5145 10429
rect -5227 10371 -5213 10423
rect -5161 10371 -5145 10423
rect -5227 10359 -5145 10371
rect -4951 10467 -4945 10501
rect -4911 10467 -4905 10501
rect -4951 10429 -4905 10467
rect -4951 10395 -4945 10429
rect -4911 10395 -4905 10429
rect -5467 10323 -5461 10357
rect -5427 10323 -5421 10357
rect -5467 10285 -5421 10323
rect -5467 10251 -5461 10285
rect -5427 10251 -5421 10285
rect -5467 10213 -5421 10251
rect -5467 10179 -5461 10213
rect -5427 10179 -5421 10213
rect -5467 10164 -5421 10179
rect -5209 10357 -5163 10359
rect -5209 10323 -5203 10357
rect -5169 10323 -5163 10357
rect -5209 10285 -5163 10323
rect -5209 10251 -5203 10285
rect -5169 10251 -5163 10285
rect -5209 10213 -5163 10251
rect -5209 10179 -5203 10213
rect -5169 10179 -5163 10213
rect -5209 10164 -5163 10179
rect -4951 10357 -4905 10395
rect -4710 10488 -4687 10501
rect -4653 10488 -4629 10501
rect -4710 10436 -4696 10488
rect -4644 10436 -4629 10488
rect -4710 10429 -4629 10436
rect -4710 10424 -4687 10429
rect -4653 10424 -4629 10429
rect -4710 10372 -4696 10424
rect -4644 10372 -4629 10424
rect -4710 10359 -4629 10372
rect -4435 10467 -4429 10501
rect -4395 10467 -4389 10501
rect -4435 10429 -4389 10467
rect -4435 10395 -4429 10429
rect -4395 10395 -4389 10429
rect -4951 10323 -4945 10357
rect -4911 10323 -4905 10357
rect -4951 10285 -4905 10323
rect -4951 10251 -4945 10285
rect -4911 10251 -4905 10285
rect -4951 10213 -4905 10251
rect -4951 10179 -4945 10213
rect -4911 10179 -4905 10213
rect -4951 10164 -4905 10179
rect -4693 10357 -4647 10359
rect -4693 10323 -4687 10357
rect -4653 10323 -4647 10357
rect -4693 10285 -4647 10323
rect -4693 10251 -4687 10285
rect -4653 10251 -4647 10285
rect -4693 10213 -4647 10251
rect -4693 10179 -4687 10213
rect -4653 10179 -4647 10213
rect -4693 10164 -4647 10179
rect -4435 10357 -4389 10395
rect -4196 10487 -4171 10501
rect -4137 10487 -4112 10501
rect -4196 10435 -4180 10487
rect -4128 10435 -4112 10487
rect -4196 10429 -4112 10435
rect -4196 10423 -4171 10429
rect -4137 10423 -4112 10429
rect -4196 10371 -4180 10423
rect -4128 10371 -4112 10423
rect -4196 10359 -4112 10371
rect -3919 10467 -3913 10501
rect -3879 10467 -3873 10501
rect -3919 10429 -3873 10467
rect -3919 10395 -3913 10429
rect -3879 10395 -3873 10429
rect -4435 10323 -4429 10357
rect -4395 10323 -4389 10357
rect -4435 10285 -4389 10323
rect -4435 10251 -4429 10285
rect -4395 10251 -4389 10285
rect -4435 10213 -4389 10251
rect -4435 10179 -4429 10213
rect -4395 10179 -4389 10213
rect -4435 10164 -4389 10179
rect -4177 10357 -4131 10359
rect -4177 10323 -4171 10357
rect -4137 10323 -4131 10357
rect -4177 10285 -4131 10323
rect -4177 10251 -4171 10285
rect -4137 10251 -4131 10285
rect -4177 10213 -4131 10251
rect -4177 10179 -4171 10213
rect -4137 10179 -4131 10213
rect -4177 10164 -4131 10179
rect -3919 10357 -3873 10395
rect -3679 10487 -3655 10501
rect -3621 10487 -3596 10501
rect -3679 10435 -3664 10487
rect -3612 10435 -3596 10487
rect -3679 10429 -3596 10435
rect -3679 10423 -3655 10429
rect -3621 10423 -3596 10429
rect -3679 10371 -3664 10423
rect -3612 10371 -3596 10423
rect -3679 10359 -3596 10371
rect 13086 10450 13746 10516
rect 13086 10416 13152 10450
rect 13186 10416 13252 10450
rect 13286 10416 13352 10450
rect 13386 10416 13452 10450
rect 13486 10416 13552 10450
rect 13586 10416 13652 10450
rect 13686 10416 13746 10450
rect 13086 10360 13746 10416
rect -3919 10323 -3913 10357
rect -3879 10323 -3873 10357
rect -3919 10285 -3873 10323
rect -3919 10251 -3913 10285
rect -3879 10251 -3873 10285
rect -3919 10213 -3873 10251
rect -3919 10179 -3913 10213
rect -3879 10179 -3873 10213
rect -3919 10164 -3873 10179
rect -3661 10357 -3615 10359
rect -3661 10323 -3655 10357
rect -3621 10323 -3615 10357
rect -3661 10285 -3615 10323
rect -3661 10251 -3655 10285
rect -3621 10251 -3615 10285
rect -3661 10213 -3615 10251
rect -3661 10179 -3655 10213
rect -3621 10179 -3615 10213
rect -3661 10164 -3615 10179
rect -8765 10126 -8573 10132
rect -8765 10092 -8722 10126
rect -8688 10092 -8650 10126
rect -8616 10092 -8573 10126
rect -8765 10086 -8573 10092
rect -8507 10126 -8315 10132
rect -8507 10092 -8464 10126
rect -8430 10092 -8392 10126
rect -8358 10092 -8315 10126
rect -8507 10086 -8315 10092
rect -8249 10126 -8057 10132
rect -8249 10092 -8206 10126
rect -8172 10092 -8134 10126
rect -8100 10092 -8057 10126
rect -8249 10086 -8057 10092
rect -7991 10126 -7799 10132
rect -7991 10092 -7948 10126
rect -7914 10092 -7876 10126
rect -7842 10092 -7799 10126
rect -7991 10086 -7799 10092
rect -7733 10126 -7541 10132
rect -7733 10092 -7690 10126
rect -7656 10092 -7618 10126
rect -7584 10092 -7541 10126
rect -7733 10086 -7541 10092
rect -7475 10126 -7283 10132
rect -7475 10092 -7432 10126
rect -7398 10092 -7360 10126
rect -7326 10092 -7283 10126
rect -7475 10086 -7283 10092
rect -7217 10126 -7025 10132
rect -7217 10092 -7174 10126
rect -7140 10092 -7102 10126
rect -7068 10092 -7025 10126
rect -7217 10086 -7025 10092
rect -6959 10126 -6767 10132
rect -6959 10092 -6916 10126
rect -6882 10092 -6844 10126
rect -6810 10092 -6767 10126
rect -6959 10086 -6767 10092
rect -6701 10126 -6509 10132
rect -6701 10092 -6658 10126
rect -6624 10092 -6586 10126
rect -6552 10092 -6509 10126
rect -6701 10086 -6509 10092
rect -6443 10126 -6251 10132
rect -6443 10092 -6400 10126
rect -6366 10092 -6328 10126
rect -6294 10092 -6251 10126
rect -6443 10086 -6251 10092
rect -6185 10126 -5993 10132
rect -6185 10092 -6142 10126
rect -6108 10092 -6070 10126
rect -6036 10092 -5993 10126
rect -6185 10086 -5993 10092
rect -5927 10126 -5735 10132
rect -5927 10092 -5884 10126
rect -5850 10092 -5812 10126
rect -5778 10092 -5735 10126
rect -5927 10086 -5735 10092
rect -5669 10126 -5477 10132
rect -5669 10092 -5626 10126
rect -5592 10092 -5554 10126
rect -5520 10092 -5477 10126
rect -5669 10086 -5477 10092
rect -5411 10126 -5219 10132
rect -5411 10092 -5368 10126
rect -5334 10092 -5296 10126
rect -5262 10092 -5219 10126
rect -5411 10086 -5219 10092
rect -5153 10126 -4961 10132
rect -5153 10092 -5110 10126
rect -5076 10092 -5038 10126
rect -5004 10092 -4961 10126
rect -5153 10086 -4961 10092
rect -4895 10126 -4703 10132
rect -4895 10092 -4852 10126
rect -4818 10092 -4780 10126
rect -4746 10092 -4703 10126
rect -4895 10086 -4703 10092
rect -4637 10126 -4445 10132
rect -4637 10092 -4594 10126
rect -4560 10092 -4522 10126
rect -4488 10092 -4445 10126
rect -4637 10086 -4445 10092
rect -4379 10126 -4187 10132
rect -4379 10092 -4336 10126
rect -4302 10092 -4264 10126
rect -4230 10092 -4187 10126
rect -4379 10086 -4187 10092
rect -4121 10126 -3929 10132
rect -4121 10092 -4078 10126
rect -4044 10092 -4006 10126
rect -3972 10092 -3929 10126
rect -4121 10086 -3929 10092
rect -3863 10126 -3671 10132
rect -3863 10092 -3820 10126
rect -3786 10092 -3748 10126
rect -3714 10092 -3671 10126
rect -3863 10086 -3671 10092
rect -9412 10026 -3671 10086
rect -9412 9928 -4750 10026
rect -10054 9882 -4750 9928
rect -9840 9877 -4750 9882
rect -7730 9871 -7482 9877
rect -7730 9837 -7687 9871
rect -7653 9837 -7615 9871
rect -7581 9837 -7482 9871
rect -7730 9831 -7482 9837
rect -7264 9871 -7072 9877
rect -7264 9837 -7221 9871
rect -7187 9837 -7149 9871
rect -7115 9837 -7072 9871
rect -7264 9831 -7072 9837
rect -7006 9871 -6814 9877
rect -7006 9837 -6963 9871
rect -6929 9837 -6891 9871
rect -6857 9837 -6814 9871
rect -7006 9831 -6814 9837
rect -6748 9871 -6556 9877
rect -6748 9837 -6705 9871
rect -6671 9837 -6633 9871
rect -6599 9837 -6556 9871
rect -6748 9831 -6556 9837
rect -6490 9871 -6298 9877
rect -6490 9837 -6447 9871
rect -6413 9837 -6375 9871
rect -6341 9837 -6298 9871
rect -6490 9831 -6298 9837
rect -6232 9871 -6040 9877
rect -6232 9837 -6189 9871
rect -6155 9837 -6117 9871
rect -6083 9837 -6040 9871
rect -6232 9831 -6040 9837
rect -5974 9871 -5782 9877
rect -5974 9837 -5931 9871
rect -5897 9837 -5859 9871
rect -5825 9837 -5782 9871
rect -5974 9831 -5782 9837
rect -5716 9871 -5524 9877
rect -5716 9837 -5673 9871
rect -5639 9837 -5601 9871
rect -5567 9837 -5524 9871
rect -5716 9831 -5524 9837
rect -5458 9871 -5266 9877
rect -5458 9837 -5415 9871
rect -5381 9837 -5343 9871
rect -5309 9837 -5266 9871
rect -5458 9831 -5266 9837
rect -5200 9871 -5008 9877
rect -5200 9837 -5157 9871
rect -5123 9837 -5085 9871
rect -5051 9837 -5008 9871
rect -5200 9831 -5008 9837
rect -4942 9871 -4750 9877
rect -4942 9837 -4899 9871
rect -4865 9837 -4827 9871
rect -4793 9837 -4750 9871
rect -4942 9831 -4750 9837
rect -7786 9788 -7740 9799
rect -7862 9784 -7740 9788
rect -7862 9750 -7780 9784
rect -7746 9750 -7740 9784
rect -7862 9712 -7740 9750
rect -7862 9678 -7780 9712
rect -7746 9678 -7740 9712
rect -7862 9640 -7740 9678
rect -7862 9606 -7780 9640
rect -7746 9606 -7740 9640
rect -7862 9568 -7740 9606
rect -7862 9534 -7780 9568
rect -7746 9534 -7740 9568
rect -7862 9496 -7740 9534
rect -7862 9462 -7780 9496
rect -7746 9462 -7740 9496
rect -7862 9424 -7740 9462
rect -7862 9390 -7780 9424
rect -7746 9390 -7740 9424
rect -7862 9352 -7740 9390
rect -7862 9318 -7780 9352
rect -7746 9318 -7740 9352
rect -7862 9280 -7740 9318
rect -7862 9246 -7780 9280
rect -7746 9246 -7740 9280
rect -7862 9208 -7740 9246
rect -7862 9174 -7780 9208
rect -7746 9174 -7740 9208
rect -7862 9136 -7740 9174
rect -7862 9102 -7780 9136
rect -7746 9102 -7740 9136
rect -7862 9064 -7740 9102
rect -7862 9030 -7780 9064
rect -7746 9030 -7740 9064
rect -7862 8992 -7740 9030
rect -7862 8958 -7780 8992
rect -7746 8958 -7740 8992
rect -7862 8920 -7740 8958
rect -7862 8886 -7780 8920
rect -7746 8886 -7740 8920
rect -7862 8848 -7740 8886
rect -7862 8814 -7780 8848
rect -7746 8814 -7740 8848
rect -7862 8799 -7740 8814
rect -7528 9784 -7482 9831
rect -7528 9750 -7522 9784
rect -7488 9750 -7482 9784
rect -7528 9712 -7482 9750
rect -7528 9678 -7522 9712
rect -7488 9678 -7482 9712
rect -7528 9640 -7482 9678
rect -7528 9606 -7522 9640
rect -7488 9606 -7482 9640
rect -7528 9568 -7482 9606
rect -7528 9534 -7522 9568
rect -7488 9534 -7482 9568
rect -7528 9496 -7482 9534
rect -7528 9462 -7522 9496
rect -7488 9462 -7482 9496
rect -7528 9424 -7482 9462
rect -7528 9390 -7522 9424
rect -7488 9390 -7482 9424
rect -7528 9352 -7482 9390
rect -7528 9318 -7522 9352
rect -7488 9318 -7482 9352
rect -7528 9280 -7482 9318
rect -7528 9246 -7522 9280
rect -7488 9246 -7482 9280
rect -7528 9208 -7482 9246
rect -7528 9174 -7522 9208
rect -7488 9174 -7482 9208
rect -7528 9136 -7482 9174
rect -7320 9784 -7274 9799
rect -7320 9750 -7314 9784
rect -7280 9750 -7274 9784
rect -7320 9712 -7274 9750
rect -7320 9678 -7314 9712
rect -7280 9678 -7274 9712
rect -7320 9640 -7274 9678
rect -7320 9606 -7314 9640
rect -7280 9606 -7274 9640
rect -7320 9568 -7274 9606
rect -7320 9534 -7314 9568
rect -7280 9534 -7274 9568
rect -7320 9496 -7274 9534
rect -7320 9462 -7314 9496
rect -7280 9462 -7274 9496
rect -7062 9784 -7016 9799
rect -7062 9750 -7056 9784
rect -7022 9750 -7016 9784
rect -7062 9712 -7016 9750
rect -7062 9678 -7056 9712
rect -7022 9678 -7016 9712
rect -7062 9640 -7016 9678
rect -7062 9606 -7056 9640
rect -7022 9606 -7016 9640
rect -7062 9568 -7016 9606
rect -7062 9534 -7056 9568
rect -7022 9534 -7016 9568
rect -7062 9496 -7016 9534
rect -7062 9495 -7056 9496
rect -7320 9424 -7274 9462
rect -7320 9390 -7314 9424
rect -7280 9390 -7274 9424
rect -7320 9352 -7274 9390
rect -7320 9318 -7314 9352
rect -7280 9318 -7274 9352
rect -7088 9478 -7056 9495
rect -7022 9495 -7016 9496
rect -6804 9784 -6758 9799
rect -6804 9750 -6798 9784
rect -6764 9750 -6758 9784
rect -6804 9712 -6758 9750
rect -6804 9678 -6798 9712
rect -6764 9678 -6758 9712
rect -6804 9640 -6758 9678
rect -6804 9606 -6798 9640
rect -6764 9606 -6758 9640
rect -6804 9568 -6758 9606
rect -6804 9534 -6798 9568
rect -6764 9534 -6758 9568
rect -6804 9496 -6758 9534
rect -7022 9478 -6991 9495
rect -7088 9426 -7065 9478
rect -7013 9426 -6991 9478
rect -7088 9424 -6991 9426
rect -7088 9414 -7056 9424
rect -7022 9414 -6991 9424
rect -7088 9362 -7065 9414
rect -7013 9362 -6991 9414
rect -7088 9352 -6991 9362
rect -7088 9343 -7056 9352
rect -7320 9280 -7274 9318
rect -7320 9246 -7314 9280
rect -7280 9246 -7274 9280
rect -7320 9208 -7274 9246
rect -7320 9174 -7314 9208
rect -7280 9174 -7274 9208
rect -7320 9164 -7274 9174
rect -7062 9318 -7056 9343
rect -7022 9343 -6991 9352
rect -6804 9462 -6798 9496
rect -6764 9462 -6758 9496
rect -6546 9784 -6500 9799
rect -6546 9750 -6540 9784
rect -6506 9750 -6500 9784
rect -6546 9712 -6500 9750
rect -6546 9678 -6540 9712
rect -6506 9678 -6500 9712
rect -6546 9640 -6500 9678
rect -6546 9606 -6540 9640
rect -6506 9606 -6500 9640
rect -6546 9568 -6500 9606
rect -6546 9534 -6540 9568
rect -6506 9534 -6500 9568
rect -6546 9496 -6500 9534
rect -6546 9495 -6540 9496
rect -6804 9424 -6758 9462
rect -6804 9390 -6798 9424
rect -6764 9390 -6758 9424
rect -6804 9352 -6758 9390
rect -7022 9318 -7016 9343
rect -7062 9280 -7016 9318
rect -7062 9246 -7056 9280
rect -7022 9246 -7016 9280
rect -7062 9208 -7016 9246
rect -7062 9174 -7056 9208
rect -7022 9174 -7016 9208
rect -7528 9102 -7522 9136
rect -7488 9102 -7482 9136
rect -7528 9064 -7482 9102
rect -7528 9030 -7522 9064
rect -7488 9030 -7482 9064
rect -7528 8992 -7482 9030
rect -7528 8958 -7522 8992
rect -7488 8958 -7482 8992
rect -7335 9136 -7257 9164
rect -7335 9128 -7314 9136
rect -7280 9128 -7257 9136
rect -7335 9076 -7322 9128
rect -7270 9076 -7257 9128
rect -7335 9064 -7257 9076
rect -7335 9012 -7322 9064
rect -7270 9012 -7257 9064
rect -7335 8992 -7257 9012
rect -7335 8979 -7314 8992
rect -7528 8920 -7482 8958
rect -7528 8886 -7522 8920
rect -7488 8886 -7482 8920
rect -7528 8848 -7482 8886
rect -7528 8814 -7522 8848
rect -7488 8814 -7482 8848
rect -7862 7700 -7778 8799
rect -7528 8767 -7482 8814
rect -7320 8958 -7314 8979
rect -7280 8979 -7257 8992
rect -7062 9136 -7016 9174
rect -6804 9318 -6798 9352
rect -6764 9318 -6758 9352
rect -6565 9475 -6540 9495
rect -6506 9495 -6500 9496
rect -6288 9784 -6242 9799
rect -6288 9750 -6282 9784
rect -6248 9750 -6242 9784
rect -6288 9712 -6242 9750
rect -6288 9678 -6282 9712
rect -6248 9678 -6242 9712
rect -6288 9640 -6242 9678
rect -6288 9606 -6282 9640
rect -6248 9606 -6242 9640
rect -6288 9568 -6242 9606
rect -6288 9534 -6282 9568
rect -6248 9534 -6242 9568
rect -6288 9496 -6242 9534
rect -6506 9475 -6481 9495
rect -6565 9423 -6549 9475
rect -6497 9423 -6481 9475
rect -6565 9411 -6540 9423
rect -6506 9411 -6481 9423
rect -6565 9359 -6549 9411
rect -6497 9359 -6481 9411
rect -6565 9352 -6481 9359
rect -6565 9343 -6540 9352
rect -6804 9280 -6758 9318
rect -6804 9246 -6798 9280
rect -6764 9246 -6758 9280
rect -6804 9208 -6758 9246
rect -6804 9174 -6798 9208
rect -6764 9174 -6758 9208
rect -6804 9164 -6758 9174
rect -6546 9318 -6540 9343
rect -6506 9343 -6481 9352
rect -6288 9462 -6282 9496
rect -6248 9462 -6242 9496
rect -6030 9784 -5984 9799
rect -6030 9750 -6024 9784
rect -5990 9750 -5984 9784
rect -6030 9712 -5984 9750
rect -6030 9678 -6024 9712
rect -5990 9678 -5984 9712
rect -6030 9640 -5984 9678
rect -6030 9606 -6024 9640
rect -5990 9606 -5984 9640
rect -6030 9568 -5984 9606
rect -6030 9534 -6024 9568
rect -5990 9534 -5984 9568
rect -6030 9496 -5984 9534
rect -6030 9495 -6024 9496
rect -6288 9424 -6242 9462
rect -6288 9390 -6282 9424
rect -6248 9390 -6242 9424
rect -6288 9352 -6242 9390
rect -6506 9318 -6500 9343
rect -6546 9280 -6500 9318
rect -6546 9246 -6540 9280
rect -6506 9246 -6500 9280
rect -6546 9208 -6500 9246
rect -6546 9174 -6540 9208
rect -6506 9174 -6500 9208
rect -7062 9102 -7056 9136
rect -7022 9102 -7016 9136
rect -7062 9064 -7016 9102
rect -7062 9030 -7056 9064
rect -7022 9030 -7016 9064
rect -7062 8992 -7016 9030
rect -7280 8958 -7274 8979
rect -7320 8920 -7274 8958
rect -7320 8886 -7314 8920
rect -7280 8886 -7274 8920
rect -7320 8848 -7274 8886
rect -7320 8814 -7314 8848
rect -7280 8814 -7274 8848
rect -7320 8799 -7274 8814
rect -7062 8958 -7056 8992
rect -7022 8958 -7016 8992
rect -6821 9136 -6737 9164
rect -6821 9127 -6798 9136
rect -6764 9127 -6737 9136
rect -6821 9075 -6805 9127
rect -6753 9075 -6737 9127
rect -6821 9064 -6737 9075
rect -6821 9063 -6798 9064
rect -6764 9063 -6737 9064
rect -6821 9011 -6805 9063
rect -6753 9011 -6737 9063
rect -6821 8992 -6737 9011
rect -6821 8979 -6798 8992
rect -7062 8920 -7016 8958
rect -7062 8886 -7056 8920
rect -7022 8886 -7016 8920
rect -7062 8848 -7016 8886
rect -7062 8814 -7056 8848
rect -7022 8814 -7016 8848
rect -7062 8799 -7016 8814
rect -6804 8958 -6798 8979
rect -6764 8979 -6737 8992
rect -6546 9136 -6500 9174
rect -6288 9318 -6282 9352
rect -6248 9318 -6242 9352
rect -6050 9477 -6024 9495
rect -5990 9495 -5984 9496
rect -5772 9784 -5726 9799
rect -5772 9750 -5766 9784
rect -5732 9750 -5726 9784
rect -5772 9712 -5726 9750
rect -5772 9678 -5766 9712
rect -5732 9678 -5726 9712
rect -5772 9640 -5726 9678
rect -5772 9606 -5766 9640
rect -5732 9606 -5726 9640
rect -5772 9568 -5726 9606
rect -5772 9534 -5766 9568
rect -5732 9534 -5726 9568
rect -5772 9496 -5726 9534
rect -5990 9477 -5962 9495
rect -6050 9425 -6033 9477
rect -5981 9425 -5962 9477
rect -6050 9424 -5962 9425
rect -6050 9413 -6024 9424
rect -5990 9413 -5962 9424
rect -6050 9361 -6033 9413
rect -5981 9361 -5962 9413
rect -6050 9352 -5962 9361
rect -6050 9343 -6024 9352
rect -6288 9280 -6242 9318
rect -6288 9246 -6282 9280
rect -6248 9246 -6242 9280
rect -6288 9208 -6242 9246
rect -6288 9174 -6282 9208
rect -6248 9174 -6242 9208
rect -6288 9164 -6242 9174
rect -6030 9318 -6024 9343
rect -5990 9343 -5962 9352
rect -5772 9462 -5766 9496
rect -5732 9462 -5726 9496
rect -5514 9784 -5468 9799
rect -5514 9750 -5508 9784
rect -5474 9750 -5468 9784
rect -5514 9712 -5468 9750
rect -5514 9678 -5508 9712
rect -5474 9678 -5468 9712
rect -5514 9640 -5468 9678
rect -5514 9606 -5508 9640
rect -5474 9606 -5468 9640
rect -5514 9568 -5468 9606
rect -5514 9534 -5508 9568
rect -5474 9534 -5468 9568
rect -5514 9496 -5468 9534
rect -5514 9495 -5508 9496
rect -5772 9424 -5726 9462
rect -5772 9390 -5766 9424
rect -5732 9390 -5726 9424
rect -5772 9352 -5726 9390
rect -5990 9318 -5984 9343
rect -6030 9280 -5984 9318
rect -6030 9246 -6024 9280
rect -5990 9246 -5984 9280
rect -6030 9208 -5984 9246
rect -6030 9174 -6024 9208
rect -5990 9174 -5984 9208
rect -6546 9102 -6540 9136
rect -6506 9102 -6500 9136
rect -6546 9064 -6500 9102
rect -6546 9030 -6540 9064
rect -6506 9030 -6500 9064
rect -6546 8992 -6500 9030
rect -6764 8958 -6758 8979
rect -6804 8920 -6758 8958
rect -6804 8886 -6798 8920
rect -6764 8886 -6758 8920
rect -6804 8848 -6758 8886
rect -6804 8814 -6798 8848
rect -6764 8814 -6758 8848
rect -6804 8799 -6758 8814
rect -6546 8958 -6540 8992
rect -6506 8958 -6500 8992
rect -6308 9136 -6223 9164
rect -6308 9129 -6282 9136
rect -6248 9129 -6223 9136
rect -6308 9077 -6292 9129
rect -6240 9077 -6223 9129
rect -6308 9065 -6223 9077
rect -6308 9013 -6292 9065
rect -6240 9013 -6223 9065
rect -6308 8992 -6223 9013
rect -6308 8979 -6282 8992
rect -6546 8920 -6500 8958
rect -6546 8886 -6540 8920
rect -6506 8886 -6500 8920
rect -6546 8848 -6500 8886
rect -6546 8814 -6540 8848
rect -6506 8814 -6500 8848
rect -6546 8799 -6500 8814
rect -6288 8958 -6282 8979
rect -6248 8979 -6223 8992
rect -6030 9136 -5984 9174
rect -5772 9318 -5766 9352
rect -5732 9318 -5726 9352
rect -5531 9475 -5508 9495
rect -5474 9495 -5468 9496
rect -5256 9784 -5210 9799
rect -5256 9750 -5250 9784
rect -5216 9750 -5210 9784
rect -5256 9712 -5210 9750
rect -5256 9678 -5250 9712
rect -5216 9678 -5210 9712
rect -5256 9640 -5210 9678
rect -5256 9606 -5250 9640
rect -5216 9606 -5210 9640
rect -5256 9568 -5210 9606
rect -5256 9534 -5250 9568
rect -5216 9534 -5210 9568
rect -5256 9496 -5210 9534
rect -5474 9475 -5449 9495
rect -5531 9423 -5516 9475
rect -5464 9423 -5449 9475
rect -5531 9411 -5508 9423
rect -5474 9411 -5449 9423
rect -5531 9359 -5516 9411
rect -5464 9359 -5449 9411
rect -5531 9352 -5449 9359
rect -5531 9343 -5508 9352
rect -5772 9280 -5726 9318
rect -5772 9246 -5766 9280
rect -5732 9246 -5726 9280
rect -5772 9208 -5726 9246
rect -5772 9174 -5766 9208
rect -5732 9174 -5726 9208
rect -5772 9164 -5726 9174
rect -5514 9318 -5508 9343
rect -5474 9343 -5449 9352
rect -5256 9462 -5250 9496
rect -5216 9462 -5210 9496
rect -4998 9784 -4952 9799
rect -4998 9750 -4992 9784
rect -4958 9750 -4952 9784
rect -4998 9712 -4952 9750
rect -4998 9678 -4992 9712
rect -4958 9678 -4952 9712
rect -4998 9640 -4952 9678
rect -4998 9606 -4992 9640
rect -4958 9606 -4952 9640
rect -4998 9568 -4952 9606
rect -4998 9534 -4992 9568
rect -4958 9534 -4952 9568
rect -4998 9496 -4952 9534
rect -4998 9495 -4992 9496
rect -5256 9424 -5210 9462
rect -5256 9390 -5250 9424
rect -5216 9390 -5210 9424
rect -5256 9352 -5210 9390
rect -5474 9318 -5468 9343
rect -5514 9280 -5468 9318
rect -5514 9246 -5508 9280
rect -5474 9246 -5468 9280
rect -5514 9208 -5468 9246
rect -5514 9174 -5508 9208
rect -5474 9174 -5468 9208
rect -6030 9102 -6024 9136
rect -5990 9102 -5984 9136
rect -6030 9064 -5984 9102
rect -6030 9030 -6024 9064
rect -5990 9030 -5984 9064
rect -6030 8992 -5984 9030
rect -6248 8958 -6242 8979
rect -6288 8920 -6242 8958
rect -6288 8886 -6282 8920
rect -6248 8886 -6242 8920
rect -6288 8848 -6242 8886
rect -6288 8814 -6282 8848
rect -6248 8814 -6242 8848
rect -6288 8799 -6242 8814
rect -6030 8958 -6024 8992
rect -5990 8958 -5984 8992
rect -5789 9136 -5706 9164
rect -5789 9128 -5766 9136
rect -5732 9128 -5706 9136
rect -5789 9076 -5774 9128
rect -5722 9076 -5706 9128
rect -5789 9064 -5706 9076
rect -5789 9012 -5774 9064
rect -5722 9012 -5706 9064
rect -5789 8992 -5706 9012
rect -5789 8979 -5766 8992
rect -6030 8920 -5984 8958
rect -6030 8886 -6024 8920
rect -5990 8886 -5984 8920
rect -6030 8848 -5984 8886
rect -6030 8814 -6024 8848
rect -5990 8814 -5984 8848
rect -6030 8799 -5984 8814
rect -5772 8958 -5766 8979
rect -5732 8979 -5706 8992
rect -5514 9136 -5468 9174
rect -5256 9318 -5250 9352
rect -5216 9318 -5210 9352
rect -5017 9476 -4992 9495
rect -4958 9495 -4952 9496
rect -4740 9784 -4694 9799
rect -4740 9750 -4734 9784
rect -4700 9750 -4694 9784
rect -4740 9712 -4694 9750
rect -4740 9678 -4734 9712
rect -4700 9678 -4694 9712
rect -4740 9640 -4694 9678
rect -4740 9606 -4734 9640
rect -4700 9606 -4694 9640
rect -4740 9568 -4694 9606
rect -4740 9534 -4734 9568
rect -4700 9534 -4694 9568
rect -4740 9496 -4694 9534
rect -4958 9476 -4930 9495
rect -5017 9424 -5002 9476
rect -4950 9424 -4930 9476
rect -5017 9412 -4992 9424
rect -4958 9412 -4930 9424
rect -5017 9360 -5002 9412
rect -4950 9360 -4930 9412
rect -5017 9352 -4930 9360
rect -5017 9343 -4992 9352
rect -5256 9280 -5210 9318
rect -5256 9246 -5250 9280
rect -5216 9246 -5210 9280
rect -5256 9208 -5210 9246
rect -5256 9174 -5250 9208
rect -5216 9174 -5210 9208
rect -5256 9164 -5210 9174
rect -4998 9318 -4992 9343
rect -4958 9343 -4930 9352
rect -4740 9462 -4734 9496
rect -4700 9462 -4694 9496
rect -4740 9424 -4694 9462
rect -4740 9390 -4734 9424
rect -4700 9390 -4694 9424
rect -4740 9352 -4694 9390
rect -4958 9318 -4952 9343
rect -4998 9280 -4952 9318
rect -4998 9246 -4992 9280
rect -4958 9246 -4952 9280
rect -4998 9208 -4952 9246
rect -4998 9174 -4992 9208
rect -4958 9174 -4952 9208
rect -5514 9102 -5508 9136
rect -5474 9102 -5468 9136
rect -5514 9064 -5468 9102
rect -5514 9030 -5508 9064
rect -5474 9030 -5468 9064
rect -5514 8992 -5468 9030
rect -5732 8958 -5726 8979
rect -5772 8920 -5726 8958
rect -5772 8886 -5766 8920
rect -5732 8886 -5726 8920
rect -5772 8848 -5726 8886
rect -5772 8814 -5766 8848
rect -5732 8814 -5726 8848
rect -5772 8799 -5726 8814
rect -5514 8958 -5508 8992
rect -5474 8958 -5468 8992
rect -5277 9136 -5186 9164
rect -5277 9128 -5250 9136
rect -5216 9128 -5186 9136
rect -5277 9076 -5257 9128
rect -5205 9076 -5186 9128
rect -5277 9064 -5186 9076
rect -5277 9012 -5257 9064
rect -5205 9012 -5186 9064
rect -5277 8992 -5186 9012
rect -5277 8979 -5250 8992
rect -5514 8920 -5468 8958
rect -5514 8886 -5508 8920
rect -5474 8886 -5468 8920
rect -5514 8848 -5468 8886
rect -5514 8814 -5508 8848
rect -5474 8814 -5468 8848
rect -5514 8799 -5468 8814
rect -5256 8958 -5250 8979
rect -5216 8979 -5186 8992
rect -4998 9136 -4952 9174
rect -4740 9318 -4734 9352
rect -4700 9318 -4694 9352
rect -4740 9280 -4694 9318
rect -4740 9246 -4734 9280
rect -4700 9246 -4694 9280
rect -4740 9208 -4694 9246
rect -4740 9174 -4734 9208
rect -4700 9174 -4694 9208
rect -4740 9164 -4694 9174
rect 13086 9460 13766 9560
rect 13086 9426 13152 9460
rect 13186 9426 13252 9460
rect 13286 9426 13352 9460
rect 13386 9426 13452 9460
rect 13486 9426 13552 9460
rect 13586 9426 13652 9460
rect 13686 9426 13766 9460
rect 13086 9360 13766 9426
rect 13086 9326 13152 9360
rect 13186 9326 13252 9360
rect 13286 9356 13352 9360
rect 13386 9356 13452 9360
rect 13486 9356 13552 9360
rect 13586 9326 13652 9360
rect 13686 9326 13766 9360
rect 13086 9260 13262 9326
rect 13570 9260 13766 9326
rect 13086 9226 13152 9260
rect 13186 9226 13252 9260
rect 13586 9226 13652 9260
rect 13686 9226 13766 9260
rect -4998 9102 -4992 9136
rect -4958 9102 -4952 9136
rect -4998 9064 -4952 9102
rect -4998 9030 -4992 9064
rect -4958 9030 -4952 9064
rect -4998 8992 -4952 9030
rect -5216 8958 -5210 8979
rect -5256 8920 -5210 8958
rect -5256 8886 -5250 8920
rect -5216 8886 -5210 8920
rect -5256 8848 -5210 8886
rect -5256 8814 -5250 8848
rect -5216 8814 -5210 8848
rect -5256 8799 -5210 8814
rect -4998 8958 -4992 8992
rect -4958 8958 -4952 8992
rect -4761 9136 -4673 9164
rect -4761 9129 -4734 9136
rect -4700 9129 -4673 9136
rect -4761 9077 -4742 9129
rect -4690 9077 -4673 9129
rect -4761 9065 -4673 9077
rect -4761 9013 -4742 9065
rect -4690 9013 -4673 9065
rect -4761 8992 -4673 9013
rect -4761 8978 -4734 8992
rect -4998 8920 -4952 8958
rect -4998 8886 -4992 8920
rect -4958 8886 -4952 8920
rect -4998 8848 -4952 8886
rect -4998 8814 -4992 8848
rect -4958 8814 -4952 8848
rect -4998 8799 -4952 8814
rect -4740 8958 -4734 8978
rect -4700 8978 -4673 8992
rect 13086 9160 13262 9226
rect 13570 9160 13766 9226
rect 13086 9126 13152 9160
rect 13186 9126 13252 9160
rect 13586 9126 13652 9160
rect 13686 9126 13766 9160
rect 13086 9060 13262 9126
rect 13570 9060 13766 9126
rect 13086 9026 13152 9060
rect 13186 9026 13252 9060
rect 13286 9026 13352 9048
rect 13386 9026 13452 9048
rect 13486 9026 13552 9048
rect 13586 9026 13652 9060
rect 13686 9026 13766 9060
rect -4700 8958 -4694 8978
rect -4740 8920 -4694 8958
rect -4740 8886 -4734 8920
rect -4700 8886 -4694 8920
rect -4740 8848 -4694 8886
rect 13086 8960 13766 9026
rect 13086 8926 13152 8960
rect 13186 8926 13252 8960
rect 13286 8926 13352 8960
rect 13386 8926 13452 8960
rect 13486 8926 13552 8960
rect 13586 8926 13652 8960
rect 13686 8926 13766 8960
rect 13086 8860 13766 8926
rect -4740 8814 -4734 8848
rect -4700 8814 -4694 8848
rect -4740 8799 -4694 8814
rect -7730 8761 -7482 8767
rect -7730 8727 -7687 8761
rect -7653 8727 -7615 8761
rect -7581 8727 -7482 8761
rect -7730 8721 -7482 8727
rect -7264 8761 -7072 8767
rect -7264 8727 -7221 8761
rect -7187 8727 -7149 8761
rect -7115 8727 -7072 8761
rect -7264 8721 -7072 8727
rect -7006 8761 -6814 8767
rect -7006 8727 -6963 8761
rect -6929 8727 -6891 8761
rect -6857 8727 -6814 8761
rect -7006 8721 -6814 8727
rect -6748 8761 -6556 8767
rect -6748 8727 -6705 8761
rect -6671 8727 -6633 8761
rect -6599 8727 -6556 8761
rect -6748 8721 -6556 8727
rect -6490 8761 -6298 8767
rect -6490 8727 -6447 8761
rect -6413 8727 -6375 8761
rect -6341 8727 -6298 8761
rect -6490 8721 -6298 8727
rect -6232 8761 -6040 8767
rect -6232 8727 -6189 8761
rect -6155 8727 -6117 8761
rect -6083 8727 -6040 8761
rect -6232 8721 -6040 8727
rect -5974 8761 -5782 8767
rect -5974 8727 -5931 8761
rect -5897 8727 -5859 8761
rect -5825 8727 -5782 8761
rect -5974 8721 -5782 8727
rect -5716 8761 -5524 8767
rect -5716 8727 -5673 8761
rect -5639 8727 -5601 8761
rect -5567 8727 -5524 8761
rect -5716 8721 -5524 8727
rect -5458 8761 -5266 8767
rect -5458 8727 -5415 8761
rect -5381 8727 -5343 8761
rect -5309 8727 -5266 8761
rect -5458 8721 -5266 8727
rect -5200 8761 -5008 8767
rect -5200 8727 -5157 8761
rect -5123 8727 -5085 8761
rect -5051 8727 -5008 8761
rect -5200 8721 -5008 8727
rect -4942 8761 -4750 8767
rect -4942 8727 -4899 8761
rect -4865 8727 -4827 8761
rect -4793 8727 -4750 8761
rect -4942 8721 -4750 8727
rect -7730 8658 -4750 8721
rect 13111 8050 13721 8095
rect 13111 8016 13142 8050
rect 13176 8016 13242 8050
rect 13276 8016 13342 8050
rect 13376 8016 13442 8050
rect 13476 8016 13542 8050
rect 13576 8016 13642 8050
rect 13676 8016 13721 8050
rect 13111 7950 13721 8016
rect 13111 7916 13142 7950
rect 13176 7916 13242 7950
rect 13276 7916 13342 7950
rect 13376 7916 13442 7950
rect 13476 7916 13542 7950
rect 13576 7916 13642 7950
rect 13676 7916 13721 7950
rect 13111 7850 13721 7916
rect 13111 7816 13142 7850
rect 13176 7816 13242 7850
rect 13276 7816 13342 7850
rect 13376 7816 13442 7850
rect 13476 7816 13542 7850
rect 13576 7816 13642 7850
rect 13676 7816 13721 7850
rect 13111 7750 13721 7816
rect 14462 7980 14682 11680
rect 16922 11391 17052 11430
rect 15852 11334 16202 11360
rect 16922 11339 16956 11391
rect 17008 11339 17052 11391
rect 16922 11334 17052 11339
rect 15004 11328 17054 11334
rect 15004 11294 15051 11328
rect 15085 11294 15123 11328
rect 15157 11294 15195 11328
rect 15229 11294 15267 11328
rect 15301 11294 15339 11328
rect 15373 11294 15411 11328
rect 15445 11294 15483 11328
rect 15517 11294 15555 11328
rect 15589 11294 15627 11328
rect 15661 11294 15699 11328
rect 15733 11294 15771 11328
rect 15805 11294 15843 11328
rect 15877 11294 15915 11328
rect 15949 11294 16109 11328
rect 16143 11294 16181 11328
rect 16215 11294 16253 11328
rect 16287 11294 16325 11328
rect 16359 11294 16397 11328
rect 16431 11294 16469 11328
rect 16503 11294 16541 11328
rect 16575 11294 16613 11328
rect 16647 11294 16685 11328
rect 16719 11294 16757 11328
rect 16791 11294 16829 11328
rect 16863 11294 16901 11328
rect 16935 11294 16973 11328
rect 17007 11294 17054 11328
rect 15004 11290 17054 11294
rect 15004 11288 15996 11290
rect 16062 11288 17054 11290
rect 14948 11204 14994 11247
rect 16006 11240 16052 11247
rect 14948 11170 14954 11204
rect 14988 11170 14994 11204
rect 14948 11132 14994 11170
rect 14948 11098 14954 11132
rect 14988 11098 14994 11132
rect 14948 11060 14994 11098
rect 14948 11026 14954 11060
rect 14988 11026 14994 11060
rect 14948 10988 14994 11026
rect 14948 10954 14954 10988
rect 14988 10954 14994 10988
rect 14948 10916 14994 10954
rect 14948 10882 14954 10916
rect 14988 10882 14994 10916
rect 15942 11204 16162 11240
rect 17064 11230 17110 11247
rect 17162 11230 17292 11690
rect 18032 11680 18635 11690
rect 18669 11680 18707 11714
rect 18741 11680 18779 11714
rect 18813 11680 18851 11714
rect 18885 11680 18923 11714
rect 18957 11680 18995 11714
rect 19029 11680 19067 11714
rect 19101 11680 19139 11714
rect 19173 11680 19211 11714
rect 19245 11680 19283 11714
rect 19317 11680 19355 11714
rect 19389 11680 19427 11714
rect 19461 11680 19499 11714
rect 19533 11680 19580 11714
rect 18032 11674 19580 11680
rect 18032 11590 18776 11674
rect 18276 11574 18776 11590
rect 17572 11414 17722 11434
rect 17536 11376 17966 11414
rect 17536 11324 17626 11376
rect 17678 11324 17966 11376
rect 17536 11308 17966 11324
rect 17528 11304 18520 11308
rect 18586 11304 19578 11308
rect 17528 11302 19578 11304
rect 17528 11268 17575 11302
rect 17609 11268 17647 11302
rect 17681 11268 17719 11302
rect 17753 11268 17791 11302
rect 17825 11268 17863 11302
rect 17897 11268 17935 11302
rect 17969 11268 18007 11302
rect 18041 11268 18079 11302
rect 18113 11268 18151 11302
rect 18185 11268 18223 11302
rect 18257 11268 18295 11302
rect 18329 11268 18367 11302
rect 18401 11268 18439 11302
rect 18473 11268 18633 11302
rect 18667 11268 18705 11302
rect 18739 11268 18777 11302
rect 18811 11268 18849 11302
rect 18883 11268 18921 11302
rect 18955 11268 18993 11302
rect 19027 11268 19065 11302
rect 19099 11268 19137 11302
rect 19171 11268 19209 11302
rect 19243 11268 19281 11302
rect 19315 11268 19353 11302
rect 19387 11268 19425 11302
rect 19459 11268 19497 11302
rect 19531 11268 19578 11302
rect 17528 11264 19578 11268
rect 17528 11262 18520 11264
rect 18586 11262 19578 11264
rect 15942 11182 16012 11204
rect 16046 11182 16162 11204
rect 15942 10938 15989 11182
rect 16105 10938 16162 11182
rect 17052 11204 17292 11230
rect 19894 11222 20250 13428
rect 17052 11170 17070 11204
rect 17104 11170 17292 11204
rect 17052 11132 17292 11170
rect 17052 11098 17070 11132
rect 17104 11098 17292 11132
rect 17052 11060 17292 11098
rect 17052 11050 17070 11060
rect 15942 10916 16162 10938
rect 15942 10890 16012 10916
rect 14948 10844 14994 10882
rect 14948 10810 14954 10844
rect 14988 10810 14994 10844
rect 14948 10772 14994 10810
rect 14948 10738 14954 10772
rect 14988 10738 14994 10772
rect 14948 10700 14994 10738
rect 14948 10666 14954 10700
rect 14988 10666 14994 10700
rect 14948 10628 14994 10666
rect 14948 10594 14954 10628
rect 14988 10594 14994 10628
rect 14948 10556 14994 10594
rect 14948 10522 14954 10556
rect 14988 10522 14994 10556
rect 14948 10484 14994 10522
rect 14948 10450 14954 10484
rect 14988 10450 14994 10484
rect 14948 10412 14994 10450
rect 14948 10378 14954 10412
rect 14988 10378 14994 10412
rect 14948 10340 14994 10378
rect 14948 10306 14954 10340
rect 14988 10306 14994 10340
rect 14948 10268 14994 10306
rect 14948 10234 14954 10268
rect 14988 10234 14994 10268
rect 14948 10196 14994 10234
rect 14948 10162 14954 10196
rect 14988 10162 14994 10196
rect 14948 10124 14994 10162
rect 14948 10090 14954 10124
rect 14988 10090 14994 10124
rect 14948 10052 14994 10090
rect 14948 10018 14954 10052
rect 14988 10018 14994 10052
rect 14948 9980 14994 10018
rect 14948 9946 14954 9980
rect 14988 9946 14994 9980
rect 14948 9908 14994 9946
rect 14948 9874 14954 9908
rect 14988 9874 14994 9908
rect 14948 9836 14994 9874
rect 14948 9802 14954 9836
rect 14988 9802 14994 9836
rect 14948 9764 14994 9802
rect 14948 9730 14954 9764
rect 14988 9730 14994 9764
rect 14948 9692 14994 9730
rect 14948 9658 14954 9692
rect 14988 9658 14994 9692
rect 14948 9620 14994 9658
rect 14948 9586 14954 9620
rect 14988 9586 14994 9620
rect 14948 9548 14994 9586
rect 14948 9514 14954 9548
rect 14988 9514 14994 9548
rect 14948 9476 14994 9514
rect 14948 9442 14954 9476
rect 14988 9442 14994 9476
rect 14948 9404 14994 9442
rect 14948 9370 14954 9404
rect 14988 9370 14994 9404
rect 14948 9332 14994 9370
rect 14948 9298 14954 9332
rect 14988 9298 14994 9332
rect 14948 9260 14994 9298
rect 14948 9226 14954 9260
rect 14988 9226 14994 9260
rect 14948 9188 14994 9226
rect 14948 9154 14954 9188
rect 14988 9154 14994 9188
rect 14948 9116 14994 9154
rect 14948 9082 14954 9116
rect 14988 9082 14994 9116
rect 14948 9044 14994 9082
rect 14948 9010 14954 9044
rect 14988 9010 14994 9044
rect 14948 8972 14994 9010
rect 14948 8938 14954 8972
rect 14988 8938 14994 8972
rect 14948 8900 14994 8938
rect 14948 8866 14954 8900
rect 14988 8866 14994 8900
rect 14948 8828 14994 8866
rect 14948 8794 14954 8828
rect 14988 8794 14994 8828
rect 14948 8756 14994 8794
rect 14948 8722 14954 8756
rect 14988 8722 14994 8756
rect 14948 8700 14994 8722
rect 16006 10882 16012 10890
rect 16046 10890 16162 10916
rect 17064 11026 17070 11050
rect 17104 11050 17292 11060
rect 17472 11178 17518 11221
rect 17472 11144 17478 11178
rect 17512 11144 17518 11178
rect 18530 11178 18576 11221
rect 18530 11174 18536 11178
rect 17472 11106 17518 11144
rect 17472 11072 17478 11106
rect 17512 11072 17518 11106
rect 17104 11026 17110 11050
rect 17064 10988 17110 11026
rect 17064 10954 17070 10988
rect 17104 10954 17110 10988
rect 17064 10916 17110 10954
rect 16046 10882 16052 10890
rect 16006 10844 16052 10882
rect 16006 10810 16012 10844
rect 16046 10810 16052 10844
rect 16006 10772 16052 10810
rect 16006 10738 16012 10772
rect 16046 10738 16052 10772
rect 16006 10700 16052 10738
rect 16006 10666 16012 10700
rect 16046 10666 16052 10700
rect 16006 10628 16052 10666
rect 16006 10594 16012 10628
rect 16046 10594 16052 10628
rect 16006 10556 16052 10594
rect 16006 10522 16012 10556
rect 16046 10522 16052 10556
rect 16006 10484 16052 10522
rect 16006 10450 16012 10484
rect 16046 10450 16052 10484
rect 16006 10412 16052 10450
rect 16006 10378 16012 10412
rect 16046 10378 16052 10412
rect 16006 10340 16052 10378
rect 16006 10306 16012 10340
rect 16046 10306 16052 10340
rect 16006 10268 16052 10306
rect 16006 10234 16012 10268
rect 16046 10234 16052 10268
rect 16006 10196 16052 10234
rect 16006 10162 16012 10196
rect 16046 10162 16052 10196
rect 16006 10124 16052 10162
rect 16006 10090 16012 10124
rect 16046 10090 16052 10124
rect 16006 10052 16052 10090
rect 16006 10018 16012 10052
rect 16046 10018 16052 10052
rect 16006 9980 16052 10018
rect 16006 9946 16012 9980
rect 16046 9946 16052 9980
rect 16006 9908 16052 9946
rect 16006 9874 16012 9908
rect 16046 9874 16052 9908
rect 16006 9836 16052 9874
rect 16006 9802 16012 9836
rect 16046 9802 16052 9836
rect 16006 9764 16052 9802
rect 16006 9730 16012 9764
rect 16046 9730 16052 9764
rect 16006 9692 16052 9730
rect 16006 9658 16012 9692
rect 16046 9658 16052 9692
rect 16006 9620 16052 9658
rect 16006 9586 16012 9620
rect 16046 9586 16052 9620
rect 16006 9548 16052 9586
rect 16006 9514 16012 9548
rect 16046 9514 16052 9548
rect 16006 9476 16052 9514
rect 16006 9442 16012 9476
rect 16046 9442 16052 9476
rect 16006 9404 16052 9442
rect 16006 9370 16012 9404
rect 16046 9370 16052 9404
rect 16006 9332 16052 9370
rect 16006 9298 16012 9332
rect 16046 9298 16052 9332
rect 16006 9260 16052 9298
rect 16006 9226 16012 9260
rect 16046 9226 16052 9260
rect 16006 9188 16052 9226
rect 16006 9154 16012 9188
rect 16046 9154 16052 9188
rect 16006 9116 16052 9154
rect 16006 9082 16012 9116
rect 16046 9082 16052 9116
rect 16006 9044 16052 9082
rect 16006 9010 16012 9044
rect 16046 9010 16052 9044
rect 16006 8972 16052 9010
rect 16006 8938 16012 8972
rect 16046 8938 16052 8972
rect 16006 8900 16052 8938
rect 16006 8866 16012 8900
rect 16046 8866 16052 8900
rect 16006 8828 16052 8866
rect 16006 8794 16012 8828
rect 16046 8794 16052 8828
rect 16006 8756 16052 8794
rect 16006 8722 16012 8756
rect 16046 8722 16052 8756
rect 14932 8684 15142 8700
rect 14932 8650 14954 8684
rect 14988 8676 15142 8684
rect 14932 8612 14979 8650
rect 14932 8578 14954 8612
rect 14932 8540 14979 8578
rect 14932 8506 14954 8540
rect 14932 8468 14979 8506
rect 14932 8434 14954 8468
rect 14932 8396 14979 8434
rect 14932 8362 14954 8396
rect 14932 8324 14979 8362
rect 14932 8290 14954 8324
rect 15095 8304 15142 8676
rect 14988 8290 15142 8304
rect 14932 8270 15142 8290
rect 16006 8684 16052 8722
rect 17064 10882 17070 10916
rect 17104 10882 17110 10916
rect 17064 10844 17110 10882
rect 17064 10810 17070 10844
rect 17104 10810 17110 10844
rect 17064 10772 17110 10810
rect 17064 10738 17070 10772
rect 17104 10738 17110 10772
rect 17064 10700 17110 10738
rect 17064 10666 17070 10700
rect 17104 10666 17110 10700
rect 17064 10628 17110 10666
rect 17064 10594 17070 10628
rect 17104 10594 17110 10628
rect 17064 10556 17110 10594
rect 17064 10522 17070 10556
rect 17104 10522 17110 10556
rect 17064 10484 17110 10522
rect 17064 10450 17070 10484
rect 17104 10450 17110 10484
rect 17064 10412 17110 10450
rect 17064 10378 17070 10412
rect 17104 10378 17110 10412
rect 17064 10340 17110 10378
rect 17064 10306 17070 10340
rect 17104 10306 17110 10340
rect 17064 10268 17110 10306
rect 17064 10234 17070 10268
rect 17104 10234 17110 10268
rect 17064 10196 17110 10234
rect 17064 10162 17070 10196
rect 17104 10162 17110 10196
rect 17064 10124 17110 10162
rect 17064 10090 17070 10124
rect 17104 10090 17110 10124
rect 17064 10052 17110 10090
rect 17064 10018 17070 10052
rect 17104 10018 17110 10052
rect 17064 9980 17110 10018
rect 17064 9946 17070 9980
rect 17104 9946 17110 9980
rect 17064 9908 17110 9946
rect 17064 9874 17070 9908
rect 17104 9874 17110 9908
rect 17064 9836 17110 9874
rect 17064 9802 17070 9836
rect 17104 9802 17110 9836
rect 17064 9764 17110 9802
rect 17064 9730 17070 9764
rect 17104 9730 17110 9764
rect 17064 9692 17110 9730
rect 17064 9658 17070 9692
rect 17104 9658 17110 9692
rect 17064 9620 17110 9658
rect 17064 9586 17070 9620
rect 17104 9586 17110 9620
rect 17064 9548 17110 9586
rect 17064 9514 17070 9548
rect 17104 9514 17110 9548
rect 17064 9476 17110 9514
rect 17064 9442 17070 9476
rect 17104 9442 17110 9476
rect 17064 9404 17110 9442
rect 17064 9370 17070 9404
rect 17104 9370 17110 9404
rect 17064 9332 17110 9370
rect 17064 9298 17070 9332
rect 17104 9298 17110 9332
rect 17064 9260 17110 9298
rect 17064 9226 17070 9260
rect 17104 9226 17110 9260
rect 17064 9188 17110 9226
rect 17064 9154 17070 9188
rect 17104 9154 17110 9188
rect 17064 9116 17110 9154
rect 17064 9082 17070 9116
rect 17104 9082 17110 9116
rect 17064 9044 17110 9082
rect 17064 9010 17070 9044
rect 17104 9010 17110 9044
rect 17064 8972 17110 9010
rect 17064 8938 17070 8972
rect 17104 8938 17110 8972
rect 17064 8900 17110 8938
rect 17064 8866 17070 8900
rect 17104 8866 17110 8900
rect 17064 8828 17110 8866
rect 17064 8794 17070 8828
rect 17104 8794 17110 8828
rect 17064 8756 17110 8794
rect 17064 8722 17070 8756
rect 17104 8722 17110 8756
rect 17064 8700 17110 8722
rect 17472 11034 17518 11072
rect 17472 11000 17478 11034
rect 17512 11000 17518 11034
rect 17472 10962 17518 11000
rect 17472 10928 17478 10962
rect 17512 10928 17518 10962
rect 17472 10890 17518 10928
rect 18466 11144 18536 11174
rect 18570 11174 18576 11178
rect 19588 11219 19634 11221
rect 19786 11219 20250 11222
rect 19588 11178 20250 11219
rect 18570 11144 18646 11174
rect 18466 11129 18646 11144
rect 18466 10949 18498 11129
rect 18614 10949 18646 11129
rect 18466 10928 18536 10949
rect 18570 10928 18646 10949
rect 18466 10904 18646 10928
rect 19588 11144 19594 11178
rect 19628 11144 20250 11178
rect 19588 11106 20250 11144
rect 19588 11072 19594 11106
rect 19628 11072 20250 11106
rect 19588 11034 20250 11072
rect 19588 11000 19594 11034
rect 19628 11000 20250 11034
rect 19588 10962 20250 11000
rect 19588 10928 19594 10962
rect 19628 10928 20250 10962
rect 17472 10856 17478 10890
rect 17512 10856 17518 10890
rect 17472 10818 17518 10856
rect 17472 10784 17478 10818
rect 17512 10784 17518 10818
rect 17472 10746 17518 10784
rect 17472 10712 17478 10746
rect 17512 10712 17518 10746
rect 17472 10674 17518 10712
rect 17472 10640 17478 10674
rect 17512 10640 17518 10674
rect 17472 10602 17518 10640
rect 17472 10568 17478 10602
rect 17512 10568 17518 10602
rect 17472 10530 17518 10568
rect 17472 10496 17478 10530
rect 17512 10496 17518 10530
rect 17472 10458 17518 10496
rect 17472 10424 17478 10458
rect 17512 10424 17518 10458
rect 17472 10386 17518 10424
rect 17472 10352 17478 10386
rect 17512 10352 17518 10386
rect 17472 10314 17518 10352
rect 17472 10280 17478 10314
rect 17512 10280 17518 10314
rect 17472 10242 17518 10280
rect 17472 10208 17478 10242
rect 17512 10208 17518 10242
rect 17472 10170 17518 10208
rect 17472 10136 17478 10170
rect 17512 10136 17518 10170
rect 17472 10098 17518 10136
rect 17472 10064 17478 10098
rect 17512 10064 17518 10098
rect 17472 10026 17518 10064
rect 17472 9992 17478 10026
rect 17512 9992 17518 10026
rect 17472 9954 17518 9992
rect 17472 9920 17478 9954
rect 17512 9920 17518 9954
rect 17472 9882 17518 9920
rect 17472 9848 17478 9882
rect 17512 9848 17518 9882
rect 17472 9810 17518 9848
rect 17472 9776 17478 9810
rect 17512 9776 17518 9810
rect 17472 9738 17518 9776
rect 17472 9704 17478 9738
rect 17512 9704 17518 9738
rect 17472 9666 17518 9704
rect 17472 9632 17478 9666
rect 17512 9632 17518 9666
rect 17472 9594 17518 9632
rect 17472 9560 17478 9594
rect 17512 9560 17518 9594
rect 17472 9522 17518 9560
rect 17472 9488 17478 9522
rect 17512 9488 17518 9522
rect 17472 9450 17518 9488
rect 17472 9416 17478 9450
rect 17512 9416 17518 9450
rect 17472 9378 17518 9416
rect 17472 9344 17478 9378
rect 17512 9344 17518 9378
rect 17472 9306 17518 9344
rect 17472 9272 17478 9306
rect 17512 9272 17518 9306
rect 17472 9234 17518 9272
rect 17472 9200 17478 9234
rect 17512 9200 17518 9234
rect 17472 9162 17518 9200
rect 17472 9128 17478 9162
rect 17512 9128 17518 9162
rect 17472 9090 17518 9128
rect 17472 9056 17478 9090
rect 17512 9056 17518 9090
rect 17472 9018 17518 9056
rect 17472 8984 17478 9018
rect 17512 8984 17518 9018
rect 17472 8946 17518 8984
rect 17472 8912 17478 8946
rect 17512 8912 17518 8946
rect 17472 8874 17518 8912
rect 17472 8840 17478 8874
rect 17512 8840 17518 8874
rect 17472 8802 17518 8840
rect 17472 8768 17478 8802
rect 17512 8768 17518 8802
rect 17472 8730 17518 8768
rect 16006 8650 16012 8684
rect 16046 8650 16052 8684
rect 16006 8612 16052 8650
rect 16006 8578 16012 8612
rect 16046 8578 16052 8612
rect 16006 8540 16052 8578
rect 16006 8506 16012 8540
rect 16046 8506 16052 8540
rect 16006 8468 16052 8506
rect 16006 8434 16012 8468
rect 16046 8434 16052 8468
rect 16006 8396 16052 8434
rect 16006 8362 16012 8396
rect 16046 8362 16052 8396
rect 16006 8324 16052 8362
rect 16006 8290 16012 8324
rect 16046 8290 16052 8324
rect 14948 8247 14994 8270
rect 16006 8247 16052 8290
rect 16912 8684 17122 8700
rect 16912 8676 17070 8684
rect 16912 8304 16959 8676
rect 17104 8650 17122 8684
rect 17472 8696 17478 8730
rect 17512 8696 17518 8730
rect 17472 8674 17518 8696
rect 18530 10890 18576 10904
rect 18530 10856 18536 10890
rect 18570 10856 18576 10890
rect 18530 10818 18576 10856
rect 18530 10784 18536 10818
rect 18570 10784 18576 10818
rect 18530 10746 18576 10784
rect 18530 10712 18536 10746
rect 18570 10712 18576 10746
rect 18530 10674 18576 10712
rect 18530 10640 18536 10674
rect 18570 10640 18576 10674
rect 18530 10602 18576 10640
rect 18530 10568 18536 10602
rect 18570 10568 18576 10602
rect 18530 10530 18576 10568
rect 18530 10496 18536 10530
rect 18570 10496 18576 10530
rect 18530 10458 18576 10496
rect 18530 10424 18536 10458
rect 18570 10424 18576 10458
rect 18530 10386 18576 10424
rect 18530 10352 18536 10386
rect 18570 10352 18576 10386
rect 18530 10314 18576 10352
rect 18530 10280 18536 10314
rect 18570 10280 18576 10314
rect 18530 10242 18576 10280
rect 18530 10208 18536 10242
rect 18570 10208 18576 10242
rect 18530 10170 18576 10208
rect 18530 10136 18536 10170
rect 18570 10136 18576 10170
rect 18530 10098 18576 10136
rect 18530 10064 18536 10098
rect 18570 10064 18576 10098
rect 18530 10026 18576 10064
rect 18530 9992 18536 10026
rect 18570 9992 18576 10026
rect 18530 9954 18576 9992
rect 18530 9920 18536 9954
rect 18570 9920 18576 9954
rect 18530 9882 18576 9920
rect 18530 9848 18536 9882
rect 18570 9848 18576 9882
rect 18530 9810 18576 9848
rect 18530 9776 18536 9810
rect 18570 9776 18576 9810
rect 18530 9738 18576 9776
rect 18530 9704 18536 9738
rect 18570 9704 18576 9738
rect 18530 9666 18576 9704
rect 18530 9632 18536 9666
rect 18570 9632 18576 9666
rect 18530 9594 18576 9632
rect 18530 9560 18536 9594
rect 18570 9560 18576 9594
rect 18530 9522 18576 9560
rect 18530 9488 18536 9522
rect 18570 9488 18576 9522
rect 18530 9450 18576 9488
rect 18530 9416 18536 9450
rect 18570 9416 18576 9450
rect 18530 9378 18576 9416
rect 18530 9344 18536 9378
rect 18570 9344 18576 9378
rect 18530 9306 18576 9344
rect 18530 9272 18536 9306
rect 18570 9272 18576 9306
rect 18530 9234 18576 9272
rect 18530 9200 18536 9234
rect 18570 9200 18576 9234
rect 18530 9162 18576 9200
rect 18530 9128 18536 9162
rect 18570 9128 18576 9162
rect 18530 9090 18576 9128
rect 18530 9056 18536 9090
rect 18570 9056 18576 9090
rect 18530 9018 18576 9056
rect 18530 8984 18536 9018
rect 18570 8984 18576 9018
rect 18530 8946 18576 8984
rect 18530 8912 18536 8946
rect 18570 8912 18576 8946
rect 18530 8874 18576 8912
rect 18530 8840 18536 8874
rect 18570 8840 18576 8874
rect 18530 8802 18576 8840
rect 18530 8768 18536 8802
rect 18570 8768 18576 8802
rect 18530 8730 18576 8768
rect 18530 8696 18536 8730
rect 18570 8696 18576 8730
rect 17075 8612 17122 8650
rect 17104 8578 17122 8612
rect 17075 8560 17122 8578
rect 17446 8658 17616 8674
rect 17446 8638 17478 8658
rect 17512 8638 17616 8658
rect 17075 8540 17382 8560
rect 17104 8506 17382 8540
rect 17075 8468 17382 8506
rect 17104 8434 17382 8468
rect 17075 8420 17382 8434
rect 17075 8396 17122 8420
rect 17104 8362 17122 8396
rect 17075 8324 17122 8362
rect 16912 8290 17070 8304
rect 17104 8290 17122 8324
rect 16912 8270 17122 8290
rect 17064 8247 17110 8270
rect 16902 8206 17058 8208
rect 15004 8200 15996 8206
rect 16062 8200 17058 8206
rect 15004 8166 15051 8200
rect 15085 8166 15123 8200
rect 15157 8166 15195 8200
rect 15229 8166 15267 8200
rect 15301 8166 15339 8200
rect 15373 8166 15411 8200
rect 15445 8166 15483 8200
rect 15517 8166 15555 8200
rect 15589 8166 15627 8200
rect 15661 8166 15699 8200
rect 15733 8166 15771 8200
rect 15805 8166 15843 8200
rect 15877 8166 15915 8200
rect 15949 8166 16109 8200
rect 16143 8166 16181 8200
rect 16215 8166 16253 8200
rect 16287 8166 16325 8200
rect 16359 8166 16397 8200
rect 16431 8166 16469 8200
rect 16503 8166 16541 8200
rect 16575 8166 16613 8200
rect 16647 8166 16685 8200
rect 16719 8166 16757 8200
rect 16791 8166 16829 8200
rect 16863 8166 16901 8200
rect 16935 8187 16973 8200
rect 17007 8187 17058 8200
rect 15004 8160 16922 8166
rect 15822 8130 16252 8160
rect 16902 8007 16922 8160
rect 17038 8007 17058 8187
rect 16412 7980 16652 7990
rect 16902 7982 17058 8007
rect 14462 7760 16662 7980
rect 16832 7877 17082 7930
rect 13111 7716 13142 7750
rect 13176 7716 13242 7750
rect 13276 7716 13342 7750
rect 13376 7716 13442 7750
rect 13476 7716 13542 7750
rect 13576 7716 13642 7750
rect 13676 7716 13721 7750
rect -7862 7626 -3668 7700
rect -7862 7610 -7538 7626
rect -7862 7576 -7687 7610
rect -7653 7576 -7615 7610
rect -7581 7576 -7538 7610
rect -7862 7570 -7538 7576
rect -7472 7610 -7280 7626
rect -7472 7576 -7429 7610
rect -7395 7576 -7357 7610
rect -7323 7576 -7280 7610
rect -7472 7570 -7280 7576
rect -7214 7610 -7022 7626
rect -7214 7576 -7171 7610
rect -7137 7576 -7099 7610
rect -7065 7576 -7022 7610
rect -7214 7570 -7022 7576
rect -6956 7616 -4442 7626
rect -6956 7610 -6764 7616
rect -6956 7576 -6913 7610
rect -6879 7576 -6841 7610
rect -6807 7576 -6764 7610
rect -6956 7570 -6764 7576
rect -6698 7610 -6506 7616
rect -6698 7576 -6655 7610
rect -6621 7576 -6583 7610
rect -6549 7576 -6506 7610
rect -6698 7570 -6506 7576
rect -6440 7610 -6248 7616
rect -6440 7576 -6397 7610
rect -6363 7576 -6325 7610
rect -6291 7576 -6248 7610
rect -6440 7570 -6248 7576
rect -6182 7610 -5990 7616
rect -6182 7576 -6139 7610
rect -6105 7576 -6067 7610
rect -6033 7576 -5990 7610
rect -6182 7570 -5990 7576
rect -5924 7610 -5732 7616
rect -5924 7576 -5881 7610
rect -5847 7576 -5809 7610
rect -5775 7576 -5732 7610
rect -5924 7570 -5732 7576
rect -5666 7610 -5474 7616
rect -5666 7576 -5623 7610
rect -5589 7576 -5551 7610
rect -5517 7576 -5474 7610
rect -5666 7570 -5474 7576
rect -5408 7610 -5216 7616
rect -5408 7576 -5365 7610
rect -5331 7576 -5293 7610
rect -5259 7576 -5216 7610
rect -5408 7570 -5216 7576
rect -5150 7610 -4958 7616
rect -5150 7576 -5107 7610
rect -5073 7576 -5035 7610
rect -5001 7576 -4958 7610
rect -5150 7570 -4958 7576
rect -4892 7610 -4700 7616
rect -4892 7576 -4849 7610
rect -4815 7576 -4777 7610
rect -4743 7576 -4700 7610
rect -4892 7570 -4700 7576
rect -4634 7610 -4442 7616
rect -4634 7576 -4591 7610
rect -4557 7576 -4519 7610
rect -4485 7576 -4442 7610
rect -4634 7570 -4442 7576
rect -4376 7610 -4184 7626
rect -4376 7576 -4333 7610
rect -4299 7576 -4261 7610
rect -4227 7576 -4184 7610
rect -4376 7570 -4184 7576
rect -4118 7610 -3926 7626
rect -4118 7576 -4075 7610
rect -4041 7576 -4003 7610
rect -3969 7576 -3926 7610
rect -4118 7570 -3926 7576
rect -3860 7610 -3668 7626
rect -3860 7576 -3817 7610
rect -3783 7576 -3745 7610
rect -3711 7576 -3668 7610
rect -3860 7570 -3668 7576
rect 13111 7650 13721 7716
rect 13111 7616 13142 7650
rect 13176 7616 13242 7650
rect 13276 7616 13342 7650
rect 13376 7616 13442 7650
rect 13476 7616 13542 7650
rect 13576 7616 13642 7650
rect 13676 7616 13721 7650
rect -7862 7491 -7740 7570
rect 13111 7550 13721 7616
rect -7862 7457 -7780 7491
rect -7746 7457 -7740 7491
rect -7862 7419 -7740 7457
rect -7862 7385 -7780 7419
rect -7746 7385 -7740 7419
rect -7862 7363 -7740 7385
rect -7786 7347 -7740 7363
rect -7786 7313 -7780 7347
rect -7746 7313 -7740 7347
rect -7786 7275 -7740 7313
rect -7786 7241 -7780 7275
rect -7746 7241 -7740 7275
rect -7786 7203 -7740 7241
rect -7786 7169 -7780 7203
rect -7746 7169 -7740 7203
rect -7786 7131 -7740 7169
rect -7786 7097 -7780 7131
rect -7746 7097 -7740 7131
rect -7786 7059 -7740 7097
rect -7786 7025 -7780 7059
rect -7746 7025 -7740 7059
rect -7786 6987 -7740 7025
rect -7786 6953 -7780 6987
rect -7746 6953 -7740 6987
rect -7786 6915 -7740 6953
rect -7786 6881 -7780 6915
rect -7746 6881 -7740 6915
rect -7786 6843 -7740 6881
rect -7786 6809 -7780 6843
rect -7746 6809 -7740 6843
rect -7786 6771 -7740 6809
rect -7786 6737 -7780 6771
rect -7746 6737 -7740 6771
rect -7786 6699 -7740 6737
rect -7786 6665 -7780 6699
rect -7746 6665 -7740 6699
rect -7786 6627 -7740 6665
rect -7786 6593 -7780 6627
rect -7746 6593 -7740 6627
rect -7786 6555 -7740 6593
rect -7786 6521 -7780 6555
rect -7746 6521 -7740 6555
rect -7786 6483 -7740 6521
rect -7786 6449 -7780 6483
rect -7746 6449 -7740 6483
rect -7786 6411 -7740 6449
rect -7786 6377 -7780 6411
rect -7746 6377 -7740 6411
rect -7786 6339 -7740 6377
rect -7786 6305 -7780 6339
rect -7746 6305 -7740 6339
rect -7786 6267 -7740 6305
rect -7786 6233 -7780 6267
rect -7746 6233 -7740 6267
rect -7786 6195 -7740 6233
rect -7786 6161 -7780 6195
rect -7746 6161 -7740 6195
rect -7786 6123 -7740 6161
rect -7786 6089 -7780 6123
rect -7746 6089 -7740 6123
rect -7786 6051 -7740 6089
rect -7786 6017 -7780 6051
rect -7746 6017 -7740 6051
rect -7786 5979 -7740 6017
rect -7786 5945 -7780 5979
rect -7746 5945 -7740 5979
rect -7786 5907 -7740 5945
rect -7997 5886 -7909 5901
rect -7997 5834 -7980 5886
rect -7928 5834 -7909 5886
rect -7997 5822 -7909 5834
rect -7997 5770 -7980 5822
rect -7928 5770 -7909 5822
rect -7997 5758 -7909 5770
rect -7997 5706 -7980 5758
rect -7928 5706 -7909 5758
rect -7997 5693 -7909 5706
rect -7786 5873 -7780 5907
rect -7746 5873 -7740 5907
rect -7528 7491 -7482 7538
rect -7528 7457 -7522 7491
rect -7488 7457 -7482 7491
rect -7528 7419 -7482 7457
rect -7528 7385 -7522 7419
rect -7488 7385 -7482 7419
rect -7528 7347 -7482 7385
rect -7528 7313 -7522 7347
rect -7488 7313 -7482 7347
rect -7528 7275 -7482 7313
rect -7528 7241 -7522 7275
rect -7488 7241 -7482 7275
rect -7528 7203 -7482 7241
rect -7528 7169 -7522 7203
rect -7488 7169 -7482 7203
rect -7528 7131 -7482 7169
rect -7528 7097 -7522 7131
rect -7488 7097 -7482 7131
rect -7528 7059 -7482 7097
rect -7528 7025 -7522 7059
rect -7488 7025 -7482 7059
rect -7528 6987 -7482 7025
rect -7528 6953 -7522 6987
rect -7488 6953 -7482 6987
rect -7528 6915 -7482 6953
rect -7528 6881 -7522 6915
rect -7488 6881 -7482 6915
rect -7528 6843 -7482 6881
rect -7528 6809 -7522 6843
rect -7488 6809 -7482 6843
rect -7270 7491 -7224 7538
rect -7270 7457 -7264 7491
rect -7230 7457 -7224 7491
rect -7270 7419 -7224 7457
rect -7270 7385 -7264 7419
rect -7230 7385 -7224 7419
rect -7270 7347 -7224 7385
rect -7270 7313 -7264 7347
rect -7230 7313 -7224 7347
rect -7270 7275 -7224 7313
rect -7270 7241 -7264 7275
rect -7230 7241 -7224 7275
rect -7270 7203 -7224 7241
rect -7270 7169 -7264 7203
rect -7230 7169 -7224 7203
rect -7270 7131 -7224 7169
rect -7270 7097 -7264 7131
rect -7230 7097 -7224 7131
rect -7270 7059 -7224 7097
rect -7270 7025 -7264 7059
rect -7230 7025 -7224 7059
rect -7270 6987 -7224 7025
rect -7270 6953 -7264 6987
rect -7230 6953 -7224 6987
rect -7270 6915 -7224 6953
rect -7270 6881 -7264 6915
rect -7230 6881 -7224 6915
rect -7270 6843 -7224 6881
rect -7270 6811 -7264 6843
rect -7528 6771 -7482 6809
rect -7528 6737 -7522 6771
rect -7488 6737 -7482 6771
rect -7528 6699 -7482 6737
rect -7528 6665 -7522 6699
rect -7488 6665 -7482 6699
rect -7528 6627 -7482 6665
rect -7528 6593 -7522 6627
rect -7488 6593 -7482 6627
rect -7290 6809 -7264 6811
rect -7230 6811 -7224 6843
rect -7012 7491 -6966 7538
rect -7012 7457 -7006 7491
rect -6972 7457 -6966 7491
rect -7012 7419 -6966 7457
rect -7012 7385 -7006 7419
rect -6972 7385 -6966 7419
rect -7012 7347 -6966 7385
rect -7012 7313 -7006 7347
rect -6972 7313 -6966 7347
rect -7012 7275 -6966 7313
rect -7012 7241 -7006 7275
rect -6972 7241 -6966 7275
rect -7012 7203 -6966 7241
rect -7012 7169 -7006 7203
rect -6972 7169 -6966 7203
rect -7012 7131 -6966 7169
rect -7012 7097 -7006 7131
rect -6972 7097 -6966 7131
rect -7012 7059 -6966 7097
rect -7012 7025 -7006 7059
rect -6972 7025 -6966 7059
rect -7012 6987 -6966 7025
rect -7012 6953 -7006 6987
rect -6972 6953 -6966 6987
rect -7012 6915 -6966 6953
rect -7012 6881 -7006 6915
rect -6972 6881 -6966 6915
rect -7012 6843 -6966 6881
rect -7230 6809 -7204 6811
rect -7290 6771 -7204 6809
rect -7290 6765 -7264 6771
rect -7230 6765 -7204 6771
rect -7290 6713 -7273 6765
rect -7221 6713 -7204 6765
rect -7290 6701 -7204 6713
rect -7290 6649 -7273 6701
rect -7221 6649 -7204 6701
rect -7290 6627 -7204 6649
rect -7290 6606 -7264 6627
rect -7528 6555 -7482 6593
rect -7528 6521 -7522 6555
rect -7488 6521 -7482 6555
rect -7528 6483 -7482 6521
rect -7528 6449 -7522 6483
rect -7488 6449 -7482 6483
rect -7528 6411 -7482 6449
rect -7528 6377 -7522 6411
rect -7488 6377 -7482 6411
rect -7528 6339 -7482 6377
rect -7528 6305 -7522 6339
rect -7488 6305 -7482 6339
rect -7528 6267 -7482 6305
rect -7528 6233 -7522 6267
rect -7488 6233 -7482 6267
rect -7528 6195 -7482 6233
rect -7528 6161 -7522 6195
rect -7488 6161 -7482 6195
rect -7528 6123 -7482 6161
rect -7528 6089 -7522 6123
rect -7488 6089 -7482 6123
rect -7528 6051 -7482 6089
rect -7528 6017 -7522 6051
rect -7488 6017 -7482 6051
rect -7528 5979 -7482 6017
rect -7528 5945 -7522 5979
rect -7488 5945 -7482 5979
rect -7528 5907 -7482 5945
rect -7528 5901 -7522 5907
rect -7786 5835 -7740 5873
rect -7786 5801 -7780 5835
rect -7746 5801 -7740 5835
rect -7786 5763 -7740 5801
rect -7786 5729 -7780 5763
rect -7746 5729 -7740 5763
rect -7786 5691 -7740 5729
rect -7536 5888 -7522 5901
rect -7488 5901 -7482 5907
rect -7270 6593 -7264 6606
rect -7230 6606 -7204 6627
rect -7012 6809 -7006 6843
rect -6972 6809 -6966 6843
rect -7012 6771 -6966 6809
rect -7012 6737 -7006 6771
rect -6972 6737 -6966 6771
rect -7012 6699 -6966 6737
rect -7012 6665 -7006 6699
rect -6972 6665 -6966 6699
rect -7012 6627 -6966 6665
rect -7230 6593 -7224 6606
rect -7270 6555 -7224 6593
rect -7270 6521 -7264 6555
rect -7230 6521 -7224 6555
rect -7270 6483 -7224 6521
rect -7270 6449 -7264 6483
rect -7230 6449 -7224 6483
rect -7270 6411 -7224 6449
rect -7270 6377 -7264 6411
rect -7230 6377 -7224 6411
rect -7270 6339 -7224 6377
rect -7270 6305 -7264 6339
rect -7230 6305 -7224 6339
rect -7270 6267 -7224 6305
rect -7270 6233 -7264 6267
rect -7230 6233 -7224 6267
rect -7270 6195 -7224 6233
rect -7270 6161 -7264 6195
rect -7230 6161 -7224 6195
rect -7270 6123 -7224 6161
rect -7270 6089 -7264 6123
rect -7230 6089 -7224 6123
rect -7270 6051 -7224 6089
rect -7270 6017 -7264 6051
rect -7230 6017 -7224 6051
rect -7270 5979 -7224 6017
rect -7270 5945 -7264 5979
rect -7230 5945 -7224 5979
rect -7270 5907 -7224 5945
rect -7488 5888 -7474 5901
rect -7536 5836 -7532 5888
rect -7480 5836 -7474 5888
rect -7536 5835 -7474 5836
rect -7536 5824 -7522 5835
rect -7488 5824 -7474 5835
rect -7536 5772 -7532 5824
rect -7480 5772 -7474 5824
rect -7536 5763 -7474 5772
rect -7536 5760 -7522 5763
rect -7488 5760 -7474 5763
rect -7536 5708 -7532 5760
rect -7480 5708 -7474 5760
rect -7536 5693 -7474 5708
rect -7270 5873 -7264 5907
rect -7230 5873 -7224 5907
rect -7012 6593 -7006 6627
rect -6972 6593 -6966 6627
rect -7012 6555 -6966 6593
rect -7012 6521 -7006 6555
rect -6972 6521 -6966 6555
rect -7012 6483 -6966 6521
rect -7012 6449 -7006 6483
rect -6972 6449 -6966 6483
rect -7012 6411 -6966 6449
rect -7012 6377 -7006 6411
rect -6972 6377 -6966 6411
rect -7012 6339 -6966 6377
rect -6754 7491 -6708 7538
rect -6754 7457 -6748 7491
rect -6714 7457 -6708 7491
rect -6754 7419 -6708 7457
rect -6754 7385 -6748 7419
rect -6714 7385 -6708 7419
rect -6754 7347 -6708 7385
rect -6754 7313 -6748 7347
rect -6714 7313 -6708 7347
rect -6754 7275 -6708 7313
rect -6754 7241 -6748 7275
rect -6714 7241 -6708 7275
rect -6754 7203 -6708 7241
rect -6754 7169 -6748 7203
rect -6714 7169 -6708 7203
rect -6754 7131 -6708 7169
rect -6754 7097 -6748 7131
rect -6714 7097 -6708 7131
rect -6754 7059 -6708 7097
rect -6754 7025 -6748 7059
rect -6714 7025 -6708 7059
rect -6754 6987 -6708 7025
rect -6754 6953 -6748 6987
rect -6714 6953 -6708 6987
rect -6754 6915 -6708 6953
rect -6754 6881 -6748 6915
rect -6714 6881 -6708 6915
rect -6754 6843 -6708 6881
rect -6754 6809 -6748 6843
rect -6714 6809 -6708 6843
rect -6754 6771 -6708 6809
rect -6754 6737 -6748 6771
rect -6714 6737 -6708 6771
rect -6754 6699 -6708 6737
rect -6754 6665 -6748 6699
rect -6714 6665 -6708 6699
rect -6754 6627 -6708 6665
rect -6754 6593 -6748 6627
rect -6714 6593 -6708 6627
rect -6754 6555 -6708 6593
rect -6754 6521 -6748 6555
rect -6714 6521 -6708 6555
rect -6754 6483 -6708 6521
rect -6754 6449 -6748 6483
rect -6714 6449 -6708 6483
rect -6754 6411 -6708 6449
rect -6754 6377 -6748 6411
rect -6714 6377 -6708 6411
rect -6754 6375 -6708 6377
rect -6496 7491 -6450 7538
rect -6496 7457 -6490 7491
rect -6456 7457 -6450 7491
rect -6496 7419 -6450 7457
rect -6496 7385 -6490 7419
rect -6456 7385 -6450 7419
rect -6496 7347 -6450 7385
rect -6496 7313 -6490 7347
rect -6456 7313 -6450 7347
rect -6496 7275 -6450 7313
rect -6496 7241 -6490 7275
rect -6456 7241 -6450 7275
rect -6496 7203 -6450 7241
rect -6496 7169 -6490 7203
rect -6456 7169 -6450 7203
rect -6496 7131 -6450 7169
rect -6496 7097 -6490 7131
rect -6456 7097 -6450 7131
rect -6496 7059 -6450 7097
rect -6496 7025 -6490 7059
rect -6456 7025 -6450 7059
rect -6496 6987 -6450 7025
rect -6496 6953 -6490 6987
rect -6456 6953 -6450 6987
rect -6496 6915 -6450 6953
rect -6496 6881 -6490 6915
rect -6456 6881 -6450 6915
rect -6496 6843 -6450 6881
rect -6496 6809 -6490 6843
rect -6456 6809 -6450 6843
rect -6496 6771 -6450 6809
rect -6496 6737 -6490 6771
rect -6456 6737 -6450 6771
rect -6496 6699 -6450 6737
rect -6496 6665 -6490 6699
rect -6456 6665 -6450 6699
rect -6496 6627 -6450 6665
rect -6496 6593 -6490 6627
rect -6456 6593 -6450 6627
rect -6496 6555 -6450 6593
rect -6496 6521 -6490 6555
rect -6456 6521 -6450 6555
rect -6496 6483 -6450 6521
rect -6496 6449 -6490 6483
rect -6456 6449 -6450 6483
rect -6496 6411 -6450 6449
rect -6496 6377 -6490 6411
rect -6456 6377 -6450 6411
rect -7012 6305 -7006 6339
rect -6972 6305 -6966 6339
rect -7012 6267 -6966 6305
rect -7012 6233 -7006 6267
rect -6972 6233 -6966 6267
rect -7012 6195 -6966 6233
rect -7012 6161 -7006 6195
rect -6972 6161 -6966 6195
rect -6790 6362 -6677 6375
rect -6790 6310 -6757 6362
rect -6705 6310 -6677 6362
rect -6790 6305 -6748 6310
rect -6714 6305 -6677 6310
rect -6790 6298 -6677 6305
rect -6790 6246 -6757 6298
rect -6705 6246 -6677 6298
rect -6790 6234 -6748 6246
rect -6714 6234 -6677 6246
rect -6790 6182 -6757 6234
rect -6705 6182 -6677 6234
rect -6790 6168 -6748 6182
rect -7012 6123 -6966 6161
rect -7012 6089 -7006 6123
rect -6972 6089 -6966 6123
rect -7012 6051 -6966 6089
rect -7012 6017 -7006 6051
rect -6972 6017 -6966 6051
rect -7012 5979 -6966 6017
rect -7012 5945 -7006 5979
rect -6972 5945 -6966 5979
rect -7012 5907 -6966 5945
rect -7012 5902 -7006 5907
rect -7270 5835 -7224 5873
rect -7270 5801 -7264 5835
rect -7230 5801 -7224 5835
rect -7270 5763 -7224 5801
rect -7270 5729 -7264 5763
rect -7230 5729 -7224 5763
rect -7786 5657 -7780 5691
rect -7746 5657 -7740 5691
rect -7786 5619 -7740 5657
rect -7786 5585 -7780 5619
rect -7746 5585 -7740 5619
rect -7786 5506 -7740 5585
rect -7528 5691 -7482 5693
rect -7528 5657 -7522 5691
rect -7488 5657 -7482 5691
rect -7528 5619 -7482 5657
rect -7528 5585 -7522 5619
rect -7488 5585 -7482 5619
rect -7528 5538 -7482 5585
rect -7270 5691 -7224 5729
rect -7025 5887 -7006 5902
rect -6972 5902 -6966 5907
rect -6754 6161 -6748 6168
rect -6714 6168 -6677 6182
rect -6496 6339 -6450 6377
rect -6238 7491 -6192 7538
rect -6238 7457 -6232 7491
rect -6198 7457 -6192 7491
rect -6238 7419 -6192 7457
rect -6238 7385 -6232 7419
rect -6198 7385 -6192 7419
rect -6238 7347 -6192 7385
rect -6238 7313 -6232 7347
rect -6198 7313 -6192 7347
rect -6238 7275 -6192 7313
rect -6238 7241 -6232 7275
rect -6198 7241 -6192 7275
rect -6238 7203 -6192 7241
rect -6238 7169 -6232 7203
rect -6198 7169 -6192 7203
rect -6238 7131 -6192 7169
rect -6238 7097 -6232 7131
rect -6198 7097 -6192 7131
rect -6238 7059 -6192 7097
rect -6238 7025 -6232 7059
rect -6198 7025 -6192 7059
rect -6238 6987 -6192 7025
rect -6238 6953 -6232 6987
rect -6198 6953 -6192 6987
rect -6238 6915 -6192 6953
rect -6238 6881 -6232 6915
rect -6198 6881 -6192 6915
rect -6238 6843 -6192 6881
rect -6238 6809 -6232 6843
rect -6198 6809 -6192 6843
rect -6238 6771 -6192 6809
rect -6238 6737 -6232 6771
rect -6198 6737 -6192 6771
rect -6238 6699 -6192 6737
rect -6238 6665 -6232 6699
rect -6198 6665 -6192 6699
rect -6238 6627 -6192 6665
rect -6238 6593 -6232 6627
rect -6198 6593 -6192 6627
rect -6238 6555 -6192 6593
rect -6238 6521 -6232 6555
rect -6198 6521 -6192 6555
rect -6238 6483 -6192 6521
rect -6238 6449 -6232 6483
rect -6198 6449 -6192 6483
rect -6238 6411 -6192 6449
rect -6238 6377 -6232 6411
rect -6198 6377 -6192 6411
rect -6238 6375 -6192 6377
rect -5980 7491 -5934 7538
rect -5980 7457 -5974 7491
rect -5940 7457 -5934 7491
rect -5980 7419 -5934 7457
rect -5980 7385 -5974 7419
rect -5940 7385 -5934 7419
rect -5980 7347 -5934 7385
rect -5980 7313 -5974 7347
rect -5940 7313 -5934 7347
rect -5980 7275 -5934 7313
rect -5980 7241 -5974 7275
rect -5940 7241 -5934 7275
rect -5980 7203 -5934 7241
rect -5980 7169 -5974 7203
rect -5940 7169 -5934 7203
rect -5980 7131 -5934 7169
rect -5980 7097 -5974 7131
rect -5940 7097 -5934 7131
rect -5980 7059 -5934 7097
rect -5980 7025 -5974 7059
rect -5940 7025 -5934 7059
rect -5980 6987 -5934 7025
rect -5980 6953 -5974 6987
rect -5940 6953 -5934 6987
rect -5980 6915 -5934 6953
rect -5980 6881 -5974 6915
rect -5940 6881 -5934 6915
rect -5980 6843 -5934 6881
rect -5980 6809 -5974 6843
rect -5940 6809 -5934 6843
rect -5980 6771 -5934 6809
rect -5980 6737 -5974 6771
rect -5940 6737 -5934 6771
rect -5980 6699 -5934 6737
rect -5980 6665 -5974 6699
rect -5940 6665 -5934 6699
rect -5980 6627 -5934 6665
rect -5980 6593 -5974 6627
rect -5940 6593 -5934 6627
rect -5980 6555 -5934 6593
rect -5980 6521 -5974 6555
rect -5940 6521 -5934 6555
rect -5980 6483 -5934 6521
rect -5980 6449 -5974 6483
rect -5940 6449 -5934 6483
rect -5980 6411 -5934 6449
rect -5980 6377 -5974 6411
rect -5940 6377 -5934 6411
rect -6496 6305 -6490 6339
rect -6456 6305 -6450 6339
rect -6496 6267 -6450 6305
rect -6496 6233 -6490 6267
rect -6456 6233 -6450 6267
rect -6496 6195 -6450 6233
rect -6714 6161 -6708 6168
rect -6754 6123 -6708 6161
rect -6754 6089 -6748 6123
rect -6714 6089 -6708 6123
rect -6754 6051 -6708 6089
rect -6754 6017 -6748 6051
rect -6714 6017 -6708 6051
rect -6754 5979 -6708 6017
rect -6754 5945 -6748 5979
rect -6714 5945 -6708 5979
rect -6754 5907 -6708 5945
rect -6972 5887 -6954 5902
rect -7025 5835 -7015 5887
rect -6963 5835 -6954 5887
rect -7025 5823 -7006 5835
rect -6972 5823 -6954 5835
rect -7025 5771 -7015 5823
rect -6963 5771 -6954 5823
rect -7025 5763 -6954 5771
rect -7025 5759 -7006 5763
rect -6972 5759 -6954 5763
rect -7025 5707 -7015 5759
rect -6963 5707 -6954 5759
rect -7025 5694 -6954 5707
rect -6754 5873 -6748 5907
rect -6714 5873 -6708 5907
rect -6496 6161 -6490 6195
rect -6456 6161 -6450 6195
rect -6260 6360 -6171 6375
rect -6260 6308 -6241 6360
rect -6189 6308 -6171 6360
rect -6260 6305 -6232 6308
rect -6198 6305 -6171 6308
rect -6260 6296 -6171 6305
rect -6260 6244 -6241 6296
rect -6189 6244 -6171 6296
rect -6260 6233 -6232 6244
rect -6198 6233 -6171 6244
rect -6260 6232 -6171 6233
rect -6260 6180 -6241 6232
rect -6189 6180 -6171 6232
rect -6260 6168 -6232 6180
rect -6496 6123 -6450 6161
rect -6496 6089 -6490 6123
rect -6456 6089 -6450 6123
rect -6496 6051 -6450 6089
rect -6496 6017 -6490 6051
rect -6456 6017 -6450 6051
rect -6496 5979 -6450 6017
rect -6496 5945 -6490 5979
rect -6456 5945 -6450 5979
rect -6496 5907 -6450 5945
rect -6496 5901 -6490 5907
rect -6754 5835 -6708 5873
rect -6754 5801 -6748 5835
rect -6714 5801 -6708 5835
rect -6754 5763 -6708 5801
rect -6754 5729 -6748 5763
rect -6714 5729 -6708 5763
rect -7270 5657 -7264 5691
rect -7230 5657 -7224 5691
rect -7270 5619 -7224 5657
rect -7270 5585 -7264 5619
rect -7230 5585 -7224 5619
rect -7270 5538 -7224 5585
rect -7012 5691 -6966 5694
rect -7012 5657 -7006 5691
rect -6972 5657 -6966 5691
rect -7012 5619 -6966 5657
rect -7012 5585 -7006 5619
rect -6972 5585 -6966 5619
rect -7012 5538 -6966 5585
rect -6754 5691 -6708 5729
rect -6511 5886 -6490 5901
rect -6456 5901 -6450 5907
rect -6238 6161 -6232 6168
rect -6198 6168 -6171 6180
rect -5980 6339 -5934 6377
rect -5722 7491 -5676 7538
rect -5722 7457 -5716 7491
rect -5682 7457 -5676 7491
rect -5722 7419 -5676 7457
rect -5722 7385 -5716 7419
rect -5682 7385 -5676 7419
rect -5722 7347 -5676 7385
rect -5722 7313 -5716 7347
rect -5682 7313 -5676 7347
rect -5722 7275 -5676 7313
rect -5722 7241 -5716 7275
rect -5682 7241 -5676 7275
rect -5722 7203 -5676 7241
rect -5722 7169 -5716 7203
rect -5682 7169 -5676 7203
rect -5722 7131 -5676 7169
rect -5722 7097 -5716 7131
rect -5682 7097 -5676 7131
rect -5722 7059 -5676 7097
rect -5722 7025 -5716 7059
rect -5682 7025 -5676 7059
rect -5722 6987 -5676 7025
rect -5722 6953 -5716 6987
rect -5682 6953 -5676 6987
rect -5722 6915 -5676 6953
rect -5722 6881 -5716 6915
rect -5682 6881 -5676 6915
rect -5722 6843 -5676 6881
rect -5722 6809 -5716 6843
rect -5682 6809 -5676 6843
rect -5722 6771 -5676 6809
rect -5722 6737 -5716 6771
rect -5682 6737 -5676 6771
rect -5722 6699 -5676 6737
rect -5722 6665 -5716 6699
rect -5682 6665 -5676 6699
rect -5722 6627 -5676 6665
rect -5722 6593 -5716 6627
rect -5682 6593 -5676 6627
rect -5722 6555 -5676 6593
rect -5722 6521 -5716 6555
rect -5682 6521 -5676 6555
rect -5722 6483 -5676 6521
rect -5722 6449 -5716 6483
rect -5682 6449 -5676 6483
rect -5722 6411 -5676 6449
rect -5722 6377 -5716 6411
rect -5682 6377 -5676 6411
rect -5722 6375 -5676 6377
rect -5464 7491 -5418 7538
rect -5464 7457 -5458 7491
rect -5424 7457 -5418 7491
rect -5464 7419 -5418 7457
rect -5464 7385 -5458 7419
rect -5424 7385 -5418 7419
rect -5464 7347 -5418 7385
rect -5464 7313 -5458 7347
rect -5424 7313 -5418 7347
rect -5464 7275 -5418 7313
rect -5464 7241 -5458 7275
rect -5424 7241 -5418 7275
rect -5464 7203 -5418 7241
rect -5464 7169 -5458 7203
rect -5424 7169 -5418 7203
rect -5464 7131 -5418 7169
rect -5464 7097 -5458 7131
rect -5424 7097 -5418 7131
rect -5464 7059 -5418 7097
rect -5464 7025 -5458 7059
rect -5424 7025 -5418 7059
rect -5464 6987 -5418 7025
rect -5464 6953 -5458 6987
rect -5424 6953 -5418 6987
rect -5464 6915 -5418 6953
rect -5464 6881 -5458 6915
rect -5424 6881 -5418 6915
rect -5464 6843 -5418 6881
rect -5464 6809 -5458 6843
rect -5424 6809 -5418 6843
rect -5464 6771 -5418 6809
rect -5464 6737 -5458 6771
rect -5424 6737 -5418 6771
rect -5464 6699 -5418 6737
rect -5464 6665 -5458 6699
rect -5424 6665 -5418 6699
rect -5464 6627 -5418 6665
rect -5464 6593 -5458 6627
rect -5424 6593 -5418 6627
rect -5464 6555 -5418 6593
rect -5464 6521 -5458 6555
rect -5424 6521 -5418 6555
rect -5464 6483 -5418 6521
rect -5464 6449 -5458 6483
rect -5424 6449 -5418 6483
rect -5464 6411 -5418 6449
rect -5464 6377 -5458 6411
rect -5424 6377 -5418 6411
rect -5980 6305 -5974 6339
rect -5940 6305 -5934 6339
rect -5980 6267 -5934 6305
rect -5980 6233 -5974 6267
rect -5940 6233 -5934 6267
rect -5980 6195 -5934 6233
rect -6198 6161 -6192 6168
rect -6238 6123 -6192 6161
rect -6238 6089 -6232 6123
rect -6198 6089 -6192 6123
rect -6238 6051 -6192 6089
rect -6238 6017 -6232 6051
rect -6198 6017 -6192 6051
rect -6238 5979 -6192 6017
rect -6238 5945 -6232 5979
rect -6198 5945 -6192 5979
rect -6238 5907 -6192 5945
rect -6456 5886 -6435 5901
rect -6511 5834 -6499 5886
rect -6447 5834 -6435 5886
rect -6511 5822 -6490 5834
rect -6456 5822 -6435 5834
rect -6511 5770 -6499 5822
rect -6447 5770 -6435 5822
rect -6511 5763 -6435 5770
rect -6511 5758 -6490 5763
rect -6456 5758 -6435 5763
rect -6511 5706 -6499 5758
rect -6447 5706 -6435 5758
rect -6511 5694 -6435 5706
rect -6238 5873 -6232 5907
rect -6198 5873 -6192 5907
rect -5980 6161 -5974 6195
rect -5940 6161 -5934 6195
rect -5746 6339 -5656 6375
rect -5746 6328 -5716 6339
rect -5682 6328 -5656 6339
rect -5746 6276 -5726 6328
rect -5674 6276 -5656 6328
rect -5746 6267 -5656 6276
rect -5746 6264 -5716 6267
rect -5682 6264 -5656 6267
rect -5746 6212 -5726 6264
rect -5674 6212 -5656 6264
rect -5746 6195 -5656 6212
rect -5746 6168 -5716 6195
rect -5980 6123 -5934 6161
rect -5980 6089 -5974 6123
rect -5940 6089 -5934 6123
rect -5980 6051 -5934 6089
rect -5980 6017 -5974 6051
rect -5940 6017 -5934 6051
rect -5980 5979 -5934 6017
rect -5980 5945 -5974 5979
rect -5940 5945 -5934 5979
rect -5980 5907 -5934 5945
rect -5980 5901 -5974 5907
rect -6238 5835 -6192 5873
rect -6238 5801 -6232 5835
rect -6198 5801 -6192 5835
rect -6238 5763 -6192 5801
rect -6238 5729 -6232 5763
rect -6198 5729 -6192 5763
rect -6754 5657 -6748 5691
rect -6714 5657 -6708 5691
rect -6754 5619 -6708 5657
rect -6754 5585 -6748 5619
rect -6714 5585 -6708 5619
rect -6754 5538 -6708 5585
rect -6496 5691 -6450 5694
rect -6496 5657 -6490 5691
rect -6456 5657 -6450 5691
rect -6496 5619 -6450 5657
rect -6496 5585 -6490 5619
rect -6456 5585 -6450 5619
rect -6496 5538 -6450 5585
rect -6238 5691 -6192 5729
rect -5997 5887 -5974 5901
rect -5940 5901 -5934 5907
rect -5722 6161 -5716 6168
rect -5682 6168 -5656 6195
rect -5464 6339 -5418 6377
rect -5206 7491 -5160 7538
rect -5206 7457 -5200 7491
rect -5166 7457 -5160 7491
rect -5206 7419 -5160 7457
rect -5206 7385 -5200 7419
rect -5166 7385 -5160 7419
rect -5206 7347 -5160 7385
rect -5206 7313 -5200 7347
rect -5166 7313 -5160 7347
rect -5206 7275 -5160 7313
rect -5206 7241 -5200 7275
rect -5166 7241 -5160 7275
rect -5206 7203 -5160 7241
rect -5206 7169 -5200 7203
rect -5166 7169 -5160 7203
rect -5206 7131 -5160 7169
rect -5206 7097 -5200 7131
rect -5166 7097 -5160 7131
rect -5206 7059 -5160 7097
rect -5206 7025 -5200 7059
rect -5166 7025 -5160 7059
rect -5206 6987 -5160 7025
rect -5206 6953 -5200 6987
rect -5166 6953 -5160 6987
rect -5206 6915 -5160 6953
rect -5206 6881 -5200 6915
rect -5166 6881 -5160 6915
rect -5206 6843 -5160 6881
rect -5206 6809 -5200 6843
rect -5166 6809 -5160 6843
rect -5206 6771 -5160 6809
rect -5206 6737 -5200 6771
rect -5166 6737 -5160 6771
rect -5206 6699 -5160 6737
rect -5206 6665 -5200 6699
rect -5166 6665 -5160 6699
rect -5206 6627 -5160 6665
rect -5206 6593 -5200 6627
rect -5166 6593 -5160 6627
rect -5206 6555 -5160 6593
rect -5206 6521 -5200 6555
rect -5166 6521 -5160 6555
rect -5206 6483 -5160 6521
rect -5206 6449 -5200 6483
rect -5166 6449 -5160 6483
rect -5206 6411 -5160 6449
rect -5206 6377 -5200 6411
rect -5166 6377 -5160 6411
rect -5206 6375 -5160 6377
rect -4948 7491 -4902 7538
rect -4948 7457 -4942 7491
rect -4908 7457 -4902 7491
rect -4948 7419 -4902 7457
rect -4948 7385 -4942 7419
rect -4908 7385 -4902 7419
rect -4948 7347 -4902 7385
rect -4948 7313 -4942 7347
rect -4908 7313 -4902 7347
rect -4948 7275 -4902 7313
rect -4948 7241 -4942 7275
rect -4908 7241 -4902 7275
rect -4948 7203 -4902 7241
rect -4948 7169 -4942 7203
rect -4908 7169 -4902 7203
rect -4948 7131 -4902 7169
rect -4948 7097 -4942 7131
rect -4908 7097 -4902 7131
rect -4948 7059 -4902 7097
rect -4948 7025 -4942 7059
rect -4908 7025 -4902 7059
rect -4948 6987 -4902 7025
rect -4948 6953 -4942 6987
rect -4908 6953 -4902 6987
rect -4948 6915 -4902 6953
rect -4948 6881 -4942 6915
rect -4908 6881 -4902 6915
rect -4948 6843 -4902 6881
rect -4948 6809 -4942 6843
rect -4908 6809 -4902 6843
rect -4948 6771 -4902 6809
rect -4948 6737 -4942 6771
rect -4908 6737 -4902 6771
rect -4948 6699 -4902 6737
rect -4948 6665 -4942 6699
rect -4908 6665 -4902 6699
rect -4948 6627 -4902 6665
rect -4948 6593 -4942 6627
rect -4908 6593 -4902 6627
rect -4948 6555 -4902 6593
rect -4948 6521 -4942 6555
rect -4908 6521 -4902 6555
rect -4948 6483 -4902 6521
rect -4948 6449 -4942 6483
rect -4908 6449 -4902 6483
rect -4948 6411 -4902 6449
rect -4948 6377 -4942 6411
rect -4908 6377 -4902 6411
rect -5464 6305 -5458 6339
rect -5424 6305 -5418 6339
rect -5464 6267 -5418 6305
rect -5464 6233 -5458 6267
rect -5424 6233 -5418 6267
rect -5464 6195 -5418 6233
rect -5682 6161 -5676 6168
rect -5722 6123 -5676 6161
rect -5722 6089 -5716 6123
rect -5682 6089 -5676 6123
rect -5722 6051 -5676 6089
rect -5722 6017 -5716 6051
rect -5682 6017 -5676 6051
rect -5722 5979 -5676 6017
rect -5722 5945 -5716 5979
rect -5682 5945 -5676 5979
rect -5722 5907 -5676 5945
rect -5940 5887 -5920 5901
rect -5997 5835 -5985 5887
rect -5933 5835 -5920 5887
rect -5997 5823 -5974 5835
rect -5940 5823 -5920 5835
rect -5997 5771 -5985 5823
rect -5933 5771 -5920 5823
rect -5997 5763 -5920 5771
rect -5997 5759 -5974 5763
rect -5940 5759 -5920 5763
rect -5997 5707 -5985 5759
rect -5933 5707 -5920 5759
rect -5997 5693 -5920 5707
rect -5722 5873 -5716 5907
rect -5682 5873 -5676 5907
rect -5464 6161 -5458 6195
rect -5424 6161 -5418 6195
rect -5227 6361 -5137 6375
rect -5227 6309 -5209 6361
rect -5157 6309 -5137 6361
rect -5227 6305 -5200 6309
rect -5166 6305 -5137 6309
rect -5227 6297 -5137 6305
rect -5227 6245 -5209 6297
rect -5157 6245 -5137 6297
rect -5227 6233 -5200 6245
rect -5166 6233 -5137 6245
rect -5227 6181 -5209 6233
rect -5157 6181 -5137 6233
rect -5227 6168 -5200 6181
rect -5464 6123 -5418 6161
rect -5464 6089 -5458 6123
rect -5424 6089 -5418 6123
rect -5464 6051 -5418 6089
rect -5464 6017 -5458 6051
rect -5424 6017 -5418 6051
rect -5464 5979 -5418 6017
rect -5464 5945 -5458 5979
rect -5424 5945 -5418 5979
rect -5464 5907 -5418 5945
rect -5464 5901 -5458 5907
rect -5722 5835 -5676 5873
rect -5722 5801 -5716 5835
rect -5682 5801 -5676 5835
rect -5722 5763 -5676 5801
rect -5722 5729 -5716 5763
rect -5682 5729 -5676 5763
rect -6238 5657 -6232 5691
rect -6198 5657 -6192 5691
rect -6238 5619 -6192 5657
rect -6238 5585 -6232 5619
rect -6198 5585 -6192 5619
rect -6238 5538 -6192 5585
rect -5980 5691 -5934 5693
rect -5980 5657 -5974 5691
rect -5940 5657 -5934 5691
rect -5980 5619 -5934 5657
rect -5980 5585 -5974 5619
rect -5940 5585 -5934 5619
rect -5980 5538 -5934 5585
rect -5722 5691 -5676 5729
rect -5483 5886 -5458 5901
rect -5424 5901 -5418 5907
rect -5206 6161 -5200 6168
rect -5166 6168 -5137 6181
rect -4948 6339 -4902 6377
rect -4690 7491 -4644 7538
rect -4690 7457 -4684 7491
rect -4650 7457 -4644 7491
rect -4690 7419 -4644 7457
rect -4690 7385 -4684 7419
rect -4650 7385 -4644 7419
rect -4690 7347 -4644 7385
rect -4690 7313 -4684 7347
rect -4650 7313 -4644 7347
rect -4690 7275 -4644 7313
rect -4690 7241 -4684 7275
rect -4650 7241 -4644 7275
rect -4690 7203 -4644 7241
rect -4690 7169 -4684 7203
rect -4650 7169 -4644 7203
rect -4690 7131 -4644 7169
rect -4690 7097 -4684 7131
rect -4650 7097 -4644 7131
rect -4690 7059 -4644 7097
rect -4690 7025 -4684 7059
rect -4650 7025 -4644 7059
rect -4690 6987 -4644 7025
rect -4690 6953 -4684 6987
rect -4650 6953 -4644 6987
rect -4690 6915 -4644 6953
rect -4690 6881 -4684 6915
rect -4650 6881 -4644 6915
rect -4690 6843 -4644 6881
rect -4690 6809 -4684 6843
rect -4650 6809 -4644 6843
rect -4690 6771 -4644 6809
rect -4690 6737 -4684 6771
rect -4650 6737 -4644 6771
rect -4690 6699 -4644 6737
rect -4690 6665 -4684 6699
rect -4650 6665 -4644 6699
rect -4690 6627 -4644 6665
rect -4690 6593 -4684 6627
rect -4650 6593 -4644 6627
rect -4690 6555 -4644 6593
rect -4690 6521 -4684 6555
rect -4650 6521 -4644 6555
rect -4690 6483 -4644 6521
rect -4690 6449 -4684 6483
rect -4650 6449 -4644 6483
rect -4690 6411 -4644 6449
rect -4690 6377 -4684 6411
rect -4650 6377 -4644 6411
rect -4690 6375 -4644 6377
rect -4432 7491 -4386 7538
rect -4432 7457 -4426 7491
rect -4392 7457 -4386 7491
rect -4432 7419 -4386 7457
rect -4432 7385 -4426 7419
rect -4392 7385 -4386 7419
rect -4432 7347 -4386 7385
rect -4432 7313 -4426 7347
rect -4392 7313 -4386 7347
rect -4432 7275 -4386 7313
rect -4432 7241 -4426 7275
rect -4392 7241 -4386 7275
rect -4432 7203 -4386 7241
rect -4432 7169 -4426 7203
rect -4392 7169 -4386 7203
rect -4432 7131 -4386 7169
rect -4432 7097 -4426 7131
rect -4392 7097 -4386 7131
rect -4432 7059 -4386 7097
rect -4432 7025 -4426 7059
rect -4392 7025 -4386 7059
rect -4432 6987 -4386 7025
rect -4432 6953 -4426 6987
rect -4392 6953 -4386 6987
rect -4432 6915 -4386 6953
rect -4432 6881 -4426 6915
rect -4392 6881 -4386 6915
rect -4432 6843 -4386 6881
rect -4432 6809 -4426 6843
rect -4392 6809 -4386 6843
rect -4174 7491 -4128 7538
rect -4174 7457 -4168 7491
rect -4134 7457 -4128 7491
rect -4174 7419 -4128 7457
rect -4174 7385 -4168 7419
rect -4134 7385 -4128 7419
rect -4174 7347 -4128 7385
rect -4174 7313 -4168 7347
rect -4134 7313 -4128 7347
rect -4174 7275 -4128 7313
rect -4174 7241 -4168 7275
rect -4134 7241 -4128 7275
rect -4174 7203 -4128 7241
rect -4174 7169 -4168 7203
rect -4134 7169 -4128 7203
rect -4174 7131 -4128 7169
rect -4174 7097 -4168 7131
rect -4134 7097 -4128 7131
rect -4174 7059 -4128 7097
rect -4174 7025 -4168 7059
rect -4134 7025 -4128 7059
rect -4174 6987 -4128 7025
rect -4174 6953 -4168 6987
rect -4134 6953 -4128 6987
rect -4174 6915 -4128 6953
rect -4174 6881 -4168 6915
rect -4134 6881 -4128 6915
rect -4174 6843 -4128 6881
rect -4174 6811 -4168 6843
rect -4432 6771 -4386 6809
rect -4432 6737 -4426 6771
rect -4392 6737 -4386 6771
rect -4432 6699 -4386 6737
rect -4432 6665 -4426 6699
rect -4392 6665 -4386 6699
rect -4432 6627 -4386 6665
rect -4432 6593 -4426 6627
rect -4392 6593 -4386 6627
rect -4194 6809 -4168 6811
rect -4134 6811 -4128 6843
rect -3916 7491 -3870 7538
rect -3916 7457 -3910 7491
rect -3876 7457 -3870 7491
rect -3916 7419 -3870 7457
rect -3916 7385 -3910 7419
rect -3876 7385 -3870 7419
rect -3916 7347 -3870 7385
rect -3916 7313 -3910 7347
rect -3876 7313 -3870 7347
rect -3916 7275 -3870 7313
rect -3916 7241 -3910 7275
rect -3876 7241 -3870 7275
rect -3916 7203 -3870 7241
rect -3916 7169 -3910 7203
rect -3876 7169 -3870 7203
rect -3916 7131 -3870 7169
rect -3916 7097 -3910 7131
rect -3876 7097 -3870 7131
rect -3916 7059 -3870 7097
rect -3916 7025 -3910 7059
rect -3876 7025 -3870 7059
rect -3916 6987 -3870 7025
rect -3916 6953 -3910 6987
rect -3876 6953 -3870 6987
rect -3916 6915 -3870 6953
rect -3916 6881 -3910 6915
rect -3876 6881 -3870 6915
rect -3916 6843 -3870 6881
rect -4134 6809 -4104 6811
rect -4194 6771 -4104 6809
rect -4194 6764 -4168 6771
rect -4134 6764 -4104 6771
rect -4194 6712 -4175 6764
rect -4123 6712 -4104 6764
rect -4194 6700 -4104 6712
rect -4194 6648 -4175 6700
rect -4123 6648 -4104 6700
rect -4194 6627 -4104 6648
rect -4194 6606 -4168 6627
rect -4432 6555 -4386 6593
rect -4432 6521 -4426 6555
rect -4392 6521 -4386 6555
rect -4432 6483 -4386 6521
rect -4432 6449 -4426 6483
rect -4392 6449 -4386 6483
rect -4432 6411 -4386 6449
rect -4432 6377 -4426 6411
rect -4392 6377 -4386 6411
rect -4948 6305 -4942 6339
rect -4908 6305 -4902 6339
rect -4948 6267 -4902 6305
rect -4948 6233 -4942 6267
rect -4908 6233 -4902 6267
rect -4948 6195 -4902 6233
rect -5166 6161 -5160 6168
rect -5206 6123 -5160 6161
rect -5206 6089 -5200 6123
rect -5166 6089 -5160 6123
rect -5206 6051 -5160 6089
rect -5206 6017 -5200 6051
rect -5166 6017 -5160 6051
rect -5206 5979 -5160 6017
rect -5206 5945 -5200 5979
rect -5166 5945 -5160 5979
rect -5206 5907 -5160 5945
rect -5424 5886 -5399 5901
rect -5483 5834 -5467 5886
rect -5415 5834 -5399 5886
rect -5483 5822 -5458 5834
rect -5424 5822 -5399 5834
rect -5483 5770 -5467 5822
rect -5415 5770 -5399 5822
rect -5483 5763 -5399 5770
rect -5483 5758 -5458 5763
rect -5424 5758 -5399 5763
rect -5483 5706 -5467 5758
rect -5415 5706 -5399 5758
rect -5483 5693 -5399 5706
rect -5206 5873 -5200 5907
rect -5166 5873 -5160 5907
rect -4948 6161 -4942 6195
rect -4908 6161 -4902 6195
rect -4708 6359 -4625 6375
rect -4708 6307 -4694 6359
rect -4642 6307 -4625 6359
rect -4708 6305 -4684 6307
rect -4650 6305 -4625 6307
rect -4708 6295 -4625 6305
rect -4708 6243 -4694 6295
rect -4642 6243 -4625 6295
rect -4708 6233 -4684 6243
rect -4650 6233 -4625 6243
rect -4708 6231 -4625 6233
rect -4708 6179 -4694 6231
rect -4642 6179 -4625 6231
rect -4708 6168 -4684 6179
rect -4948 6123 -4902 6161
rect -4948 6089 -4942 6123
rect -4908 6089 -4902 6123
rect -4948 6051 -4902 6089
rect -4948 6017 -4942 6051
rect -4908 6017 -4902 6051
rect -4948 5979 -4902 6017
rect -4948 5945 -4942 5979
rect -4908 5945 -4902 5979
rect -4948 5907 -4902 5945
rect -4948 5901 -4942 5907
rect -5206 5835 -5160 5873
rect -5206 5801 -5200 5835
rect -5166 5801 -5160 5835
rect -5206 5763 -5160 5801
rect -5206 5729 -5200 5763
rect -5166 5729 -5160 5763
rect -5722 5657 -5716 5691
rect -5682 5657 -5676 5691
rect -5722 5619 -5676 5657
rect -5722 5585 -5716 5619
rect -5682 5585 -5676 5619
rect -5722 5538 -5676 5585
rect -5464 5691 -5418 5693
rect -5464 5657 -5458 5691
rect -5424 5657 -5418 5691
rect -5464 5619 -5418 5657
rect -5464 5585 -5458 5619
rect -5424 5585 -5418 5619
rect -5464 5538 -5418 5585
rect -5206 5691 -5160 5729
rect -4965 5887 -4942 5901
rect -4908 5901 -4902 5907
rect -4690 6161 -4684 6168
rect -4650 6168 -4625 6179
rect -4432 6339 -4386 6377
rect -4432 6305 -4426 6339
rect -4392 6305 -4386 6339
rect -4432 6267 -4386 6305
rect -4432 6233 -4426 6267
rect -4392 6233 -4386 6267
rect -4432 6195 -4386 6233
rect -4650 6161 -4644 6168
rect -4690 6123 -4644 6161
rect -4690 6089 -4684 6123
rect -4650 6089 -4644 6123
rect -4690 6051 -4644 6089
rect -4690 6017 -4684 6051
rect -4650 6017 -4644 6051
rect -4690 5979 -4644 6017
rect -4690 5945 -4684 5979
rect -4650 5945 -4644 5979
rect -4690 5907 -4644 5945
rect -4908 5887 -4885 5901
rect -4965 5835 -4952 5887
rect -4900 5835 -4885 5887
rect -4965 5823 -4942 5835
rect -4908 5823 -4885 5835
rect -4965 5771 -4952 5823
rect -4900 5771 -4885 5823
rect -4965 5763 -4885 5771
rect -4965 5759 -4942 5763
rect -4908 5759 -4885 5763
rect -4965 5707 -4952 5759
rect -4900 5707 -4885 5759
rect -4965 5693 -4885 5707
rect -4690 5873 -4684 5907
rect -4650 5873 -4644 5907
rect -4432 6161 -4426 6195
rect -4392 6161 -4386 6195
rect -4432 6123 -4386 6161
rect -4432 6089 -4426 6123
rect -4392 6089 -4386 6123
rect -4432 6051 -4386 6089
rect -4432 6017 -4426 6051
rect -4392 6017 -4386 6051
rect -4432 5979 -4386 6017
rect -4432 5945 -4426 5979
rect -4392 5945 -4386 5979
rect -4432 5907 -4386 5945
rect -4432 5901 -4426 5907
rect -4690 5835 -4644 5873
rect -4690 5801 -4684 5835
rect -4650 5801 -4644 5835
rect -4690 5763 -4644 5801
rect -4690 5729 -4684 5763
rect -4650 5729 -4644 5763
rect -5206 5657 -5200 5691
rect -5166 5657 -5160 5691
rect -5206 5619 -5160 5657
rect -5206 5585 -5200 5619
rect -5166 5585 -5160 5619
rect -5206 5538 -5160 5585
rect -4948 5691 -4902 5693
rect -4948 5657 -4942 5691
rect -4908 5657 -4902 5691
rect -4948 5619 -4902 5657
rect -4948 5585 -4942 5619
rect -4908 5585 -4902 5619
rect -4948 5538 -4902 5585
rect -4690 5691 -4644 5729
rect -4449 5887 -4426 5901
rect -4392 5901 -4386 5907
rect -4174 6593 -4168 6606
rect -4134 6606 -4104 6627
rect -3916 6809 -3910 6843
rect -3876 6809 -3870 6843
rect -3658 7491 -3612 7538
rect 13111 7530 13142 7550
rect -3658 7457 -3652 7491
rect -3618 7457 -3612 7491
rect -3658 7419 -3612 7457
rect -3658 7385 -3652 7419
rect -3618 7385 -3612 7419
rect -3658 7347 -3612 7385
rect -3658 7313 -3652 7347
rect -3618 7313 -3612 7347
rect -3658 7275 -3612 7313
rect -3658 7241 -3652 7275
rect -3618 7241 -3612 7275
rect -3658 7203 -3612 7241
rect -3658 7169 -3652 7203
rect -3618 7169 -3612 7203
rect -3658 7131 -3612 7169
rect -3658 7097 -3652 7131
rect -3618 7097 -3612 7131
rect -3658 7059 -3612 7097
rect -3658 7025 -3652 7059
rect -3618 7025 -3612 7059
rect -3658 6987 -3612 7025
rect -3658 6953 -3652 6987
rect -3618 6953 -3612 6987
rect -3658 6915 -3612 6953
rect -3658 6881 -3652 6915
rect -3618 6881 -3612 6915
rect -3658 6843 -3612 6881
rect -3658 6811 -3652 6843
rect -3916 6771 -3870 6809
rect -3916 6737 -3910 6771
rect -3876 6737 -3870 6771
rect -3916 6699 -3870 6737
rect -3916 6665 -3910 6699
rect -3876 6665 -3870 6699
rect -3916 6627 -3870 6665
rect -4134 6593 -4128 6606
rect -4174 6555 -4128 6593
rect -4174 6521 -4168 6555
rect -4134 6521 -4128 6555
rect -4174 6483 -4128 6521
rect -4174 6449 -4168 6483
rect -4134 6449 -4128 6483
rect -4174 6411 -4128 6449
rect -4174 6377 -4168 6411
rect -4134 6377 -4128 6411
rect -4174 6339 -4128 6377
rect -4174 6305 -4168 6339
rect -4134 6305 -4128 6339
rect -4174 6267 -4128 6305
rect -4174 6233 -4168 6267
rect -4134 6233 -4128 6267
rect -4174 6195 -4128 6233
rect -4174 6161 -4168 6195
rect -4134 6161 -4128 6195
rect -4174 6123 -4128 6161
rect -4174 6089 -4168 6123
rect -4134 6089 -4128 6123
rect -4174 6051 -4128 6089
rect -4174 6017 -4168 6051
rect -4134 6017 -4128 6051
rect -4174 5979 -4128 6017
rect -4174 5945 -4168 5979
rect -4134 5945 -4128 5979
rect -4174 5907 -4128 5945
rect -4392 5887 -4370 5901
rect -4449 5835 -4435 5887
rect -4383 5835 -4370 5887
rect -4449 5823 -4426 5835
rect -4392 5823 -4370 5835
rect -4449 5771 -4435 5823
rect -4383 5771 -4370 5823
rect -4449 5763 -4370 5771
rect -4449 5759 -4426 5763
rect -4392 5759 -4370 5763
rect -4449 5707 -4435 5759
rect -4383 5707 -4370 5759
rect -4449 5693 -4370 5707
rect -4174 5873 -4168 5907
rect -4134 5873 -4128 5907
rect -3916 6593 -3910 6627
rect -3876 6593 -3870 6627
rect -3675 6809 -3652 6811
rect -3618 6811 -3612 6843
rect 13066 7516 13142 7530
rect 13176 7516 13242 7550
rect 13276 7516 13342 7550
rect 13376 7516 13442 7550
rect 13476 7516 13542 7550
rect 13576 7516 13642 7550
rect 13676 7530 13721 7550
rect 16412 7560 16652 7760
rect 16832 7633 16872 7877
rect 17052 7660 17082 7877
rect 17242 7910 17382 8420
rect 17446 8330 17468 8638
rect 17584 8330 17616 8638
rect 17446 8298 17616 8330
rect 17446 8294 17478 8298
rect 17472 8264 17478 8294
rect 17512 8294 17616 8298
rect 18530 8658 18576 8696
rect 19588 10890 20250 10928
rect 19588 10856 19594 10890
rect 19628 10856 20250 10890
rect 19588 10818 20250 10856
rect 19588 10784 19594 10818
rect 19628 10784 20250 10818
rect 19588 10746 20250 10784
rect 19588 10712 19594 10746
rect 19628 10712 20250 10746
rect 19588 10690 20250 10712
rect 19588 10674 20246 10690
rect 19588 10640 19594 10674
rect 19628 10654 20246 10674
rect 19628 10650 19876 10654
rect 19628 10640 19634 10650
rect 19588 10602 19634 10640
rect 19588 10568 19594 10602
rect 19628 10568 19634 10602
rect 19588 10530 19634 10568
rect 19588 10496 19594 10530
rect 19628 10496 19634 10530
rect 19588 10458 19634 10496
rect 19588 10424 19594 10458
rect 19628 10424 19634 10458
rect 19588 10386 19634 10424
rect 19588 10352 19594 10386
rect 19628 10352 19634 10386
rect 19588 10314 19634 10352
rect 19588 10280 19594 10314
rect 19628 10280 19634 10314
rect 19588 10242 19634 10280
rect 19588 10208 19594 10242
rect 19628 10208 19634 10242
rect 19588 10170 19634 10208
rect 19588 10136 19594 10170
rect 19628 10136 19634 10170
rect 19588 10098 19634 10136
rect 19588 10064 19594 10098
rect 19628 10064 19634 10098
rect 19588 10026 19634 10064
rect 19588 9992 19594 10026
rect 19628 9992 19634 10026
rect 19588 9954 19634 9992
rect 19588 9920 19594 9954
rect 19628 9920 19634 9954
rect 19588 9882 19634 9920
rect 19588 9848 19594 9882
rect 19628 9848 19634 9882
rect 19588 9810 19634 9848
rect 19588 9776 19594 9810
rect 19628 9776 19634 9810
rect 19588 9738 19634 9776
rect 19588 9704 19594 9738
rect 19628 9704 19634 9738
rect 19588 9666 19634 9704
rect 19588 9632 19594 9666
rect 19628 9632 19634 9666
rect 19588 9594 19634 9632
rect 19588 9560 19594 9594
rect 19628 9560 19634 9594
rect 19588 9522 19634 9560
rect 19588 9488 19594 9522
rect 19628 9488 19634 9522
rect 19588 9450 19634 9488
rect 19588 9416 19594 9450
rect 19628 9416 19634 9450
rect 19588 9378 19634 9416
rect 19588 9344 19594 9378
rect 19628 9344 19634 9378
rect 19588 9306 19634 9344
rect 19588 9272 19594 9306
rect 19628 9272 19634 9306
rect 19588 9234 19634 9272
rect 19588 9200 19594 9234
rect 19628 9200 19634 9234
rect 19588 9162 19634 9200
rect 19588 9128 19594 9162
rect 19628 9128 19634 9162
rect 19588 9090 19634 9128
rect 19588 9056 19594 9090
rect 19628 9056 19634 9090
rect 19588 9018 19634 9056
rect 19588 8984 19594 9018
rect 19628 8984 19634 9018
rect 21086 9398 21300 14056
rect 21476 14450 21526 14464
rect 21476 14416 21484 14450
rect 21518 14416 21526 14450
rect 21476 14378 21526 14416
rect 21476 14344 21484 14378
rect 21518 14344 21526 14378
rect 21476 14306 21526 14344
rect 21476 14272 21484 14306
rect 21518 14272 21526 14306
rect 21476 14234 21526 14272
rect 21476 14200 21484 14234
rect 21518 14200 21526 14234
rect 21476 14162 21526 14200
rect 21476 14128 21484 14162
rect 21518 14128 21526 14162
rect 21476 14090 21526 14128
rect 21476 14056 21484 14090
rect 21518 14056 21526 14090
rect 21476 14043 21526 14056
rect 28974 14171 29024 14185
rect 28974 14137 28982 14171
rect 29016 14137 29024 14171
rect 28974 14099 29024 14137
rect 28974 14065 28982 14099
rect 29016 14065 29024 14099
rect 28974 14027 29024 14065
rect 28974 13993 28982 14027
rect 29016 13993 29024 14027
rect 28974 13955 29024 13993
rect 28974 13921 28982 13955
rect 29016 13921 29024 13955
rect 28974 13883 29024 13921
rect 28974 13849 28982 13883
rect 29016 13849 29024 13883
rect 28974 13811 29024 13849
rect 28974 13777 28982 13811
rect 29016 13777 29024 13811
rect 28974 13764 29024 13777
rect 29200 14171 29466 14204
rect 29200 14137 29300 14171
rect 29334 14137 29466 14171
rect 29200 14099 29466 14137
rect 29200 14065 29300 14099
rect 29334 14065 29466 14099
rect 29200 14027 29466 14065
rect 29200 13993 29300 14027
rect 29334 13993 29466 14027
rect 29200 13955 29466 13993
rect 29200 13921 29300 13955
rect 29334 13921 29466 13955
rect 29200 13883 29466 13921
rect 29200 13849 29300 13883
rect 29334 13849 29466 13883
rect 29200 13811 29466 13849
rect 29200 13777 29300 13811
rect 29334 13777 29466 13811
rect 29200 13673 29466 13777
rect 29610 14171 29660 14185
rect 29610 14137 29618 14171
rect 29652 14137 29660 14171
rect 29610 14099 29660 14137
rect 29610 14065 29618 14099
rect 29652 14065 29660 14099
rect 29610 14027 29660 14065
rect 29610 13993 29618 14027
rect 29652 13993 29660 14027
rect 29610 13955 29660 13993
rect 29610 13921 29618 13955
rect 29652 13921 29660 13955
rect 29610 13883 29660 13921
rect 29610 13849 29618 13883
rect 29652 13849 29660 13883
rect 29610 13811 29660 13849
rect 29610 13777 29618 13811
rect 29652 13777 29660 13811
rect 29610 13764 29660 13777
rect 36395 13673 36661 15695
rect 38454 15653 38878 15747
rect 38454 15652 38877 15653
rect 39497 15625 39895 15747
rect 40126 15694 40366 15714
rect 40126 15642 40155 15694
rect 40207 15642 40219 15694
rect 40271 15642 40283 15694
rect 40335 15642 40366 15694
rect 40531 15659 40679 15747
rect 40126 15624 40366 15642
rect 41643 15635 41816 16686
rect 41643 15601 41730 15635
rect 41764 15601 41816 15635
rect 38127 15538 38173 15585
rect 38127 15504 38133 15538
rect 38167 15504 38173 15538
rect 38127 15466 38173 15504
rect 38127 15432 38133 15466
rect 38167 15432 38173 15466
rect 38127 15394 38173 15432
rect 38127 15360 38133 15394
rect 38167 15360 38173 15394
rect 38127 15322 38173 15360
rect 38127 15288 38133 15322
rect 38167 15288 38173 15322
rect 38127 15250 38173 15288
rect 38127 15216 38133 15250
rect 38167 15216 38173 15250
rect 38127 15178 38173 15216
rect 38127 15144 38133 15178
rect 38167 15144 38173 15178
rect 38127 15106 38173 15144
rect 38127 15072 38133 15106
rect 38167 15072 38173 15106
rect 38127 15034 38173 15072
rect 38127 15000 38133 15034
rect 38167 15000 38173 15034
rect 38127 14962 38173 15000
rect 38127 14928 38133 14962
rect 38167 14928 38173 14962
rect 38127 14890 38173 14928
rect 38127 14856 38133 14890
rect 38167 14856 38173 14890
rect 38127 14818 38173 14856
rect 38127 14784 38133 14818
rect 38167 14784 38173 14818
rect 38127 14746 38173 14784
rect 38127 14712 38133 14746
rect 38167 14712 38173 14746
rect 38127 14674 38173 14712
rect 38127 14640 38133 14674
rect 38167 14640 38173 14674
rect 38127 14602 38173 14640
rect 38127 14568 38133 14602
rect 38167 14568 38173 14602
rect 38127 14530 38173 14568
rect 38127 14496 38133 14530
rect 38167 14496 38173 14530
rect 38127 14458 38173 14496
rect 38127 14424 38133 14458
rect 38167 14424 38173 14458
rect 38127 14386 38173 14424
rect 38127 14352 38133 14386
rect 38167 14352 38173 14386
rect 38127 14314 38173 14352
rect 38127 14280 38133 14314
rect 38167 14280 38173 14314
rect 38127 14242 38173 14280
rect 38127 14208 38133 14242
rect 38167 14208 38173 14242
rect 38127 14170 38173 14208
rect 38127 14136 38133 14170
rect 38167 14136 38173 14170
rect 38127 14098 38173 14136
rect 38127 14064 38133 14098
rect 38167 14064 38173 14098
rect 38127 14026 38173 14064
rect 38127 13992 38133 14026
rect 38167 13992 38173 14026
rect 38127 13954 38173 13992
rect 38127 13920 38133 13954
rect 38167 13920 38173 13954
rect 38127 13882 38173 13920
rect 38127 13869 38133 13882
rect 38092 13848 38133 13869
rect 38167 13869 38173 13882
rect 38385 15538 38431 15585
rect 38643 15572 38689 15585
rect 38385 15504 38391 15538
rect 38425 15504 38431 15538
rect 38385 15466 38431 15504
rect 38385 15432 38391 15466
rect 38425 15432 38431 15466
rect 38385 15394 38431 15432
rect 38385 15360 38391 15394
rect 38425 15360 38431 15394
rect 38385 15322 38431 15360
rect 38385 15288 38391 15322
rect 38425 15288 38431 15322
rect 38385 15250 38431 15288
rect 38598 15538 38748 15572
rect 38598 15518 38649 15538
rect 38683 15518 38748 15538
rect 38598 15466 38645 15518
rect 38697 15466 38748 15518
rect 38598 15454 38649 15466
rect 38683 15454 38748 15466
rect 38598 15402 38645 15454
rect 38697 15402 38748 15454
rect 38598 15394 38748 15402
rect 38598 15390 38649 15394
rect 38683 15390 38748 15394
rect 38598 15338 38645 15390
rect 38697 15338 38748 15390
rect 38598 15322 38748 15338
rect 38598 15288 38649 15322
rect 38683 15288 38748 15322
rect 38598 15286 38748 15288
rect 38901 15538 38947 15585
rect 38901 15504 38907 15538
rect 38941 15504 38947 15538
rect 38901 15466 38947 15504
rect 38901 15432 38907 15466
rect 38941 15432 38947 15466
rect 38901 15394 38947 15432
rect 38901 15360 38907 15394
rect 38941 15360 38947 15394
rect 38901 15322 38947 15360
rect 38901 15288 38907 15322
rect 38941 15288 38947 15322
rect 38385 15216 38391 15250
rect 38425 15216 38431 15250
rect 38385 15178 38431 15216
rect 38385 15144 38391 15178
rect 38425 15144 38431 15178
rect 38385 15106 38431 15144
rect 38385 15072 38391 15106
rect 38425 15072 38431 15106
rect 38385 15034 38431 15072
rect 38385 15000 38391 15034
rect 38425 15000 38431 15034
rect 38385 14962 38431 15000
rect 38385 14928 38391 14962
rect 38425 14928 38431 14962
rect 38385 14890 38431 14928
rect 38385 14856 38391 14890
rect 38425 14856 38431 14890
rect 38385 14818 38431 14856
rect 38385 14784 38391 14818
rect 38425 14784 38431 14818
rect 38385 14746 38431 14784
rect 38385 14712 38391 14746
rect 38425 14712 38431 14746
rect 38385 14674 38431 14712
rect 38385 14640 38391 14674
rect 38425 14640 38431 14674
rect 38385 14602 38431 14640
rect 38385 14568 38391 14602
rect 38425 14568 38431 14602
rect 38385 14530 38431 14568
rect 38385 14496 38391 14530
rect 38425 14496 38431 14530
rect 38385 14458 38431 14496
rect 38385 14424 38391 14458
rect 38425 14424 38431 14458
rect 38385 14386 38431 14424
rect 38385 14352 38391 14386
rect 38425 14352 38431 14386
rect 38385 14314 38431 14352
rect 38385 14280 38391 14314
rect 38425 14280 38431 14314
rect 38385 14242 38431 14280
rect 38385 14208 38391 14242
rect 38425 14208 38431 14242
rect 38385 14170 38431 14208
rect 38385 14136 38391 14170
rect 38425 14136 38431 14170
rect 38385 14098 38431 14136
rect 38385 14064 38391 14098
rect 38425 14064 38431 14098
rect 38385 14026 38431 14064
rect 38385 13992 38391 14026
rect 38425 13992 38431 14026
rect 38385 13954 38431 13992
rect 38385 13920 38391 13954
rect 38425 13920 38431 13954
rect 38385 13882 38431 13920
rect 38167 13848 38242 13869
rect 38092 13815 38242 13848
rect 38092 13810 38139 13815
rect 38092 13776 38133 13810
rect 38092 13763 38139 13776
rect 38191 13763 38242 13815
rect 38092 13751 38242 13763
rect 38092 13738 38139 13751
rect 38092 13704 38133 13738
rect 38092 13699 38139 13704
rect 38191 13699 38242 13751
rect 38092 13687 38242 13699
rect 29200 13407 36662 13673
rect 38092 13666 38139 13687
rect 38092 13632 38133 13666
rect 38191 13635 38242 13687
rect 38167 13632 38242 13635
rect 38092 13583 38242 13632
rect 38385 13848 38391 13882
rect 38425 13848 38431 13882
rect 38385 13810 38431 13848
rect 38385 13776 38391 13810
rect 38425 13776 38431 13810
rect 38385 13738 38431 13776
rect 38385 13704 38391 13738
rect 38425 13704 38431 13738
rect 38385 13666 38431 13704
rect 38385 13632 38391 13666
rect 38425 13632 38431 13666
rect 38385 13585 38431 13632
rect 38643 15250 38689 15286
rect 38643 15216 38649 15250
rect 38683 15216 38689 15250
rect 38643 15178 38689 15216
rect 38643 15144 38649 15178
rect 38683 15144 38689 15178
rect 38643 15106 38689 15144
rect 38643 15072 38649 15106
rect 38683 15072 38689 15106
rect 38643 15034 38689 15072
rect 38643 15000 38649 15034
rect 38683 15000 38689 15034
rect 38643 14962 38689 15000
rect 38643 14928 38649 14962
rect 38683 14928 38689 14962
rect 38643 14890 38689 14928
rect 38643 14856 38649 14890
rect 38683 14856 38689 14890
rect 38643 14818 38689 14856
rect 38643 14784 38649 14818
rect 38683 14784 38689 14818
rect 38643 14746 38689 14784
rect 38643 14712 38649 14746
rect 38683 14712 38689 14746
rect 38643 14674 38689 14712
rect 38643 14640 38649 14674
rect 38683 14640 38689 14674
rect 38643 14602 38689 14640
rect 38643 14568 38649 14602
rect 38683 14568 38689 14602
rect 38643 14530 38689 14568
rect 38643 14496 38649 14530
rect 38683 14496 38689 14530
rect 38643 14458 38689 14496
rect 38643 14424 38649 14458
rect 38683 14424 38689 14458
rect 38643 14386 38689 14424
rect 38643 14352 38649 14386
rect 38683 14352 38689 14386
rect 38643 14314 38689 14352
rect 38643 14280 38649 14314
rect 38683 14280 38689 14314
rect 38643 14242 38689 14280
rect 38643 14208 38649 14242
rect 38683 14208 38689 14242
rect 38643 14170 38689 14208
rect 38643 14136 38649 14170
rect 38683 14136 38689 14170
rect 38643 14098 38689 14136
rect 38643 14064 38649 14098
rect 38683 14064 38689 14098
rect 38643 14026 38689 14064
rect 38643 13992 38649 14026
rect 38683 13992 38689 14026
rect 38643 13954 38689 13992
rect 38643 13920 38649 13954
rect 38683 13920 38689 13954
rect 38643 13882 38689 13920
rect 38643 13848 38649 13882
rect 38683 13848 38689 13882
rect 38643 13810 38689 13848
rect 38643 13776 38649 13810
rect 38683 13776 38689 13810
rect 38643 13738 38689 13776
rect 38643 13704 38649 13738
rect 38683 13704 38689 13738
rect 38643 13666 38689 13704
rect 38643 13632 38649 13666
rect 38683 13632 38689 13666
rect 38643 13585 38689 13632
rect 38901 15250 38947 15288
rect 38901 15216 38907 15250
rect 38941 15216 38947 15250
rect 38901 15178 38947 15216
rect 38901 15144 38907 15178
rect 38941 15144 38947 15178
rect 38901 15106 38947 15144
rect 38901 15072 38907 15106
rect 38941 15072 38947 15106
rect 38901 15034 38947 15072
rect 38901 15000 38907 15034
rect 38941 15000 38947 15034
rect 38901 14962 38947 15000
rect 38901 14928 38907 14962
rect 38941 14928 38947 14962
rect 38901 14890 38947 14928
rect 38901 14856 38907 14890
rect 38941 14856 38947 14890
rect 38901 14818 38947 14856
rect 38901 14784 38907 14818
rect 38941 14784 38947 14818
rect 38901 14746 38947 14784
rect 38901 14712 38907 14746
rect 38941 14712 38947 14746
rect 38901 14674 38947 14712
rect 38901 14640 38907 14674
rect 38941 14640 38947 14674
rect 38901 14602 38947 14640
rect 38901 14568 38907 14602
rect 38941 14568 38947 14602
rect 38901 14530 38947 14568
rect 38901 14496 38907 14530
rect 38941 14496 38947 14530
rect 38901 14458 38947 14496
rect 38901 14424 38907 14458
rect 38941 14424 38947 14458
rect 38901 14386 38947 14424
rect 38901 14352 38907 14386
rect 38941 14352 38947 14386
rect 38901 14314 38947 14352
rect 38901 14280 38907 14314
rect 38941 14280 38947 14314
rect 38901 14242 38947 14280
rect 38901 14208 38907 14242
rect 38941 14208 38947 14242
rect 38901 14170 38947 14208
rect 38901 14136 38907 14170
rect 38941 14136 38947 14170
rect 38901 14098 38947 14136
rect 38901 14064 38907 14098
rect 38941 14064 38947 14098
rect 38901 14026 38947 14064
rect 38901 13992 38907 14026
rect 38941 13992 38947 14026
rect 38901 13954 38947 13992
rect 38901 13920 38907 13954
rect 38941 13920 38947 13954
rect 38901 13882 38947 13920
rect 38901 13848 38907 13882
rect 38941 13848 38947 13882
rect 39159 15538 39205 15585
rect 39159 15504 39165 15538
rect 39199 15504 39205 15538
rect 39159 15466 39205 15504
rect 39159 15432 39165 15466
rect 39199 15432 39205 15466
rect 39159 15394 39205 15432
rect 39159 15360 39165 15394
rect 39199 15360 39205 15394
rect 39159 15322 39205 15360
rect 39159 15288 39165 15322
rect 39199 15288 39205 15322
rect 39159 15250 39205 15288
rect 39159 15216 39165 15250
rect 39199 15216 39205 15250
rect 39159 15178 39205 15216
rect 39159 15144 39165 15178
rect 39199 15144 39205 15178
rect 39159 15106 39205 15144
rect 39159 15072 39165 15106
rect 39199 15072 39205 15106
rect 39159 15034 39205 15072
rect 39159 15000 39165 15034
rect 39199 15000 39205 15034
rect 39159 14962 39205 15000
rect 39159 14928 39165 14962
rect 39199 14928 39205 14962
rect 39159 14890 39205 14928
rect 39159 14856 39165 14890
rect 39199 14856 39205 14890
rect 39159 14818 39205 14856
rect 39159 14784 39165 14818
rect 39199 14784 39205 14818
rect 39159 14746 39205 14784
rect 39159 14712 39165 14746
rect 39199 14712 39205 14746
rect 39159 14674 39205 14712
rect 39159 14640 39165 14674
rect 39199 14640 39205 14674
rect 39159 14602 39205 14640
rect 39159 14568 39165 14602
rect 39199 14568 39205 14602
rect 39159 14530 39205 14568
rect 39159 14496 39165 14530
rect 39199 14496 39205 14530
rect 39159 14458 39205 14496
rect 39159 14424 39165 14458
rect 39199 14424 39205 14458
rect 39159 14386 39205 14424
rect 39159 14352 39165 14386
rect 39199 14352 39205 14386
rect 39159 14314 39205 14352
rect 39159 14280 39165 14314
rect 39199 14280 39205 14314
rect 39159 14242 39205 14280
rect 39159 14208 39165 14242
rect 39199 14208 39205 14242
rect 39159 14170 39205 14208
rect 39159 14136 39165 14170
rect 39199 14136 39205 14170
rect 39159 14098 39205 14136
rect 39159 14064 39165 14098
rect 39199 14064 39205 14098
rect 39159 14026 39205 14064
rect 39159 13992 39165 14026
rect 39199 13992 39205 14026
rect 39159 13954 39205 13992
rect 39159 13920 39165 13954
rect 39199 13920 39205 13954
rect 39159 13882 39205 13920
rect 39159 13880 39165 13882
rect 38901 13810 38947 13848
rect 38901 13776 38907 13810
rect 38941 13776 38947 13810
rect 38901 13738 38947 13776
rect 38901 13704 38907 13738
rect 38941 13704 38947 13738
rect 38901 13666 38947 13704
rect 38901 13632 38907 13666
rect 38941 13632 38947 13666
rect 38901 13585 38947 13632
rect 39111 13848 39165 13880
rect 39199 13880 39205 13882
rect 39417 15538 39463 15585
rect 39675 15559 39721 15585
rect 39417 15504 39423 15538
rect 39457 15504 39463 15538
rect 39417 15466 39463 15504
rect 39417 15432 39423 15466
rect 39457 15432 39463 15466
rect 39417 15394 39463 15432
rect 39417 15360 39423 15394
rect 39457 15360 39463 15394
rect 39417 15322 39463 15360
rect 39417 15288 39423 15322
rect 39457 15288 39463 15322
rect 39417 15250 39463 15288
rect 39609 15538 39759 15559
rect 39609 15505 39681 15538
rect 39609 15453 39656 15505
rect 39715 15504 39759 15538
rect 39708 15466 39759 15504
rect 39609 15441 39681 15453
rect 39609 15389 39656 15441
rect 39715 15432 39759 15466
rect 39708 15394 39759 15432
rect 39609 15377 39681 15389
rect 39609 15325 39656 15377
rect 39715 15360 39759 15394
rect 39708 15325 39759 15360
rect 39609 15322 39759 15325
rect 39609 15288 39681 15322
rect 39715 15288 39759 15322
rect 39609 15273 39759 15288
rect 39933 15538 39979 15585
rect 39933 15504 39939 15538
rect 39973 15504 39979 15538
rect 39933 15466 39979 15504
rect 39933 15432 39939 15466
rect 39973 15432 39979 15466
rect 39933 15394 39979 15432
rect 39933 15360 39939 15394
rect 39973 15360 39979 15394
rect 39933 15322 39979 15360
rect 39933 15288 39939 15322
rect 39973 15288 39979 15322
rect 39417 15216 39423 15250
rect 39457 15216 39463 15250
rect 39417 15178 39463 15216
rect 39417 15144 39423 15178
rect 39457 15144 39463 15178
rect 39417 15106 39463 15144
rect 39417 15072 39423 15106
rect 39457 15072 39463 15106
rect 39417 15034 39463 15072
rect 39417 15000 39423 15034
rect 39457 15000 39463 15034
rect 39417 14962 39463 15000
rect 39417 14928 39423 14962
rect 39457 14928 39463 14962
rect 39417 14890 39463 14928
rect 39417 14856 39423 14890
rect 39457 14856 39463 14890
rect 39417 14818 39463 14856
rect 39417 14784 39423 14818
rect 39457 14784 39463 14818
rect 39417 14746 39463 14784
rect 39417 14712 39423 14746
rect 39457 14712 39463 14746
rect 39417 14674 39463 14712
rect 39417 14640 39423 14674
rect 39457 14640 39463 14674
rect 39417 14602 39463 14640
rect 39417 14568 39423 14602
rect 39457 14568 39463 14602
rect 39417 14530 39463 14568
rect 39417 14496 39423 14530
rect 39457 14496 39463 14530
rect 39417 14458 39463 14496
rect 39417 14424 39423 14458
rect 39457 14424 39463 14458
rect 39417 14386 39463 14424
rect 39417 14352 39423 14386
rect 39457 14352 39463 14386
rect 39417 14314 39463 14352
rect 39417 14280 39423 14314
rect 39457 14280 39463 14314
rect 39417 14242 39463 14280
rect 39417 14208 39423 14242
rect 39457 14208 39463 14242
rect 39417 14170 39463 14208
rect 39417 14136 39423 14170
rect 39457 14136 39463 14170
rect 39417 14098 39463 14136
rect 39417 14064 39423 14098
rect 39457 14064 39463 14098
rect 39417 14026 39463 14064
rect 39417 13992 39423 14026
rect 39457 13992 39463 14026
rect 39417 13954 39463 13992
rect 39417 13920 39423 13954
rect 39457 13920 39463 13954
rect 39417 13882 39463 13920
rect 39199 13848 39261 13880
rect 39111 13826 39261 13848
rect 39111 13774 39158 13826
rect 39210 13774 39261 13826
rect 39111 13762 39261 13774
rect 39111 13710 39158 13762
rect 39210 13710 39261 13762
rect 39111 13704 39165 13710
rect 39199 13704 39261 13710
rect 39111 13698 39261 13704
rect 39111 13646 39158 13698
rect 39210 13646 39261 13698
rect 39111 13632 39165 13646
rect 39199 13632 39261 13646
rect 39111 13594 39261 13632
rect 39417 13848 39423 13882
rect 39457 13848 39463 13882
rect 39417 13810 39463 13848
rect 39417 13776 39423 13810
rect 39457 13776 39463 13810
rect 39417 13738 39463 13776
rect 39417 13704 39423 13738
rect 39457 13704 39463 13738
rect 39417 13666 39463 13704
rect 39417 13632 39423 13666
rect 39457 13632 39463 13666
rect 39159 13585 39205 13594
rect 39417 13585 39463 13632
rect 39675 15250 39721 15273
rect 39675 15216 39681 15250
rect 39715 15216 39721 15250
rect 39675 15178 39721 15216
rect 39675 15144 39681 15178
rect 39715 15144 39721 15178
rect 39675 15106 39721 15144
rect 39675 15072 39681 15106
rect 39715 15072 39721 15106
rect 39675 15034 39721 15072
rect 39675 15000 39681 15034
rect 39715 15000 39721 15034
rect 39675 14962 39721 15000
rect 39675 14928 39681 14962
rect 39715 14928 39721 14962
rect 39675 14890 39721 14928
rect 39675 14856 39681 14890
rect 39715 14856 39721 14890
rect 39675 14818 39721 14856
rect 39675 14784 39681 14818
rect 39715 14784 39721 14818
rect 39675 14746 39721 14784
rect 39675 14712 39681 14746
rect 39715 14712 39721 14746
rect 39675 14674 39721 14712
rect 39675 14640 39681 14674
rect 39715 14640 39721 14674
rect 39675 14602 39721 14640
rect 39675 14568 39681 14602
rect 39715 14568 39721 14602
rect 39675 14530 39721 14568
rect 39675 14496 39681 14530
rect 39715 14496 39721 14530
rect 39675 14458 39721 14496
rect 39675 14424 39681 14458
rect 39715 14424 39721 14458
rect 39675 14386 39721 14424
rect 39675 14352 39681 14386
rect 39715 14352 39721 14386
rect 39675 14314 39721 14352
rect 39675 14280 39681 14314
rect 39715 14280 39721 14314
rect 39675 14242 39721 14280
rect 39675 14208 39681 14242
rect 39715 14208 39721 14242
rect 39675 14170 39721 14208
rect 39675 14136 39681 14170
rect 39715 14136 39721 14170
rect 39675 14098 39721 14136
rect 39675 14064 39681 14098
rect 39715 14064 39721 14098
rect 39675 14026 39721 14064
rect 39675 13992 39681 14026
rect 39715 13992 39721 14026
rect 39675 13954 39721 13992
rect 39675 13920 39681 13954
rect 39715 13920 39721 13954
rect 39675 13882 39721 13920
rect 39675 13848 39681 13882
rect 39715 13848 39721 13882
rect 39675 13810 39721 13848
rect 39675 13776 39681 13810
rect 39715 13776 39721 13810
rect 39675 13738 39721 13776
rect 39675 13704 39681 13738
rect 39715 13704 39721 13738
rect 39675 13666 39721 13704
rect 39675 13632 39681 13666
rect 39715 13632 39721 13666
rect 39675 13585 39721 13632
rect 39933 15250 39979 15288
rect 39933 15216 39939 15250
rect 39973 15216 39979 15250
rect 39933 15178 39979 15216
rect 39933 15144 39939 15178
rect 39973 15144 39979 15178
rect 39933 15106 39979 15144
rect 39933 15072 39939 15106
rect 39973 15072 39979 15106
rect 39933 15034 39979 15072
rect 39933 15000 39939 15034
rect 39973 15000 39979 15034
rect 39933 14962 39979 15000
rect 39933 14928 39939 14962
rect 39973 14928 39979 14962
rect 39933 14890 39979 14928
rect 39933 14856 39939 14890
rect 39973 14856 39979 14890
rect 39933 14818 39979 14856
rect 39933 14784 39939 14818
rect 39973 14784 39979 14818
rect 39933 14746 39979 14784
rect 39933 14712 39939 14746
rect 39973 14712 39979 14746
rect 39933 14674 39979 14712
rect 39933 14640 39939 14674
rect 39973 14640 39979 14674
rect 39933 14602 39979 14640
rect 39933 14568 39939 14602
rect 39973 14568 39979 14602
rect 39933 14530 39979 14568
rect 39933 14496 39939 14530
rect 39973 14496 39979 14530
rect 39933 14458 39979 14496
rect 39933 14424 39939 14458
rect 39973 14424 39979 14458
rect 39933 14386 39979 14424
rect 39933 14352 39939 14386
rect 39973 14352 39979 14386
rect 39933 14314 39979 14352
rect 39933 14280 39939 14314
rect 39973 14280 39979 14314
rect 39933 14242 39979 14280
rect 39933 14208 39939 14242
rect 39973 14208 39979 14242
rect 39933 14170 39979 14208
rect 39933 14136 39939 14170
rect 39973 14136 39979 14170
rect 39933 14098 39979 14136
rect 39933 14064 39939 14098
rect 39973 14064 39979 14098
rect 39933 14026 39979 14064
rect 39933 13992 39939 14026
rect 39973 13992 39979 14026
rect 39933 13954 39979 13992
rect 39933 13920 39939 13954
rect 39973 13920 39979 13954
rect 39933 13882 39979 13920
rect 40191 15538 40237 15585
rect 40191 15504 40197 15538
rect 40231 15504 40237 15538
rect 40191 15466 40237 15504
rect 40191 15432 40197 15466
rect 40231 15432 40237 15466
rect 40191 15394 40237 15432
rect 40191 15360 40197 15394
rect 40231 15360 40237 15394
rect 40191 15322 40237 15360
rect 40191 15288 40197 15322
rect 40231 15288 40237 15322
rect 40191 15250 40237 15288
rect 40191 15216 40197 15250
rect 40231 15216 40237 15250
rect 40191 15178 40237 15216
rect 40191 15144 40197 15178
rect 40231 15144 40237 15178
rect 40191 15106 40237 15144
rect 40191 15072 40197 15106
rect 40231 15072 40237 15106
rect 40191 15034 40237 15072
rect 40191 15000 40197 15034
rect 40231 15000 40237 15034
rect 40191 14962 40237 15000
rect 40191 14928 40197 14962
rect 40231 14928 40237 14962
rect 40191 14890 40237 14928
rect 40191 14856 40197 14890
rect 40231 14856 40237 14890
rect 40191 14818 40237 14856
rect 40191 14784 40197 14818
rect 40231 14784 40237 14818
rect 40191 14746 40237 14784
rect 40191 14712 40197 14746
rect 40231 14712 40237 14746
rect 40191 14674 40237 14712
rect 40191 14640 40197 14674
rect 40231 14640 40237 14674
rect 40191 14602 40237 14640
rect 40191 14568 40197 14602
rect 40231 14568 40237 14602
rect 40191 14530 40237 14568
rect 40191 14496 40197 14530
rect 40231 14496 40237 14530
rect 40191 14458 40237 14496
rect 40191 14424 40197 14458
rect 40231 14424 40237 14458
rect 40191 14386 40237 14424
rect 40191 14352 40197 14386
rect 40231 14352 40237 14386
rect 40191 14314 40237 14352
rect 40191 14280 40197 14314
rect 40231 14280 40237 14314
rect 40191 14242 40237 14280
rect 40191 14208 40197 14242
rect 40231 14208 40237 14242
rect 40191 14170 40237 14208
rect 40191 14136 40197 14170
rect 40231 14136 40237 14170
rect 40191 14098 40237 14136
rect 40191 14064 40197 14098
rect 40231 14064 40237 14098
rect 40191 14026 40237 14064
rect 40191 13992 40197 14026
rect 40231 13992 40237 14026
rect 40191 13954 40237 13992
rect 40191 13920 40197 13954
rect 40231 13920 40237 13954
rect 40191 13890 40237 13920
rect 40449 15538 40495 15585
rect 40707 15559 40753 15585
rect 41643 15563 41816 15601
rect 40449 15504 40455 15538
rect 40489 15504 40495 15538
rect 40449 15466 40495 15504
rect 40449 15432 40455 15466
rect 40489 15432 40495 15466
rect 40449 15394 40495 15432
rect 40449 15360 40455 15394
rect 40489 15360 40495 15394
rect 40449 15322 40495 15360
rect 40449 15288 40455 15322
rect 40489 15288 40495 15322
rect 40449 15250 40495 15288
rect 40646 15538 40796 15559
rect 40646 15505 40713 15538
rect 40646 15453 40693 15505
rect 40747 15504 40796 15538
rect 40745 15466 40796 15504
rect 40646 15441 40713 15453
rect 40646 15389 40693 15441
rect 40747 15432 40796 15466
rect 40745 15394 40796 15432
rect 40646 15377 40713 15389
rect 40646 15325 40693 15377
rect 40747 15360 40796 15394
rect 40745 15325 40796 15360
rect 40646 15322 40796 15325
rect 40646 15288 40713 15322
rect 40747 15288 40796 15322
rect 40646 15273 40796 15288
rect 41643 15529 41730 15563
rect 41764 15529 41816 15563
rect 41643 15491 41816 15529
rect 41643 15457 41730 15491
rect 41764 15457 41816 15491
rect 41643 15419 41816 15457
rect 41643 15385 41730 15419
rect 41764 15385 41816 15419
rect 41643 15347 41816 15385
rect 41643 15313 41730 15347
rect 41764 15313 41816 15347
rect 41643 15275 41816 15313
rect 40449 15216 40455 15250
rect 40489 15216 40495 15250
rect 40449 15178 40495 15216
rect 40449 15144 40455 15178
rect 40489 15144 40495 15178
rect 40449 15106 40495 15144
rect 40449 15072 40455 15106
rect 40489 15072 40495 15106
rect 40449 15034 40495 15072
rect 40449 15000 40455 15034
rect 40489 15000 40495 15034
rect 40449 14962 40495 15000
rect 40449 14928 40455 14962
rect 40489 14928 40495 14962
rect 40449 14890 40495 14928
rect 40449 14856 40455 14890
rect 40489 14856 40495 14890
rect 40449 14818 40495 14856
rect 40449 14784 40455 14818
rect 40489 14784 40495 14818
rect 40449 14746 40495 14784
rect 40449 14712 40455 14746
rect 40489 14712 40495 14746
rect 40449 14674 40495 14712
rect 40449 14640 40455 14674
rect 40489 14640 40495 14674
rect 40449 14602 40495 14640
rect 40449 14568 40455 14602
rect 40489 14568 40495 14602
rect 40449 14530 40495 14568
rect 40449 14496 40455 14530
rect 40489 14496 40495 14530
rect 40449 14458 40495 14496
rect 40449 14424 40455 14458
rect 40489 14424 40495 14458
rect 40449 14386 40495 14424
rect 40449 14352 40455 14386
rect 40489 14352 40495 14386
rect 40449 14314 40495 14352
rect 40449 14280 40455 14314
rect 40489 14280 40495 14314
rect 40449 14242 40495 14280
rect 40449 14208 40455 14242
rect 40489 14208 40495 14242
rect 40449 14170 40495 14208
rect 40449 14136 40455 14170
rect 40489 14136 40495 14170
rect 40449 14098 40495 14136
rect 40449 14064 40455 14098
rect 40489 14064 40495 14098
rect 40449 14026 40495 14064
rect 40449 13992 40455 14026
rect 40489 13992 40495 14026
rect 40449 13954 40495 13992
rect 40449 13920 40455 13954
rect 40489 13920 40495 13954
rect 39933 13848 39939 13882
rect 39973 13848 39979 13882
rect 39933 13810 39979 13848
rect 39933 13776 39939 13810
rect 39973 13776 39979 13810
rect 39933 13738 39979 13776
rect 39933 13704 39939 13738
rect 39973 13704 39979 13738
rect 39933 13666 39979 13704
rect 39933 13632 39939 13666
rect 39973 13632 39979 13666
rect 39933 13585 39979 13632
rect 40141 13882 40291 13890
rect 40141 13848 40197 13882
rect 40231 13848 40291 13882
rect 40141 13836 40291 13848
rect 40141 13784 40188 13836
rect 40240 13784 40291 13836
rect 40141 13776 40197 13784
rect 40231 13776 40291 13784
rect 40141 13772 40291 13776
rect 40141 13720 40188 13772
rect 40240 13720 40291 13772
rect 40141 13708 40197 13720
rect 40231 13708 40291 13720
rect 40141 13656 40188 13708
rect 40240 13656 40291 13708
rect 40141 13632 40197 13656
rect 40231 13632 40291 13656
rect 40141 13604 40291 13632
rect 40449 13882 40495 13920
rect 40449 13848 40455 13882
rect 40489 13848 40495 13882
rect 40449 13810 40495 13848
rect 40449 13776 40455 13810
rect 40489 13776 40495 13810
rect 40449 13738 40495 13776
rect 40449 13704 40455 13738
rect 40489 13704 40495 13738
rect 40449 13666 40495 13704
rect 40449 13632 40455 13666
rect 40489 13632 40495 13666
rect 40191 13585 40237 13604
rect 40449 13585 40495 13632
rect 40707 15250 40753 15273
rect 40707 15216 40713 15250
rect 40747 15216 40753 15250
rect 40707 15178 40753 15216
rect 41643 15241 41730 15275
rect 41764 15241 41816 15275
rect 41643 15209 41816 15241
rect 40707 15144 40713 15178
rect 40747 15144 40753 15178
rect 40707 15106 40753 15144
rect 40707 15072 40713 15106
rect 40747 15072 40753 15106
rect 40707 15034 40753 15072
rect 40707 15000 40713 15034
rect 40747 15000 40753 15034
rect 40707 14962 40753 15000
rect 40707 14928 40713 14962
rect 40747 14928 40753 14962
rect 40707 14890 40753 14928
rect 40707 14856 40713 14890
rect 40747 14856 40753 14890
rect 40707 14818 40753 14856
rect 40707 14784 40713 14818
rect 40747 14784 40753 14818
rect 40707 14746 40753 14784
rect 40707 14712 40713 14746
rect 40747 14712 40753 14746
rect 40707 14674 40753 14712
rect 40707 14640 40713 14674
rect 40747 14640 40753 14674
rect 40707 14602 40753 14640
rect 40707 14568 40713 14602
rect 40747 14568 40753 14602
rect 40707 14530 40753 14568
rect 40707 14496 40713 14530
rect 40747 14496 40753 14530
rect 40707 14458 40753 14496
rect 40707 14424 40713 14458
rect 40747 14424 40753 14458
rect 40707 14386 40753 14424
rect 40707 14352 40713 14386
rect 40747 14352 40753 14386
rect 40707 14314 40753 14352
rect 40707 14280 40713 14314
rect 40747 14280 40753 14314
rect 40707 14242 40753 14280
rect 40707 14208 40713 14242
rect 40747 14208 40753 14242
rect 40707 14170 40753 14208
rect 40707 14136 40713 14170
rect 40747 14136 40753 14170
rect 40707 14098 40753 14136
rect 40707 14064 40713 14098
rect 40747 14064 40753 14098
rect 40707 14026 40753 14064
rect 40707 13992 40713 14026
rect 40747 13992 40753 14026
rect 40707 13954 40753 13992
rect 40707 13920 40713 13954
rect 40747 13920 40753 13954
rect 40707 13882 40753 13920
rect 40707 13848 40713 13882
rect 40747 13848 40753 13882
rect 40707 13810 40753 13848
rect 40707 13776 40713 13810
rect 40747 13776 40753 13810
rect 40707 13738 40753 13776
rect 40707 13704 40713 13738
rect 40747 13704 40753 13738
rect 40707 13666 40753 13704
rect 40707 13632 40713 13666
rect 40747 13632 40753 13666
rect 40707 13585 40753 13632
rect 41653 13604 41818 13625
rect 37112 13547 37678 13582
rect 37112 13422 37145 13547
rect 23209 13356 24209 13362
rect 24792 13356 24912 13362
rect 23209 13322 23224 13356
rect 23258 13322 23296 13356
rect 23330 13322 23368 13356
rect 23402 13322 23440 13356
rect 23474 13322 23512 13356
rect 23546 13322 23584 13356
rect 23618 13322 23656 13356
rect 23690 13322 23728 13356
rect 23762 13322 23800 13356
rect 23834 13322 23872 13356
rect 23906 13322 23944 13356
rect 23978 13322 24016 13356
rect 24050 13322 24088 13356
rect 24122 13322 24160 13356
rect 24194 13322 24209 13356
rect 23209 13316 24209 13322
rect 24769 13350 25769 13356
rect 24769 13316 24784 13350
rect 24818 13348 24856 13350
rect 24818 13316 24826 13348
rect 24890 13316 24928 13350
rect 24962 13316 25000 13350
rect 25034 13316 25072 13350
rect 25106 13316 25144 13350
rect 25178 13316 25216 13350
rect 25250 13316 25288 13350
rect 25322 13316 25360 13350
rect 25394 13316 25432 13350
rect 25466 13316 25504 13350
rect 25538 13316 25576 13350
rect 25610 13316 25648 13350
rect 25682 13316 25720 13350
rect 25754 13316 25769 13350
rect 24769 13310 24826 13316
rect 23122 13259 23168 13306
rect 23122 13225 23128 13259
rect 23162 13225 23168 13259
rect 23122 13187 23168 13225
rect 23122 13153 23128 13187
rect 23162 13153 23168 13187
rect 23122 13115 23168 13153
rect 23122 13081 23128 13115
rect 23162 13081 23168 13115
rect 23122 13043 23168 13081
rect 23122 13009 23128 13043
rect 23162 13009 23168 13043
rect 23122 12971 23168 13009
rect 23122 12937 23128 12971
rect 23162 12937 23168 12971
rect 23122 12899 23168 12937
rect 23122 12865 23128 12899
rect 23162 12865 23168 12899
rect 23122 12827 23168 12865
rect 23122 12793 23128 12827
rect 23162 12793 23168 12827
rect 23122 12755 23168 12793
rect 23122 12721 23128 12755
rect 23162 12721 23168 12755
rect 23122 12683 23168 12721
rect 23122 12649 23128 12683
rect 23162 12649 23168 12683
rect 23122 12611 23168 12649
rect 23122 12577 23128 12611
rect 23162 12577 23168 12611
rect 23122 12539 23168 12577
rect 23122 12505 23128 12539
rect 23162 12505 23168 12539
rect 23122 12467 23168 12505
rect 23122 12433 23128 12467
rect 23162 12433 23168 12467
rect 23122 12395 23168 12433
rect 23122 12361 23128 12395
rect 23162 12361 23168 12395
rect 23122 12314 23168 12361
rect 24250 13259 24296 13306
rect 24250 13225 24256 13259
rect 24290 13225 24296 13259
rect 24250 13187 24296 13225
rect 24250 13153 24256 13187
rect 24290 13153 24296 13187
rect 24250 13115 24296 13153
rect 24250 13081 24256 13115
rect 24290 13081 24296 13115
rect 24250 13043 24296 13081
rect 24250 13009 24256 13043
rect 24290 13009 24296 13043
rect 24250 12971 24296 13009
rect 24250 12937 24256 12971
rect 24290 12937 24296 12971
rect 24250 12899 24296 12937
rect 24250 12865 24256 12899
rect 24290 12872 24296 12899
rect 24682 13253 24728 13300
rect 24792 13296 24826 13310
rect 24878 13310 25769 13316
rect 26538 13324 26588 13338
rect 24878 13296 24912 13310
rect 24792 13272 24912 13296
rect 24682 13219 24688 13253
rect 24722 13219 24728 13253
rect 24682 13181 24728 13219
rect 24682 13147 24688 13181
rect 24722 13147 24728 13181
rect 24682 13109 24728 13147
rect 24682 13075 24688 13109
rect 24722 13075 24728 13109
rect 24682 13037 24728 13075
rect 24682 13003 24688 13037
rect 24722 13003 24728 13037
rect 24682 12965 24728 13003
rect 24682 12931 24688 12965
rect 24722 12931 24728 12965
rect 24682 12893 24728 12931
rect 24682 12872 24688 12893
rect 24290 12865 24688 12872
rect 24250 12859 24688 12865
rect 24722 12859 24728 12893
rect 24250 12827 24728 12859
rect 24250 12793 24256 12827
rect 24290 12821 24728 12827
rect 24290 12793 24688 12821
rect 24250 12787 24688 12793
rect 24722 12787 24728 12821
rect 24250 12755 24728 12787
rect 24250 12721 24256 12755
rect 24290 12749 24728 12755
rect 24290 12721 24688 12749
rect 24250 12715 24688 12721
rect 24722 12715 24728 12749
rect 24250 12683 24728 12715
rect 24250 12649 24256 12683
rect 24290 12677 24728 12683
rect 24290 12649 24688 12677
rect 24250 12643 24688 12649
rect 24722 12643 24728 12677
rect 24250 12642 24728 12643
rect 24250 12611 24296 12642
rect 24250 12577 24256 12611
rect 24290 12577 24296 12611
rect 24250 12539 24296 12577
rect 24250 12505 24256 12539
rect 24290 12505 24296 12539
rect 24250 12467 24296 12505
rect 24250 12433 24256 12467
rect 24290 12433 24296 12467
rect 24250 12395 24296 12433
rect 24250 12361 24256 12395
rect 24290 12361 24296 12395
rect 24682 12605 24728 12642
rect 24682 12571 24688 12605
rect 24722 12571 24728 12605
rect 24682 12533 24728 12571
rect 24682 12499 24688 12533
rect 24722 12499 24728 12533
rect 24682 12461 24728 12499
rect 24682 12427 24688 12461
rect 24722 12427 24728 12461
rect 24682 12389 24728 12427
rect 24682 12382 24688 12389
rect 23209 12298 24209 12304
rect 24250 12298 24296 12361
rect 23209 12264 23224 12298
rect 23258 12264 23296 12298
rect 23330 12264 23368 12298
rect 23402 12264 23440 12298
rect 23474 12264 23512 12298
rect 23546 12264 23584 12298
rect 23618 12264 23656 12298
rect 23690 12264 23728 12298
rect 23762 12264 23800 12298
rect 23834 12264 23872 12298
rect 23906 12264 23944 12298
rect 23978 12264 24016 12298
rect 24050 12264 24088 12298
rect 24122 12264 24160 12298
rect 24194 12264 24296 12298
rect 24652 12355 24688 12382
rect 24722 12355 24728 12389
rect 24652 12308 24728 12355
rect 25810 13253 25856 13300
rect 25810 13219 25816 13253
rect 25850 13219 25856 13253
rect 25810 13181 25856 13219
rect 25810 13147 25816 13181
rect 25850 13147 25856 13181
rect 25810 13109 25856 13147
rect 25810 13075 25816 13109
rect 25850 13075 25856 13109
rect 25810 13037 25856 13075
rect 25810 13003 25816 13037
rect 25850 13003 25856 13037
rect 25810 12965 25856 13003
rect 25810 12931 25816 12965
rect 25850 12931 25856 12965
rect 25810 12893 25856 12931
rect 26538 13290 26546 13324
rect 26580 13290 26588 13324
rect 26856 13324 26906 13338
rect 26856 13322 26864 13324
rect 26538 13252 26588 13290
rect 26538 13218 26546 13252
rect 26580 13218 26588 13252
rect 26538 13180 26588 13218
rect 26538 13146 26546 13180
rect 26580 13146 26588 13180
rect 26538 13108 26588 13146
rect 26538 13074 26546 13108
rect 26580 13074 26588 13108
rect 26538 13036 26588 13074
rect 26538 13002 26546 13036
rect 26580 13002 26588 13036
rect 26538 12964 26588 13002
rect 26538 12930 26546 12964
rect 26580 12930 26588 12964
rect 26538 12917 26588 12930
rect 26672 13298 26864 13322
rect 26898 13322 26906 13324
rect 27174 13324 27224 13338
rect 26672 12926 26697 13298
rect 26898 13290 26912 13322
rect 26877 13252 26912 13290
rect 26898 13218 26912 13252
rect 26877 13180 26912 13218
rect 26898 13146 26912 13180
rect 26877 13108 26912 13146
rect 26898 13074 26912 13108
rect 26877 13036 26912 13074
rect 26898 13002 26912 13036
rect 26877 12964 26912 13002
rect 26898 12930 26912 12964
rect 26877 12926 26912 12930
rect 26672 12902 26912 12926
rect 27174 13290 27182 13324
rect 27216 13290 27224 13324
rect 27174 13252 27224 13290
rect 27174 13218 27182 13252
rect 27216 13218 27224 13252
rect 27174 13180 27224 13218
rect 27174 13146 27182 13180
rect 27216 13146 27224 13180
rect 27174 13108 27224 13146
rect 27174 13074 27182 13108
rect 27216 13074 27224 13108
rect 27174 13036 27224 13074
rect 27174 13002 27182 13036
rect 27216 13002 27224 13036
rect 27174 12964 27224 13002
rect 27174 12930 27182 12964
rect 27216 12930 27224 12964
rect 27174 12917 27224 12930
rect 27710 13308 27760 13322
rect 27710 13274 27718 13308
rect 27752 13274 27760 13308
rect 27710 13236 27760 13274
rect 27710 13202 27718 13236
rect 27752 13202 27760 13236
rect 27710 13164 27760 13202
rect 27710 13130 27718 13164
rect 27752 13130 27760 13164
rect 27710 13092 27760 13130
rect 27710 13058 27718 13092
rect 27752 13058 27760 13092
rect 27710 13020 27760 13058
rect 27710 12986 27718 13020
rect 27752 12986 27760 13020
rect 27710 12948 27760 12986
rect 27710 12914 27718 12948
rect 27752 12914 27760 12948
rect 27710 12901 27760 12914
rect 28024 13308 28414 13332
rect 28024 13274 28036 13308
rect 28070 13274 28354 13308
rect 28388 13274 28414 13308
rect 28024 13236 28414 13274
rect 28024 13202 28036 13236
rect 28070 13202 28354 13236
rect 28388 13202 28414 13236
rect 28024 13164 28414 13202
rect 28024 13130 28036 13164
rect 28070 13130 28354 13164
rect 28388 13130 28414 13164
rect 28024 13092 28414 13130
rect 28024 13058 28036 13092
rect 28070 13058 28354 13092
rect 28388 13058 28414 13092
rect 28024 13020 28414 13058
rect 28024 12986 28036 13020
rect 28070 12986 28354 13020
rect 28388 12986 28414 13020
rect 28024 12948 28414 12986
rect 28024 12914 28036 12948
rect 28070 12914 28354 12948
rect 28388 12914 28414 12948
rect 28024 12902 28414 12914
rect 28660 13308 29050 13332
rect 28660 13274 28672 13308
rect 28706 13274 28990 13308
rect 29024 13274 29050 13308
rect 28660 13236 29050 13274
rect 28660 13202 28672 13236
rect 28706 13202 28990 13236
rect 29024 13202 29050 13236
rect 28660 13164 29050 13202
rect 28660 13130 28672 13164
rect 28706 13130 28990 13164
rect 29024 13130 29050 13164
rect 28660 13092 29050 13130
rect 28660 13058 28672 13092
rect 28706 13058 28990 13092
rect 29024 13058 29050 13092
rect 28660 13020 29050 13058
rect 28660 12986 28672 13020
rect 28706 12986 28990 13020
rect 29024 12986 29050 13020
rect 28660 12948 29050 12986
rect 28660 12914 28672 12948
rect 28706 12914 28990 12948
rect 29024 12914 29050 12948
rect 28660 12902 29050 12914
rect 29200 13308 29466 13407
rect 29200 13274 29308 13308
rect 29342 13274 29466 13308
rect 29200 13236 29466 13274
rect 29200 13202 29308 13236
rect 29342 13202 29466 13236
rect 29200 13164 29466 13202
rect 29200 13130 29308 13164
rect 29342 13130 29466 13164
rect 29200 13092 29466 13130
rect 29200 13058 29308 13092
rect 29342 13058 29466 13092
rect 29200 13020 29466 13058
rect 29200 12986 29308 13020
rect 29342 12986 29466 13020
rect 29200 12948 29466 12986
rect 29200 12914 29308 12948
rect 29342 12914 29466 12948
rect 28028 12901 28078 12902
rect 28346 12901 28396 12902
rect 28664 12901 28714 12902
rect 28982 12901 29032 12902
rect 29200 12894 29466 12914
rect 29618 13308 29668 13322
rect 29618 13274 29626 13308
rect 29660 13274 29668 13308
rect 29618 13236 29668 13274
rect 29618 13202 29626 13236
rect 29660 13202 29668 13236
rect 29618 13164 29668 13202
rect 29618 13130 29626 13164
rect 29660 13130 29668 13164
rect 37111 13175 37145 13422
rect 37645 13422 37678 13547
rect 41653 13571 41730 13604
rect 41764 13571 41818 13604
rect 38720 13517 38894 13537
rect 38720 13465 38747 13517
rect 38799 13465 38811 13517
rect 38863 13465 38894 13517
rect 38720 13451 38894 13465
rect 37645 13320 40431 13422
rect 37645 13312 40330 13320
rect 37645 13310 39282 13312
rect 37645 13302 39042 13310
rect 37645 13268 38253 13302
rect 38287 13276 39042 13302
rect 39076 13278 39282 13310
rect 39316 13307 40330 13312
rect 39316 13278 40061 13307
rect 39076 13276 40061 13278
rect 38287 13273 40061 13276
rect 40095 13286 40330 13307
rect 40364 13286 40431 13320
rect 40095 13273 40431 13286
rect 38287 13268 40431 13273
rect 37645 13248 40431 13268
rect 37645 13240 40330 13248
rect 37645 13238 39282 13240
rect 37645 13230 39042 13238
rect 37645 13196 38253 13230
rect 38287 13204 39042 13230
rect 39076 13206 39282 13238
rect 39316 13235 40330 13240
rect 39316 13206 40061 13235
rect 39076 13204 40061 13206
rect 38287 13201 40061 13204
rect 40095 13214 40330 13235
rect 40364 13214 40431 13248
rect 40095 13201 40431 13214
rect 38287 13196 40431 13201
rect 37645 13175 40431 13196
rect 37111 13152 40431 13175
rect 41653 13199 41674 13571
rect 41790 13199 41818 13571
rect 41653 13154 41818 13199
rect 37112 13142 37678 13152
rect 29618 13092 29668 13130
rect 29618 13058 29626 13092
rect 29660 13058 29668 13092
rect 29618 13020 29668 13058
rect 29618 12986 29626 13020
rect 29660 12986 29668 13020
rect 29618 12948 29668 12986
rect 29618 12914 29626 12948
rect 29660 12914 29668 12948
rect 29618 12901 29668 12914
rect 25810 12859 25816 12893
rect 25850 12859 25856 12893
rect 25810 12821 25856 12859
rect 25810 12787 25816 12821
rect 25850 12787 25856 12821
rect 25810 12749 25856 12787
rect 25810 12715 25816 12749
rect 25850 12715 25856 12749
rect 25810 12677 25856 12715
rect 25810 12643 25816 12677
rect 25850 12643 25856 12677
rect 25810 12605 25856 12643
rect 25810 12571 25816 12605
rect 25850 12571 25856 12605
rect 25810 12533 25856 12571
rect 25810 12499 25816 12533
rect 25850 12499 25856 12533
rect 25810 12461 25856 12499
rect 25810 12427 25816 12461
rect 25850 12427 25856 12461
rect 25810 12389 25856 12427
rect 25810 12355 25816 12389
rect 25850 12355 25856 12389
rect 23209 12258 24209 12264
rect 23222 11822 23432 12258
rect 24652 12242 24682 12308
rect 25632 12298 25762 12312
rect 25810 12308 25856 12355
rect 24769 12292 25666 12298
rect 25718 12292 25769 12298
rect 24769 12258 24784 12292
rect 24818 12258 24856 12292
rect 24890 12258 24928 12292
rect 24962 12258 25000 12292
rect 25034 12258 25072 12292
rect 25106 12258 25144 12292
rect 25178 12258 25216 12292
rect 25250 12258 25288 12292
rect 25322 12258 25360 12292
rect 25394 12258 25432 12292
rect 25466 12258 25504 12292
rect 25538 12258 25576 12292
rect 25610 12258 25648 12292
rect 25718 12258 25720 12292
rect 25754 12258 25769 12292
rect 24769 12252 25666 12258
rect 25632 12246 25666 12252
rect 25718 12252 25769 12258
rect 25718 12246 25762 12252
rect 24652 12195 24728 12242
rect 25632 12232 25762 12246
rect 24652 12192 24688 12195
rect 24682 12161 24688 12192
rect 24722 12161 24728 12195
rect 24682 12123 24728 12161
rect 24682 12089 24688 12123
rect 24722 12089 24728 12123
rect 24682 12051 24728 12089
rect 24682 12017 24688 12051
rect 24722 12017 24728 12051
rect 24682 11979 24728 12017
rect 24682 11945 24688 11979
rect 24722 11945 24728 11979
rect 24682 11907 24728 11945
rect 24682 11873 24688 11907
rect 24722 11873 24728 11907
rect 24682 11835 24728 11873
rect 23130 11816 24130 11822
rect 23130 11782 23145 11816
rect 23179 11782 23217 11816
rect 23251 11782 23289 11816
rect 23323 11782 23361 11816
rect 23395 11782 23433 11816
rect 23467 11782 23505 11816
rect 23539 11782 23577 11816
rect 23611 11782 23649 11816
rect 23683 11782 23721 11816
rect 23755 11782 23793 11816
rect 23827 11782 23865 11816
rect 23899 11782 23937 11816
rect 23971 11782 24009 11816
rect 24043 11782 24081 11816
rect 24115 11782 24130 11816
rect 23130 11776 24130 11782
rect 24682 11801 24688 11835
rect 24722 11801 24728 11835
rect 23052 11719 23098 11766
rect 23052 11685 23058 11719
rect 23092 11685 23098 11719
rect 23052 11647 23098 11685
rect 23052 11613 23058 11647
rect 23092 11613 23098 11647
rect 23052 11575 23098 11613
rect 23052 11541 23058 11575
rect 23092 11541 23098 11575
rect 23052 11503 23098 11541
rect 23052 11469 23058 11503
rect 23092 11469 23098 11503
rect 23052 11431 23098 11469
rect 23052 11397 23058 11431
rect 23092 11397 23098 11431
rect 23052 11359 23098 11397
rect 23052 11325 23058 11359
rect 23092 11325 23098 11359
rect 23052 11287 23098 11325
rect 23052 11253 23058 11287
rect 23092 11253 23098 11287
rect 23052 11215 23098 11253
rect 23052 11181 23058 11215
rect 23092 11181 23098 11215
rect 23052 11143 23098 11181
rect 23052 11109 23058 11143
rect 23092 11109 23098 11143
rect 23052 11092 23098 11109
rect 22632 11071 23098 11092
rect 22632 11037 23058 11071
rect 23092 11037 23098 11071
rect 22632 10999 23098 11037
rect 22632 10965 23058 10999
rect 23092 10965 23098 10999
rect 22632 10927 23098 10965
rect 22632 10893 23058 10927
rect 23092 10893 23098 10927
rect 22632 10855 23098 10893
rect 22632 10821 23058 10855
rect 23092 10821 23098 10855
rect 22632 10774 23098 10821
rect 24162 11719 24208 11766
rect 24162 11685 24168 11719
rect 24202 11685 24208 11719
rect 24162 11647 24208 11685
rect 24162 11613 24168 11647
rect 24202 11613 24208 11647
rect 24162 11575 24208 11613
rect 24162 11541 24168 11575
rect 24202 11541 24208 11575
rect 24162 11503 24208 11541
rect 24162 11469 24168 11503
rect 24202 11469 24208 11503
rect 24162 11431 24208 11469
rect 24162 11397 24168 11431
rect 24202 11397 24208 11431
rect 24162 11359 24208 11397
rect 24162 11325 24168 11359
rect 24202 11325 24208 11359
rect 24162 11287 24208 11325
rect 24682 11763 24728 11801
rect 24682 11729 24688 11763
rect 24722 11729 24728 11763
rect 24682 11691 24728 11729
rect 24682 11657 24688 11691
rect 24722 11657 24728 11691
rect 24682 11619 24728 11657
rect 24682 11585 24688 11619
rect 24722 11585 24728 11619
rect 24682 11547 24728 11585
rect 24682 11513 24688 11547
rect 24722 11513 24728 11547
rect 24682 11475 24728 11513
rect 24682 11441 24688 11475
rect 24722 11441 24728 11475
rect 24682 11403 24728 11441
rect 24682 11369 24688 11403
rect 24722 11369 24728 11403
rect 24682 11331 24728 11369
rect 24682 11312 24688 11331
rect 24162 11253 24168 11287
rect 24202 11253 24208 11287
rect 24162 11215 24208 11253
rect 24162 11181 24168 11215
rect 24202 11181 24208 11215
rect 24162 11143 24208 11181
rect 24162 11109 24168 11143
rect 24202 11109 24208 11143
rect 24652 11297 24688 11312
rect 24722 11297 24728 11331
rect 24652 11250 24728 11297
rect 25810 12195 25856 12242
rect 25810 12161 25816 12195
rect 25850 12161 25856 12195
rect 25810 12123 25856 12161
rect 25810 12089 25816 12123
rect 25850 12089 25856 12123
rect 25810 12051 25856 12089
rect 25810 12017 25816 12051
rect 25850 12017 25856 12051
rect 25810 11979 25856 12017
rect 25810 11945 25816 11979
rect 25850 11945 25856 11979
rect 36827 11992 41925 12052
rect 36827 11986 37019 11992
rect 36827 11952 36870 11986
rect 36904 11952 36942 11986
rect 36976 11952 37019 11986
rect 36827 11946 37019 11952
rect 37085 11986 37277 11992
rect 37085 11952 37128 11986
rect 37162 11952 37200 11986
rect 37234 11952 37277 11986
rect 37085 11946 37277 11952
rect 37343 11986 37535 11992
rect 37343 11952 37386 11986
rect 37420 11952 37458 11986
rect 37492 11952 37535 11986
rect 37343 11946 37535 11952
rect 37601 11986 37793 11992
rect 37601 11952 37644 11986
rect 37678 11952 37716 11986
rect 37750 11952 37793 11986
rect 37601 11946 37793 11952
rect 37859 11986 38051 11992
rect 37859 11952 37902 11986
rect 37936 11952 37974 11986
rect 38008 11952 38051 11986
rect 37859 11946 38051 11952
rect 38117 11986 38309 11992
rect 38117 11952 38160 11986
rect 38194 11952 38232 11986
rect 38266 11952 38309 11986
rect 38117 11946 38309 11952
rect 38375 11986 38567 11992
rect 38375 11952 38418 11986
rect 38452 11952 38490 11986
rect 38524 11952 38567 11986
rect 38375 11946 38567 11952
rect 38633 11986 38825 11992
rect 38633 11952 38676 11986
rect 38710 11952 38748 11986
rect 38782 11952 38825 11986
rect 38633 11946 38825 11952
rect 38891 11986 39083 11992
rect 38891 11952 38934 11986
rect 38968 11952 39006 11986
rect 39040 11952 39083 11986
rect 38891 11946 39083 11952
rect 39149 11986 39341 11992
rect 39149 11952 39192 11986
rect 39226 11952 39264 11986
rect 39298 11952 39341 11986
rect 39149 11946 39341 11952
rect 39407 11986 39599 11992
rect 39407 11952 39450 11986
rect 39484 11952 39522 11986
rect 39556 11952 39599 11986
rect 39407 11946 39599 11952
rect 39665 11986 39857 11992
rect 39665 11952 39708 11986
rect 39742 11952 39780 11986
rect 39814 11952 39857 11986
rect 39665 11946 39857 11952
rect 39923 11986 40115 11992
rect 39923 11952 39966 11986
rect 40000 11952 40038 11986
rect 40072 11952 40115 11986
rect 39923 11946 40115 11952
rect 40181 11986 40373 11992
rect 40181 11952 40224 11986
rect 40258 11952 40296 11986
rect 40330 11952 40373 11986
rect 40181 11946 40373 11952
rect 40439 11986 40631 11992
rect 40439 11952 40482 11986
rect 40516 11952 40554 11986
rect 40588 11952 40631 11986
rect 40439 11946 40631 11952
rect 40697 11986 40889 11992
rect 40697 11952 40740 11986
rect 40774 11952 40812 11986
rect 40846 11952 40889 11986
rect 40697 11946 40889 11952
rect 40955 11986 41147 11992
rect 40955 11952 40998 11986
rect 41032 11952 41070 11986
rect 41104 11952 41147 11986
rect 40955 11946 41147 11952
rect 41213 11986 41405 11992
rect 41213 11952 41256 11986
rect 41290 11952 41328 11986
rect 41362 11952 41405 11986
rect 41213 11946 41405 11952
rect 41471 11986 41663 11992
rect 41471 11952 41514 11986
rect 41548 11952 41586 11986
rect 41620 11952 41663 11986
rect 41471 11946 41663 11952
rect 41729 11986 41921 11992
rect 41729 11952 41772 11986
rect 41806 11952 41844 11986
rect 41878 11952 41921 11986
rect 41729 11946 41921 11952
rect 25810 11907 25856 11945
rect 25810 11873 25816 11907
rect 25850 11873 25856 11907
rect 25810 11835 25856 11873
rect 25810 11801 25816 11835
rect 25850 11801 25856 11835
rect 25810 11763 25856 11801
rect 25810 11729 25816 11763
rect 25850 11729 25856 11763
rect 25810 11691 25856 11729
rect 25810 11657 25816 11691
rect 25850 11657 25856 11691
rect 25810 11619 25856 11657
rect 25810 11585 25816 11619
rect 25850 11585 25856 11619
rect 25810 11547 25856 11585
rect 25810 11513 25816 11547
rect 25850 11513 25856 11547
rect 25810 11475 25856 11513
rect 25810 11441 25816 11475
rect 25850 11441 25856 11475
rect 25810 11403 25856 11441
rect 25810 11369 25816 11403
rect 25850 11369 25856 11403
rect 25810 11331 25856 11369
rect 25810 11297 25816 11331
rect 25850 11297 25856 11331
rect 24652 11184 24682 11250
rect 24792 11243 24912 11282
rect 25810 11250 25856 11297
rect 36771 11899 36817 11914
rect 36771 11865 36777 11899
rect 36811 11865 36817 11899
rect 36771 11827 36817 11865
rect 36771 11793 36777 11827
rect 36811 11793 36817 11827
rect 36771 11755 36817 11793
rect 36771 11721 36777 11755
rect 36811 11721 36817 11755
rect 36771 11683 36817 11721
rect 36771 11649 36777 11683
rect 36811 11649 36817 11683
rect 36771 11611 36817 11649
rect 36771 11577 36777 11611
rect 36811 11577 36817 11611
rect 36771 11539 36817 11577
rect 36771 11505 36777 11539
rect 36811 11505 36817 11539
rect 37029 11899 37075 11914
rect 37029 11865 37035 11899
rect 37069 11865 37075 11899
rect 37029 11827 37075 11865
rect 37029 11793 37035 11827
rect 37069 11793 37075 11827
rect 37029 11755 37075 11793
rect 37029 11721 37035 11755
rect 37069 11721 37075 11755
rect 37029 11683 37075 11721
rect 37029 11649 37035 11683
rect 37069 11649 37075 11683
rect 37029 11611 37075 11649
rect 37029 11577 37035 11611
rect 37069 11577 37075 11611
rect 37029 11539 37075 11577
rect 37029 11523 37035 11539
rect 36771 11467 36817 11505
rect 36771 11433 36777 11467
rect 36811 11433 36817 11467
rect 36771 11395 36817 11433
rect 36771 11361 36777 11395
rect 36811 11361 36817 11395
rect 37007 11516 37035 11523
rect 37069 11523 37075 11539
rect 37287 11899 37333 11914
rect 37287 11865 37293 11899
rect 37327 11865 37333 11899
rect 37287 11827 37333 11865
rect 37287 11793 37293 11827
rect 37327 11793 37333 11827
rect 37287 11755 37333 11793
rect 37287 11721 37293 11755
rect 37327 11721 37333 11755
rect 37287 11683 37333 11721
rect 37287 11649 37293 11683
rect 37327 11649 37333 11683
rect 37287 11611 37333 11649
rect 37287 11577 37293 11611
rect 37327 11577 37333 11611
rect 37287 11539 37333 11577
rect 37069 11516 37096 11523
rect 37007 11464 37026 11516
rect 37078 11464 37096 11516
rect 37007 11452 37035 11464
rect 37069 11452 37096 11464
rect 37007 11400 37026 11452
rect 37078 11400 37096 11452
rect 37007 11395 37096 11400
rect 37007 11390 37035 11395
rect 36771 11323 36817 11361
rect 36771 11289 36777 11323
rect 36811 11289 36817 11323
rect 36771 11251 36817 11289
rect 37029 11361 37035 11390
rect 37069 11390 37096 11395
rect 37287 11505 37293 11539
rect 37327 11505 37333 11539
rect 37545 11899 37591 11914
rect 37545 11865 37551 11899
rect 37585 11865 37591 11899
rect 37545 11827 37591 11865
rect 37545 11793 37551 11827
rect 37585 11793 37591 11827
rect 37545 11755 37591 11793
rect 37545 11721 37551 11755
rect 37585 11721 37591 11755
rect 37545 11683 37591 11721
rect 37545 11649 37551 11683
rect 37585 11649 37591 11683
rect 37545 11611 37591 11649
rect 37545 11577 37551 11611
rect 37585 11577 37591 11611
rect 37545 11539 37591 11577
rect 37545 11523 37551 11539
rect 37287 11467 37333 11505
rect 37287 11433 37293 11467
rect 37327 11433 37333 11467
rect 37287 11395 37333 11433
rect 37069 11361 37075 11390
rect 37029 11323 37075 11361
rect 37029 11289 37035 11323
rect 37069 11289 37075 11323
rect 37029 11251 37075 11289
rect 37287 11361 37293 11395
rect 37327 11361 37333 11395
rect 37525 11505 37551 11523
rect 37585 11523 37591 11539
rect 37803 11899 37849 11914
rect 37803 11865 37809 11899
rect 37843 11865 37849 11899
rect 37803 11827 37849 11865
rect 37803 11793 37809 11827
rect 37843 11793 37849 11827
rect 37803 11755 37849 11793
rect 37803 11721 37809 11755
rect 37843 11721 37849 11755
rect 37803 11683 37849 11721
rect 37803 11649 37809 11683
rect 37843 11649 37849 11683
rect 37803 11611 37849 11649
rect 37803 11577 37809 11611
rect 37843 11577 37849 11611
rect 37803 11539 37849 11577
rect 37585 11505 37611 11523
rect 37525 11483 37611 11505
rect 37525 11431 37541 11483
rect 37593 11431 37611 11483
rect 37525 11395 37611 11431
rect 37525 11390 37551 11395
rect 37287 11323 37333 11361
rect 37287 11289 37293 11323
rect 37327 11289 37333 11323
rect 37287 11251 37333 11289
rect 37545 11361 37551 11390
rect 37585 11390 37611 11395
rect 37803 11505 37809 11539
rect 37843 11505 37849 11539
rect 38061 11899 38107 11914
rect 38061 11865 38067 11899
rect 38101 11865 38107 11899
rect 38061 11827 38107 11865
rect 38061 11793 38067 11827
rect 38101 11793 38107 11827
rect 38061 11755 38107 11793
rect 38061 11721 38067 11755
rect 38101 11721 38107 11755
rect 38061 11683 38107 11721
rect 38061 11649 38067 11683
rect 38101 11649 38107 11683
rect 38061 11611 38107 11649
rect 38061 11577 38067 11611
rect 38101 11577 38107 11611
rect 38061 11539 38107 11577
rect 38061 11523 38067 11539
rect 37803 11467 37849 11505
rect 37803 11433 37809 11467
rect 37843 11433 37849 11467
rect 37803 11395 37849 11433
rect 37585 11361 37591 11390
rect 37545 11323 37591 11361
rect 37545 11289 37551 11323
rect 37585 11289 37591 11323
rect 37545 11251 37591 11289
rect 37803 11361 37809 11395
rect 37843 11361 37849 11395
rect 38043 11505 38067 11523
rect 38101 11523 38107 11539
rect 38319 11899 38365 11914
rect 38319 11865 38325 11899
rect 38359 11865 38365 11899
rect 38319 11827 38365 11865
rect 38319 11793 38325 11827
rect 38359 11793 38365 11827
rect 38319 11755 38365 11793
rect 38319 11721 38325 11755
rect 38359 11721 38365 11755
rect 38319 11683 38365 11721
rect 38319 11649 38325 11683
rect 38359 11649 38365 11683
rect 38319 11611 38365 11649
rect 38319 11577 38325 11611
rect 38359 11577 38365 11611
rect 38319 11539 38365 11577
rect 38101 11505 38126 11523
rect 38043 11482 38126 11505
rect 38043 11430 38058 11482
rect 38110 11430 38126 11482
rect 38043 11395 38126 11430
rect 38043 11390 38067 11395
rect 37803 11323 37849 11361
rect 37803 11289 37809 11323
rect 37843 11289 37849 11323
rect 37803 11251 37849 11289
rect 38061 11361 38067 11390
rect 38101 11390 38126 11395
rect 38319 11505 38325 11539
rect 38359 11505 38365 11539
rect 38577 11899 38623 11914
rect 38577 11865 38583 11899
rect 38617 11865 38623 11899
rect 38577 11827 38623 11865
rect 38577 11793 38583 11827
rect 38617 11793 38623 11827
rect 38577 11755 38623 11793
rect 38577 11721 38583 11755
rect 38617 11721 38623 11755
rect 38577 11683 38623 11721
rect 38577 11649 38583 11683
rect 38617 11649 38623 11683
rect 38577 11611 38623 11649
rect 38577 11577 38583 11611
rect 38617 11577 38623 11611
rect 38577 11539 38623 11577
rect 38577 11523 38583 11539
rect 38319 11467 38365 11505
rect 38319 11433 38325 11467
rect 38359 11433 38365 11467
rect 38319 11395 38365 11433
rect 38101 11361 38107 11390
rect 38061 11323 38107 11361
rect 38061 11289 38067 11323
rect 38101 11289 38107 11323
rect 38061 11251 38107 11289
rect 38319 11361 38325 11395
rect 38359 11361 38365 11395
rect 38558 11505 38583 11523
rect 38617 11523 38623 11539
rect 38835 11899 38881 11914
rect 38835 11865 38841 11899
rect 38875 11865 38881 11899
rect 38835 11827 38881 11865
rect 38835 11793 38841 11827
rect 38875 11793 38881 11827
rect 38835 11755 38881 11793
rect 38835 11721 38841 11755
rect 38875 11721 38881 11755
rect 38835 11683 38881 11721
rect 38835 11649 38841 11683
rect 38875 11649 38881 11683
rect 38835 11611 38881 11649
rect 38835 11577 38841 11611
rect 38875 11577 38881 11611
rect 38835 11539 38881 11577
rect 38617 11505 38643 11523
rect 38558 11483 38643 11505
rect 38558 11431 38574 11483
rect 38626 11431 38643 11483
rect 38558 11395 38643 11431
rect 38558 11390 38583 11395
rect 38319 11323 38365 11361
rect 38319 11289 38325 11323
rect 38359 11289 38365 11323
rect 38319 11251 38365 11289
rect 38577 11361 38583 11390
rect 38617 11390 38643 11395
rect 38835 11505 38841 11539
rect 38875 11505 38881 11539
rect 39093 11899 39139 11914
rect 39093 11865 39099 11899
rect 39133 11865 39139 11899
rect 39093 11827 39139 11865
rect 39093 11793 39099 11827
rect 39133 11793 39139 11827
rect 39093 11755 39139 11793
rect 39093 11721 39099 11755
rect 39133 11721 39139 11755
rect 39093 11683 39139 11721
rect 39093 11649 39099 11683
rect 39133 11649 39139 11683
rect 39093 11611 39139 11649
rect 39093 11577 39099 11611
rect 39133 11577 39139 11611
rect 39093 11539 39139 11577
rect 39093 11523 39099 11539
rect 38835 11467 38881 11505
rect 38835 11433 38841 11467
rect 38875 11433 38881 11467
rect 38835 11395 38881 11433
rect 38617 11361 38623 11390
rect 38577 11323 38623 11361
rect 38577 11289 38583 11323
rect 38617 11289 38623 11323
rect 38577 11251 38623 11289
rect 38835 11361 38841 11395
rect 38875 11361 38881 11395
rect 39074 11505 39099 11523
rect 39133 11523 39139 11539
rect 39351 11899 39397 11914
rect 39351 11865 39357 11899
rect 39391 11865 39397 11899
rect 39351 11827 39397 11865
rect 39351 11793 39357 11827
rect 39391 11793 39397 11827
rect 39351 11755 39397 11793
rect 39351 11721 39357 11755
rect 39391 11721 39397 11755
rect 39351 11683 39397 11721
rect 39351 11649 39357 11683
rect 39391 11649 39397 11683
rect 39351 11611 39397 11649
rect 39351 11577 39357 11611
rect 39391 11577 39397 11611
rect 39351 11539 39397 11577
rect 39133 11505 39160 11523
rect 39074 11481 39160 11505
rect 39074 11429 39090 11481
rect 39142 11429 39160 11481
rect 39074 11395 39160 11429
rect 39074 11390 39099 11395
rect 38835 11323 38881 11361
rect 38835 11289 38841 11323
rect 38875 11289 38881 11323
rect 38835 11251 38881 11289
rect 39093 11361 39099 11390
rect 39133 11390 39160 11395
rect 39351 11505 39357 11539
rect 39391 11505 39397 11539
rect 39609 11899 39655 11914
rect 39609 11865 39615 11899
rect 39649 11865 39655 11899
rect 39609 11827 39655 11865
rect 39609 11793 39615 11827
rect 39649 11793 39655 11827
rect 39609 11755 39655 11793
rect 39609 11721 39615 11755
rect 39649 11721 39655 11755
rect 39609 11683 39655 11721
rect 39609 11649 39615 11683
rect 39649 11649 39655 11683
rect 39609 11611 39655 11649
rect 39609 11577 39615 11611
rect 39649 11577 39655 11611
rect 39609 11539 39655 11577
rect 39609 11523 39615 11539
rect 39351 11467 39397 11505
rect 39351 11433 39357 11467
rect 39391 11433 39397 11467
rect 39351 11395 39397 11433
rect 39133 11361 39139 11390
rect 39093 11323 39139 11361
rect 39093 11289 39099 11323
rect 39133 11289 39139 11323
rect 39093 11251 39139 11289
rect 39351 11361 39357 11395
rect 39391 11361 39397 11395
rect 39592 11505 39615 11523
rect 39649 11523 39655 11539
rect 39867 11899 39913 11914
rect 39867 11865 39873 11899
rect 39907 11865 39913 11899
rect 39867 11827 39913 11865
rect 39867 11793 39873 11827
rect 39907 11793 39913 11827
rect 39867 11755 39913 11793
rect 39867 11721 39873 11755
rect 39907 11721 39913 11755
rect 39867 11683 39913 11721
rect 39867 11649 39873 11683
rect 39907 11649 39913 11683
rect 39867 11611 39913 11649
rect 39867 11577 39873 11611
rect 39907 11577 39913 11611
rect 39867 11539 39913 11577
rect 39649 11505 39672 11523
rect 39592 11482 39672 11505
rect 39592 11430 39606 11482
rect 39658 11430 39672 11482
rect 39592 11395 39672 11430
rect 39592 11390 39615 11395
rect 39351 11323 39397 11361
rect 39351 11289 39357 11323
rect 39391 11289 39397 11323
rect 39351 11251 39397 11289
rect 39609 11361 39615 11390
rect 39649 11390 39672 11395
rect 39867 11505 39873 11539
rect 39907 11505 39913 11539
rect 40125 11899 40171 11914
rect 40125 11865 40131 11899
rect 40165 11865 40171 11899
rect 40125 11827 40171 11865
rect 40125 11793 40131 11827
rect 40165 11793 40171 11827
rect 40125 11755 40171 11793
rect 40125 11721 40131 11755
rect 40165 11721 40171 11755
rect 40125 11683 40171 11721
rect 40125 11649 40131 11683
rect 40165 11649 40171 11683
rect 40125 11611 40171 11649
rect 40125 11577 40131 11611
rect 40165 11577 40171 11611
rect 40125 11539 40171 11577
rect 40125 11523 40131 11539
rect 39867 11467 39913 11505
rect 39867 11433 39873 11467
rect 39907 11433 39913 11467
rect 39867 11395 39913 11433
rect 39649 11361 39655 11390
rect 39609 11323 39655 11361
rect 39609 11289 39615 11323
rect 39649 11289 39655 11323
rect 39609 11251 39655 11289
rect 39867 11361 39873 11395
rect 39907 11361 39913 11395
rect 40108 11505 40131 11523
rect 40165 11523 40171 11539
rect 40383 11899 40429 11914
rect 40383 11865 40389 11899
rect 40423 11865 40429 11899
rect 40383 11827 40429 11865
rect 40383 11793 40389 11827
rect 40423 11793 40429 11827
rect 40383 11755 40429 11793
rect 40383 11721 40389 11755
rect 40423 11721 40429 11755
rect 40383 11683 40429 11721
rect 40383 11649 40389 11683
rect 40423 11649 40429 11683
rect 40383 11611 40429 11649
rect 40383 11577 40389 11611
rect 40423 11577 40429 11611
rect 40383 11539 40429 11577
rect 40165 11505 40188 11523
rect 40108 11481 40188 11505
rect 40108 11429 40122 11481
rect 40174 11429 40188 11481
rect 40108 11395 40188 11429
rect 40108 11390 40131 11395
rect 39867 11323 39913 11361
rect 39867 11289 39873 11323
rect 39907 11289 39913 11323
rect 39867 11251 39913 11289
rect 40125 11361 40131 11390
rect 40165 11390 40188 11395
rect 40383 11505 40389 11539
rect 40423 11505 40429 11539
rect 40641 11899 40687 11914
rect 40641 11865 40647 11899
rect 40681 11865 40687 11899
rect 40641 11827 40687 11865
rect 40641 11793 40647 11827
rect 40681 11793 40687 11827
rect 40641 11755 40687 11793
rect 40641 11721 40647 11755
rect 40681 11721 40687 11755
rect 40641 11683 40687 11721
rect 40641 11649 40647 11683
rect 40681 11649 40687 11683
rect 40641 11611 40687 11649
rect 40641 11577 40647 11611
rect 40681 11577 40687 11611
rect 40641 11539 40687 11577
rect 40641 11523 40647 11539
rect 40383 11467 40429 11505
rect 40383 11433 40389 11467
rect 40423 11433 40429 11467
rect 40383 11395 40429 11433
rect 40165 11361 40171 11390
rect 40125 11323 40171 11361
rect 40125 11289 40131 11323
rect 40165 11289 40171 11323
rect 40125 11251 40171 11289
rect 40383 11361 40389 11395
rect 40423 11361 40429 11395
rect 40623 11505 40647 11523
rect 40681 11523 40687 11539
rect 40899 11899 40945 11914
rect 40899 11865 40905 11899
rect 40939 11865 40945 11899
rect 40899 11827 40945 11865
rect 40899 11793 40905 11827
rect 40939 11793 40945 11827
rect 40899 11755 40945 11793
rect 40899 11721 40905 11755
rect 40939 11721 40945 11755
rect 40899 11683 40945 11721
rect 40899 11649 40905 11683
rect 40939 11649 40945 11683
rect 40899 11611 40945 11649
rect 40899 11577 40905 11611
rect 40939 11577 40945 11611
rect 40899 11539 40945 11577
rect 40681 11505 40705 11523
rect 40623 11482 40705 11505
rect 40623 11430 40638 11482
rect 40690 11430 40705 11482
rect 40623 11395 40705 11430
rect 40623 11390 40647 11395
rect 40383 11323 40429 11361
rect 40383 11289 40389 11323
rect 40423 11289 40429 11323
rect 40383 11251 40429 11289
rect 40641 11361 40647 11390
rect 40681 11390 40705 11395
rect 40899 11505 40905 11539
rect 40939 11505 40945 11539
rect 41157 11899 41203 11914
rect 41157 11865 41163 11899
rect 41197 11865 41203 11899
rect 41157 11827 41203 11865
rect 41157 11793 41163 11827
rect 41197 11793 41203 11827
rect 41157 11755 41203 11793
rect 41157 11721 41163 11755
rect 41197 11721 41203 11755
rect 41157 11683 41203 11721
rect 41157 11649 41163 11683
rect 41197 11649 41203 11683
rect 41157 11611 41203 11649
rect 41157 11577 41163 11611
rect 41197 11577 41203 11611
rect 41157 11539 41203 11577
rect 41157 11523 41163 11539
rect 40899 11467 40945 11505
rect 40899 11433 40905 11467
rect 40939 11433 40945 11467
rect 40899 11395 40945 11433
rect 40681 11361 40687 11390
rect 40641 11323 40687 11361
rect 40641 11289 40647 11323
rect 40681 11289 40687 11323
rect 40641 11251 40687 11289
rect 40899 11361 40905 11395
rect 40939 11361 40945 11395
rect 41141 11505 41163 11523
rect 41197 11523 41203 11539
rect 41415 11899 41461 11914
rect 41415 11865 41421 11899
rect 41455 11865 41461 11899
rect 41415 11827 41461 11865
rect 41415 11793 41421 11827
rect 41455 11793 41461 11827
rect 41415 11755 41461 11793
rect 41415 11721 41421 11755
rect 41455 11721 41461 11755
rect 41415 11683 41461 11721
rect 41415 11649 41421 11683
rect 41455 11649 41461 11683
rect 41415 11611 41461 11649
rect 41415 11577 41421 11611
rect 41455 11577 41461 11611
rect 41415 11539 41461 11577
rect 41197 11505 41220 11523
rect 41141 11482 41220 11505
rect 41141 11430 41154 11482
rect 41206 11430 41220 11482
rect 41141 11395 41220 11430
rect 41141 11390 41163 11395
rect 40899 11323 40945 11361
rect 40899 11289 40905 11323
rect 40939 11289 40945 11323
rect 40899 11251 40945 11289
rect 41157 11361 41163 11390
rect 41197 11390 41220 11395
rect 41415 11505 41421 11539
rect 41455 11505 41461 11539
rect 41673 11899 41719 11914
rect 41673 11865 41679 11899
rect 41713 11865 41719 11899
rect 41673 11827 41719 11865
rect 41673 11793 41679 11827
rect 41713 11793 41719 11827
rect 41673 11755 41719 11793
rect 41673 11721 41679 11755
rect 41713 11721 41719 11755
rect 41673 11683 41719 11721
rect 41673 11649 41679 11683
rect 41713 11649 41719 11683
rect 41673 11611 41719 11649
rect 41673 11577 41679 11611
rect 41713 11577 41719 11611
rect 41673 11539 41719 11577
rect 41673 11523 41679 11539
rect 41415 11467 41461 11505
rect 41415 11433 41421 11467
rect 41455 11433 41461 11467
rect 41415 11395 41461 11433
rect 41197 11361 41203 11390
rect 41157 11323 41203 11361
rect 41157 11289 41163 11323
rect 41197 11289 41203 11323
rect 41157 11251 41203 11289
rect 41415 11361 41421 11395
rect 41455 11361 41461 11395
rect 41656 11505 41679 11523
rect 41713 11523 41719 11539
rect 41931 11899 41977 11914
rect 41931 11865 41937 11899
rect 41971 11865 41977 11899
rect 41931 11827 41977 11865
rect 41931 11793 41937 11827
rect 41971 11793 41977 11827
rect 41931 11755 41977 11793
rect 41931 11721 41937 11755
rect 41971 11721 41977 11755
rect 41931 11683 41977 11721
rect 41931 11649 41937 11683
rect 41971 11649 41977 11683
rect 41931 11611 41977 11649
rect 41931 11577 41937 11611
rect 41971 11577 41977 11611
rect 41931 11539 41977 11577
rect 41713 11505 41737 11523
rect 41656 11482 41737 11505
rect 41656 11430 41670 11482
rect 41722 11430 41737 11482
rect 41656 11395 41737 11430
rect 41656 11390 41679 11395
rect 41415 11323 41461 11361
rect 41415 11289 41421 11323
rect 41455 11289 41461 11323
rect 41415 11251 41461 11289
rect 41673 11361 41679 11390
rect 41713 11390 41737 11395
rect 41931 11505 41937 11539
rect 41971 11505 41977 11539
rect 41931 11467 41977 11505
rect 41931 11433 41937 11467
rect 41971 11433 41977 11467
rect 41931 11395 41977 11433
rect 41713 11361 41719 11390
rect 41673 11323 41719 11361
rect 41673 11289 41679 11323
rect 41713 11289 41719 11323
rect 41673 11251 41719 11289
rect 41931 11361 41937 11395
rect 41971 11361 41977 11395
rect 41931 11323 41977 11361
rect 41931 11289 41937 11323
rect 41971 11289 41977 11323
rect 41931 11251 41977 11289
rect 24792 11240 24826 11243
rect 24769 11234 24826 11240
rect 24878 11240 24912 11243
rect 24878 11234 25769 11240
rect 24769 11200 24784 11234
rect 24818 11200 24826 11234
rect 24890 11200 24928 11234
rect 24962 11200 25000 11234
rect 25034 11200 25072 11234
rect 25106 11200 25144 11234
rect 25178 11200 25216 11234
rect 25250 11200 25288 11234
rect 25322 11200 25360 11234
rect 25394 11200 25432 11234
rect 25466 11200 25504 11234
rect 25538 11200 25576 11234
rect 25610 11200 25648 11234
rect 25682 11200 25720 11234
rect 25754 11200 25769 11234
rect 24769 11194 24826 11200
rect 24792 11191 24826 11194
rect 24878 11194 25769 11200
rect 36736 11236 36777 11251
rect 36811 11236 36838 11251
rect 24878 11191 24912 11194
rect 24652 11137 24728 11184
rect 24792 11152 24912 11191
rect 36736 11184 36768 11236
rect 36820 11184 36838 11236
rect 24652 11122 24688 11137
rect 24162 11071 24208 11109
rect 24162 11037 24168 11071
rect 24202 11037 24208 11071
rect 24162 10999 24208 11037
rect 24162 10965 24168 10999
rect 24202 10965 24208 10999
rect 24162 10927 24208 10965
rect 24162 10893 24168 10927
rect 24202 10893 24208 10927
rect 24162 10855 24208 10893
rect 24162 10821 24168 10855
rect 24202 10821 24208 10855
rect 24162 10774 24208 10821
rect 24682 11103 24688 11122
rect 24722 11103 24728 11137
rect 24682 11065 24728 11103
rect 24682 11031 24688 11065
rect 24722 11031 24728 11065
rect 24682 10993 24728 11031
rect 24682 10959 24688 10993
rect 24722 10959 24728 10993
rect 24682 10921 24728 10959
rect 24682 10887 24688 10921
rect 24722 10887 24728 10921
rect 24682 10849 24728 10887
rect 24682 10815 24688 10849
rect 24722 10815 24728 10849
rect 24682 10777 24728 10815
rect 22632 10391 23062 10774
rect 23912 10764 24112 10772
rect 23130 10758 24130 10764
rect 23130 10724 23145 10758
rect 23179 10724 23217 10758
rect 23251 10724 23289 10758
rect 23323 10724 23361 10758
rect 23395 10724 23433 10758
rect 23467 10724 23505 10758
rect 23539 10724 23577 10758
rect 23611 10724 23649 10758
rect 23683 10724 23721 10758
rect 23755 10724 23793 10758
rect 23827 10724 23865 10758
rect 23899 10724 23937 10758
rect 23971 10724 24009 10758
rect 24043 10724 24081 10758
rect 24115 10724 24130 10758
rect 23130 10718 24130 10724
rect 24682 10743 24688 10777
rect 24722 10743 24728 10777
rect 21086 9346 21302 9398
rect 21086 9038 21137 9346
rect 21253 9038 21302 9346
rect 22632 9251 22655 10391
rect 23027 9251 23062 10391
rect 22632 9202 23062 9251
rect 21086 8995 21302 9038
rect 21088 8994 21302 8995
rect 19588 8946 19634 8984
rect 19588 8912 19594 8946
rect 19628 8912 19634 8946
rect 19588 8874 19634 8912
rect 19588 8840 19594 8874
rect 19628 8840 19634 8874
rect 19588 8802 19634 8840
rect 19588 8768 19594 8802
rect 19628 8768 19634 8802
rect 19588 8730 19634 8768
rect 19588 8696 19594 8730
rect 19628 8696 19634 8730
rect 19588 8674 19634 8696
rect 18530 8624 18536 8658
rect 18570 8624 18576 8658
rect 18530 8586 18576 8624
rect 18530 8552 18536 8586
rect 18570 8552 18576 8586
rect 18530 8514 18576 8552
rect 18530 8480 18536 8514
rect 18570 8480 18576 8514
rect 18530 8442 18576 8480
rect 18530 8408 18536 8442
rect 18570 8408 18576 8442
rect 18530 8370 18576 8408
rect 18530 8336 18536 8370
rect 18570 8336 18576 8370
rect 18530 8298 18576 8336
rect 17512 8264 17518 8294
rect 17472 8221 17518 8264
rect 18530 8264 18536 8298
rect 18570 8264 18576 8298
rect 19456 8658 19634 8674
rect 19456 8638 19594 8658
rect 19456 8330 19478 8638
rect 19628 8624 19634 8658
rect 19594 8586 19634 8624
rect 19628 8552 19634 8586
rect 19594 8514 19634 8552
rect 19628 8480 19634 8514
rect 19594 8442 19634 8480
rect 19628 8408 19634 8442
rect 19594 8370 19634 8408
rect 19628 8336 19634 8370
rect 19594 8330 19634 8336
rect 19456 8298 19634 8330
rect 19456 8294 19594 8298
rect 18530 8221 18576 8264
rect 19588 8264 19594 8294
rect 19628 8264 19634 8298
rect 19588 8221 19634 8264
rect 17862 8180 18152 8200
rect 17528 8174 18520 8180
rect 18586 8174 19578 8180
rect 17528 8140 17575 8174
rect 17609 8140 17647 8174
rect 17681 8140 17719 8174
rect 17753 8140 17791 8174
rect 17825 8140 17863 8174
rect 17897 8166 17935 8174
rect 17969 8166 18007 8174
rect 18041 8166 18079 8174
rect 18113 8166 18151 8174
rect 18001 8140 18007 8166
rect 17528 8134 17885 8140
rect 17862 8114 17885 8134
rect 17937 8114 17949 8140
rect 18001 8114 18013 8140
rect 18065 8114 18077 8166
rect 18129 8140 18151 8166
rect 18185 8140 18223 8174
rect 18257 8140 18295 8174
rect 18329 8140 18367 8174
rect 18401 8140 18439 8174
rect 18473 8140 18633 8174
rect 18667 8140 18705 8174
rect 18739 8140 18777 8174
rect 18811 8140 18849 8174
rect 18883 8140 18921 8174
rect 18955 8140 18993 8174
rect 19027 8140 19065 8174
rect 19099 8140 19137 8174
rect 19171 8140 19209 8174
rect 19243 8140 19281 8174
rect 19315 8140 19353 8174
rect 19387 8140 19425 8174
rect 19459 8140 19497 8174
rect 19531 8140 19578 8174
rect 18129 8134 19578 8140
rect 18129 8114 18152 8134
rect 17862 8080 18152 8114
rect 17242 7770 20152 7910
rect 23642 7886 23812 7892
rect 23912 7886 24112 10718
rect 24682 10705 24728 10743
rect 24682 10671 24688 10705
rect 24722 10671 24728 10705
rect 24682 10633 24728 10671
rect 24682 10599 24688 10633
rect 24722 10599 24728 10633
rect 24682 10561 24728 10599
rect 24682 10527 24688 10561
rect 24722 10527 24728 10561
rect 24682 10489 24728 10527
rect 24682 10455 24688 10489
rect 24722 10455 24728 10489
rect 24682 10417 24728 10455
rect 24682 10383 24688 10417
rect 24722 10383 24728 10417
rect 24682 10345 24728 10383
rect 24682 10311 24688 10345
rect 24722 10311 24728 10345
rect 24682 10273 24728 10311
rect 24682 10252 24688 10273
rect 24652 10239 24688 10252
rect 24722 10239 24728 10273
rect 24652 10192 24728 10239
rect 25810 11137 25856 11184
rect 25810 11103 25816 11137
rect 25850 11103 25856 11137
rect 36736 11179 36838 11184
rect 36736 11172 36777 11179
rect 36811 11172 36838 11179
rect 36736 11120 36768 11172
rect 36820 11120 36838 11172
rect 36736 11109 36838 11120
rect 37029 11217 37035 11251
rect 37069 11217 37075 11251
rect 37029 11179 37075 11217
rect 37029 11145 37035 11179
rect 37069 11145 37075 11179
rect 25810 11065 25856 11103
rect 25810 11031 25816 11065
rect 25850 11031 25856 11065
rect 25810 10993 25856 11031
rect 25810 10959 25816 10993
rect 25850 10959 25856 10993
rect 25810 10921 25856 10959
rect 25810 10887 25816 10921
rect 25850 10887 25856 10921
rect 36771 11107 36817 11109
rect 36771 11073 36777 11107
rect 36811 11073 36817 11107
rect 36771 11035 36817 11073
rect 36771 11001 36777 11035
rect 36811 11001 36817 11035
rect 36771 10963 36817 11001
rect 36771 10929 36777 10963
rect 36811 10929 36817 10963
rect 36771 10914 36817 10929
rect 37029 11107 37075 11145
rect 37268 11238 37293 11251
rect 37327 11238 37353 11251
rect 37268 11186 37284 11238
rect 37336 11186 37353 11238
rect 37268 11179 37353 11186
rect 37268 11174 37293 11179
rect 37327 11174 37353 11179
rect 37268 11122 37284 11174
rect 37336 11122 37353 11174
rect 37268 11109 37353 11122
rect 37545 11217 37551 11251
rect 37585 11217 37591 11251
rect 37545 11179 37591 11217
rect 37545 11145 37551 11179
rect 37585 11145 37591 11179
rect 37029 11073 37035 11107
rect 37069 11073 37075 11107
rect 37029 11035 37075 11073
rect 37029 11001 37035 11035
rect 37069 11001 37075 11035
rect 37029 10963 37075 11001
rect 37029 10929 37035 10963
rect 37069 10929 37075 10963
rect 37029 10914 37075 10929
rect 37287 11107 37333 11109
rect 37287 11073 37293 11107
rect 37327 11073 37333 11107
rect 37287 11035 37333 11073
rect 37287 11001 37293 11035
rect 37327 11001 37333 11035
rect 37287 10963 37333 11001
rect 37287 10929 37293 10963
rect 37327 10929 37333 10963
rect 37287 10914 37333 10929
rect 37545 11107 37591 11145
rect 37784 11238 37809 11251
rect 37843 11238 37869 11251
rect 37784 11186 37800 11238
rect 37852 11186 37869 11238
rect 37784 11179 37869 11186
rect 37784 11174 37809 11179
rect 37843 11174 37869 11179
rect 37784 11122 37800 11174
rect 37852 11122 37869 11174
rect 37784 11109 37869 11122
rect 38061 11217 38067 11251
rect 38101 11217 38107 11251
rect 38061 11179 38107 11217
rect 38061 11145 38067 11179
rect 38101 11145 38107 11179
rect 37545 11073 37551 11107
rect 37585 11073 37591 11107
rect 37545 11035 37591 11073
rect 37545 11001 37551 11035
rect 37585 11001 37591 11035
rect 37545 10963 37591 11001
rect 37545 10929 37551 10963
rect 37585 10929 37591 10963
rect 37545 10914 37591 10929
rect 37803 11107 37849 11109
rect 37803 11073 37809 11107
rect 37843 11073 37849 11107
rect 37803 11035 37849 11073
rect 37803 11001 37809 11035
rect 37843 11001 37849 11035
rect 37803 10963 37849 11001
rect 37803 10929 37809 10963
rect 37843 10929 37849 10963
rect 37803 10914 37849 10929
rect 38061 11107 38107 11145
rect 38302 11237 38325 11251
rect 38359 11237 38383 11251
rect 38302 11185 38316 11237
rect 38368 11185 38383 11237
rect 38302 11179 38383 11185
rect 38302 11173 38325 11179
rect 38359 11173 38383 11179
rect 38302 11121 38316 11173
rect 38368 11121 38383 11173
rect 38302 11109 38383 11121
rect 38577 11217 38583 11251
rect 38617 11217 38623 11251
rect 38577 11179 38623 11217
rect 38577 11145 38583 11179
rect 38617 11145 38623 11179
rect 38061 11073 38067 11107
rect 38101 11073 38107 11107
rect 38061 11035 38107 11073
rect 38061 11001 38067 11035
rect 38101 11001 38107 11035
rect 38061 10963 38107 11001
rect 38061 10929 38067 10963
rect 38101 10929 38107 10963
rect 38061 10914 38107 10929
rect 38319 11107 38365 11109
rect 38319 11073 38325 11107
rect 38359 11073 38365 11107
rect 38319 11035 38365 11073
rect 38319 11001 38325 11035
rect 38359 11001 38365 11035
rect 38319 10963 38365 11001
rect 38319 10929 38325 10963
rect 38359 10929 38365 10963
rect 38319 10914 38365 10929
rect 38577 11107 38623 11145
rect 38816 11238 38841 11251
rect 38875 11238 38900 11251
rect 38816 11186 38832 11238
rect 38884 11186 38900 11238
rect 38816 11179 38900 11186
rect 38816 11174 38841 11179
rect 38875 11174 38900 11179
rect 38816 11122 38832 11174
rect 38884 11122 38900 11174
rect 38816 11109 38900 11122
rect 39093 11217 39099 11251
rect 39133 11217 39139 11251
rect 39093 11179 39139 11217
rect 39093 11145 39099 11179
rect 39133 11145 39139 11179
rect 38577 11073 38583 11107
rect 38617 11073 38623 11107
rect 38577 11035 38623 11073
rect 38577 11001 38583 11035
rect 38617 11001 38623 11035
rect 38577 10963 38623 11001
rect 38577 10929 38583 10963
rect 38617 10929 38623 10963
rect 38577 10914 38623 10929
rect 38835 11107 38881 11109
rect 38835 11073 38841 11107
rect 38875 11073 38881 11107
rect 38835 11035 38881 11073
rect 38835 11001 38841 11035
rect 38875 11001 38881 11035
rect 38835 10963 38881 11001
rect 38835 10929 38841 10963
rect 38875 10929 38881 10963
rect 38835 10914 38881 10929
rect 39093 11107 39139 11145
rect 39332 11239 39357 11251
rect 39391 11239 39416 11251
rect 39332 11187 39349 11239
rect 39401 11187 39416 11239
rect 39332 11179 39416 11187
rect 39332 11175 39357 11179
rect 39391 11175 39416 11179
rect 39332 11123 39349 11175
rect 39401 11123 39416 11175
rect 39332 11109 39416 11123
rect 39609 11217 39615 11251
rect 39649 11217 39655 11251
rect 39609 11179 39655 11217
rect 39609 11145 39615 11179
rect 39649 11145 39655 11179
rect 39093 11073 39099 11107
rect 39133 11073 39139 11107
rect 39093 11035 39139 11073
rect 39093 11001 39099 11035
rect 39133 11001 39139 11035
rect 39093 10963 39139 11001
rect 39093 10929 39099 10963
rect 39133 10929 39139 10963
rect 39093 10914 39139 10929
rect 39351 11107 39397 11109
rect 39351 11073 39357 11107
rect 39391 11073 39397 11107
rect 39351 11035 39397 11073
rect 39351 11001 39357 11035
rect 39391 11001 39397 11035
rect 39351 10963 39397 11001
rect 39351 10929 39357 10963
rect 39391 10929 39397 10963
rect 39351 10914 39397 10929
rect 39609 11107 39655 11145
rect 39850 11236 39873 11251
rect 39907 11236 39935 11251
rect 39850 11184 39864 11236
rect 39916 11184 39935 11236
rect 39850 11179 39935 11184
rect 39850 11172 39873 11179
rect 39907 11172 39935 11179
rect 39850 11120 39864 11172
rect 39916 11120 39935 11172
rect 39850 11109 39935 11120
rect 40125 11217 40131 11251
rect 40165 11217 40171 11251
rect 40125 11179 40171 11217
rect 40125 11145 40131 11179
rect 40165 11145 40171 11179
rect 39609 11073 39615 11107
rect 39649 11073 39655 11107
rect 39609 11035 39655 11073
rect 39609 11001 39615 11035
rect 39649 11001 39655 11035
rect 39609 10963 39655 11001
rect 39609 10929 39615 10963
rect 39649 10929 39655 10963
rect 39609 10914 39655 10929
rect 39867 11107 39913 11109
rect 39867 11073 39873 11107
rect 39907 11073 39913 11107
rect 39867 11035 39913 11073
rect 39867 11001 39873 11035
rect 39907 11001 39913 11035
rect 39867 10963 39913 11001
rect 39867 10929 39873 10963
rect 39907 10929 39913 10963
rect 39867 10914 39913 10929
rect 40125 11107 40171 11145
rect 40365 11237 40389 11251
rect 40423 11237 40447 11251
rect 40365 11185 40379 11237
rect 40431 11185 40447 11237
rect 40365 11179 40447 11185
rect 40365 11173 40389 11179
rect 40423 11173 40447 11179
rect 40365 11121 40379 11173
rect 40431 11121 40447 11173
rect 40365 11109 40447 11121
rect 40641 11217 40647 11251
rect 40681 11217 40687 11251
rect 40641 11179 40687 11217
rect 40641 11145 40647 11179
rect 40681 11145 40687 11179
rect 40125 11073 40131 11107
rect 40165 11073 40171 11107
rect 40125 11035 40171 11073
rect 40125 11001 40131 11035
rect 40165 11001 40171 11035
rect 40125 10963 40171 11001
rect 40125 10929 40131 10963
rect 40165 10929 40171 10963
rect 40125 10914 40171 10929
rect 40383 11107 40429 11109
rect 40383 11073 40389 11107
rect 40423 11073 40429 11107
rect 40383 11035 40429 11073
rect 40383 11001 40389 11035
rect 40423 11001 40429 11035
rect 40383 10963 40429 11001
rect 40383 10929 40389 10963
rect 40423 10929 40429 10963
rect 40383 10914 40429 10929
rect 40641 11107 40687 11145
rect 40882 11238 40905 11251
rect 40939 11238 40963 11251
rect 40882 11186 40896 11238
rect 40948 11186 40963 11238
rect 40882 11179 40963 11186
rect 40882 11174 40905 11179
rect 40939 11174 40963 11179
rect 40882 11122 40896 11174
rect 40948 11122 40963 11174
rect 40882 11109 40963 11122
rect 41157 11217 41163 11251
rect 41197 11217 41203 11251
rect 41157 11179 41203 11217
rect 41157 11145 41163 11179
rect 41197 11145 41203 11179
rect 40641 11073 40647 11107
rect 40681 11073 40687 11107
rect 40641 11035 40687 11073
rect 40641 11001 40647 11035
rect 40681 11001 40687 11035
rect 40641 10963 40687 11001
rect 40641 10929 40647 10963
rect 40681 10929 40687 10963
rect 40641 10914 40687 10929
rect 40899 11107 40945 11109
rect 40899 11073 40905 11107
rect 40939 11073 40945 11107
rect 40899 11035 40945 11073
rect 40899 11001 40905 11035
rect 40939 11001 40945 11035
rect 40899 10963 40945 11001
rect 40899 10929 40905 10963
rect 40939 10929 40945 10963
rect 40899 10914 40945 10929
rect 41157 11107 41203 11145
rect 41396 11237 41421 11251
rect 41455 11237 41480 11251
rect 41396 11185 41412 11237
rect 41464 11185 41480 11237
rect 41396 11179 41480 11185
rect 41396 11173 41421 11179
rect 41455 11173 41480 11179
rect 41396 11121 41412 11173
rect 41464 11121 41480 11173
rect 41396 11109 41480 11121
rect 41673 11217 41679 11251
rect 41713 11217 41719 11251
rect 41673 11179 41719 11217
rect 41673 11145 41679 11179
rect 41713 11145 41719 11179
rect 41157 11073 41163 11107
rect 41197 11073 41203 11107
rect 41157 11035 41203 11073
rect 41157 11001 41163 11035
rect 41197 11001 41203 11035
rect 41157 10963 41203 11001
rect 41157 10929 41163 10963
rect 41197 10929 41203 10963
rect 41157 10914 41203 10929
rect 41415 11107 41461 11109
rect 41415 11073 41421 11107
rect 41455 11073 41461 11107
rect 41415 11035 41461 11073
rect 41415 11001 41421 11035
rect 41455 11001 41461 11035
rect 41415 10963 41461 11001
rect 41415 10929 41421 10963
rect 41455 10929 41461 10963
rect 41415 10914 41461 10929
rect 41673 11107 41719 11145
rect 41913 11237 41937 11251
rect 41971 11237 41996 11251
rect 41913 11185 41928 11237
rect 41980 11185 41996 11237
rect 41913 11179 41996 11185
rect 41913 11173 41937 11179
rect 41971 11173 41996 11179
rect 41913 11121 41928 11173
rect 41980 11121 41996 11173
rect 41913 11109 41996 11121
rect 41673 11073 41679 11107
rect 41713 11073 41719 11107
rect 41673 11035 41719 11073
rect 41673 11001 41679 11035
rect 41713 11001 41719 11035
rect 41673 10963 41719 11001
rect 41673 10929 41679 10963
rect 41713 10929 41719 10963
rect 41673 10914 41719 10929
rect 41931 11107 41977 11109
rect 41931 11073 41937 11107
rect 41971 11073 41977 11107
rect 41931 11035 41977 11073
rect 41931 11001 41937 11035
rect 41971 11001 41977 11035
rect 41931 10963 41977 11001
rect 41931 10929 41937 10963
rect 41971 10929 41977 10963
rect 41931 10914 41977 10929
rect 25810 10849 25856 10887
rect 25810 10815 25816 10849
rect 25850 10815 25856 10849
rect 36827 10876 37019 10882
rect 36827 10842 36870 10876
rect 36904 10842 36942 10876
rect 36976 10842 37019 10876
rect 36827 10836 37019 10842
rect 37085 10876 37277 10882
rect 37085 10842 37128 10876
rect 37162 10842 37200 10876
rect 37234 10842 37277 10876
rect 37085 10836 37277 10842
rect 37343 10876 37535 10882
rect 37343 10842 37386 10876
rect 37420 10842 37458 10876
rect 37492 10842 37535 10876
rect 37343 10836 37535 10842
rect 37601 10876 37793 10882
rect 37601 10842 37644 10876
rect 37678 10842 37716 10876
rect 37750 10842 37793 10876
rect 37601 10836 37793 10842
rect 37859 10876 38051 10882
rect 37859 10842 37902 10876
rect 37936 10842 37974 10876
rect 38008 10842 38051 10876
rect 37859 10836 38051 10842
rect 38117 10876 38309 10882
rect 38117 10842 38160 10876
rect 38194 10842 38232 10876
rect 38266 10842 38309 10876
rect 38117 10836 38309 10842
rect 38375 10876 38567 10882
rect 38375 10842 38418 10876
rect 38452 10842 38490 10876
rect 38524 10842 38567 10876
rect 38375 10836 38567 10842
rect 38633 10876 38825 10882
rect 38633 10842 38676 10876
rect 38710 10842 38748 10876
rect 38782 10842 38825 10876
rect 38633 10836 38825 10842
rect 38891 10876 39083 10882
rect 38891 10842 38934 10876
rect 38968 10842 39006 10876
rect 39040 10842 39083 10876
rect 38891 10836 39083 10842
rect 39149 10876 39341 10882
rect 39149 10842 39192 10876
rect 39226 10842 39264 10876
rect 39298 10842 39341 10876
rect 39149 10836 39341 10842
rect 39407 10876 39599 10882
rect 39407 10842 39450 10876
rect 39484 10842 39522 10876
rect 39556 10842 39599 10876
rect 39407 10836 39599 10842
rect 39665 10876 39857 10882
rect 39665 10842 39708 10876
rect 39742 10842 39780 10876
rect 39814 10842 39857 10876
rect 39665 10836 39857 10842
rect 39923 10876 40115 10882
rect 39923 10842 39966 10876
rect 40000 10842 40038 10876
rect 40072 10842 40115 10876
rect 39923 10836 40115 10842
rect 40181 10876 40373 10882
rect 40181 10842 40224 10876
rect 40258 10842 40296 10876
rect 40330 10842 40373 10876
rect 40181 10836 40373 10842
rect 40439 10876 40631 10882
rect 40439 10842 40482 10876
rect 40516 10842 40554 10876
rect 40588 10842 40631 10876
rect 40439 10836 40631 10842
rect 40697 10876 40889 10882
rect 40697 10842 40740 10876
rect 40774 10842 40812 10876
rect 40846 10842 40889 10876
rect 40697 10836 40889 10842
rect 40955 10876 41147 10882
rect 40955 10842 40998 10876
rect 41032 10842 41070 10876
rect 41104 10842 41147 10876
rect 40955 10836 41147 10842
rect 41213 10876 41405 10882
rect 41213 10842 41256 10876
rect 41290 10842 41328 10876
rect 41362 10842 41405 10876
rect 41213 10836 41405 10842
rect 41471 10876 41663 10882
rect 41471 10842 41514 10876
rect 41548 10842 41586 10876
rect 41620 10842 41663 10876
rect 41471 10836 41663 10842
rect 41729 10876 41921 10882
rect 41729 10842 41772 10876
rect 41806 10842 41844 10876
rect 41878 10842 41921 10876
rect 41729 10836 41921 10842
rect 25810 10777 25856 10815
rect 25810 10743 25816 10777
rect 25850 10743 25856 10777
rect 36823 10776 41921 10836
rect 25810 10705 25856 10743
rect 25810 10671 25816 10705
rect 25850 10671 25856 10705
rect 25810 10633 25856 10671
rect 25810 10599 25816 10633
rect 25850 10599 25856 10633
rect 25810 10561 25856 10599
rect 37862 10627 40842 10776
rect 37862 10621 38110 10627
rect 37862 10587 37905 10621
rect 37939 10587 37977 10621
rect 38011 10587 38110 10621
rect 37862 10581 38110 10587
rect 38328 10621 38520 10627
rect 38328 10587 38371 10621
rect 38405 10587 38443 10621
rect 38477 10587 38520 10621
rect 38328 10581 38520 10587
rect 38586 10621 38778 10627
rect 38586 10587 38629 10621
rect 38663 10587 38701 10621
rect 38735 10587 38778 10621
rect 38586 10581 38778 10587
rect 38844 10621 39036 10627
rect 38844 10587 38887 10621
rect 38921 10587 38959 10621
rect 38993 10587 39036 10621
rect 38844 10581 39036 10587
rect 39102 10621 39294 10627
rect 39102 10587 39145 10621
rect 39179 10587 39217 10621
rect 39251 10587 39294 10621
rect 39102 10581 39294 10587
rect 39360 10621 39552 10627
rect 39360 10587 39403 10621
rect 39437 10587 39475 10621
rect 39509 10587 39552 10621
rect 39360 10581 39552 10587
rect 39618 10621 39810 10627
rect 39618 10587 39661 10621
rect 39695 10587 39733 10621
rect 39767 10587 39810 10621
rect 39618 10581 39810 10587
rect 39876 10621 40068 10627
rect 39876 10587 39919 10621
rect 39953 10587 39991 10621
rect 40025 10587 40068 10621
rect 39876 10581 40068 10587
rect 40134 10621 40326 10627
rect 40134 10587 40177 10621
rect 40211 10587 40249 10621
rect 40283 10587 40326 10621
rect 40134 10581 40326 10587
rect 40392 10621 40584 10627
rect 40392 10587 40435 10621
rect 40469 10587 40507 10621
rect 40541 10587 40584 10621
rect 40392 10581 40584 10587
rect 40650 10621 40842 10627
rect 40650 10587 40693 10621
rect 40727 10587 40765 10621
rect 40799 10587 40842 10621
rect 40650 10581 40842 10587
rect 25810 10527 25816 10561
rect 25850 10527 25856 10561
rect 37806 10538 37852 10549
rect 25810 10489 25856 10527
rect 25810 10455 25816 10489
rect 25850 10455 25856 10489
rect 25810 10417 25856 10455
rect 25810 10383 25816 10417
rect 25850 10383 25856 10417
rect 25810 10345 25856 10383
rect 25810 10311 25816 10345
rect 25850 10311 25856 10345
rect 25810 10273 25856 10311
rect 25810 10239 25816 10273
rect 25850 10239 25856 10273
rect 25632 10198 25762 10232
rect 24652 10126 24682 10192
rect 25632 10182 25671 10198
rect 24769 10176 25671 10182
rect 25723 10182 25762 10198
rect 25810 10192 25856 10239
rect 37730 10534 37852 10538
rect 37730 10500 37812 10534
rect 37846 10500 37852 10534
rect 37730 10462 37852 10500
rect 37730 10428 37812 10462
rect 37846 10428 37852 10462
rect 37730 10390 37852 10428
rect 37730 10356 37812 10390
rect 37846 10356 37852 10390
rect 37730 10318 37852 10356
rect 37730 10284 37812 10318
rect 37846 10284 37852 10318
rect 37730 10246 37852 10284
rect 37730 10212 37812 10246
rect 37846 10212 37852 10246
rect 25723 10176 25769 10182
rect 24769 10142 24784 10176
rect 24818 10142 24856 10176
rect 24890 10142 24928 10176
rect 24962 10142 25000 10176
rect 25034 10142 25072 10176
rect 25106 10142 25144 10176
rect 25178 10142 25216 10176
rect 25250 10142 25288 10176
rect 25322 10142 25360 10176
rect 25394 10142 25432 10176
rect 25466 10142 25504 10176
rect 25538 10142 25576 10176
rect 25610 10142 25648 10176
rect 25682 10142 25720 10146
rect 25754 10142 25769 10176
rect 24769 10136 25769 10142
rect 37730 10174 37852 10212
rect 37730 10140 37812 10174
rect 37846 10140 37852 10174
rect 25632 10132 25762 10136
rect 24652 10079 24728 10126
rect 24652 10062 24688 10079
rect 24682 10045 24688 10062
rect 24722 10045 24728 10079
rect 24682 10007 24728 10045
rect 24682 9973 24688 10007
rect 24722 9973 24728 10007
rect 24682 9935 24728 9973
rect 24682 9901 24688 9935
rect 24722 9901 24728 9935
rect 24682 9863 24728 9901
rect 24682 9829 24688 9863
rect 24722 9829 24728 9863
rect 24682 9791 24728 9829
rect 24682 9757 24688 9791
rect 24722 9757 24728 9791
rect 24682 9719 24728 9757
rect 24682 9685 24688 9719
rect 24722 9685 24728 9719
rect 24682 9647 24728 9685
rect 24682 9613 24688 9647
rect 24722 9613 24728 9647
rect 24682 9575 24728 9613
rect 24682 9541 24688 9575
rect 24722 9541 24728 9575
rect 24682 9503 24728 9541
rect 24682 9469 24688 9503
rect 24722 9469 24728 9503
rect 24682 9431 24728 9469
rect 24682 9397 24688 9431
rect 24722 9397 24728 9431
rect 24682 9359 24728 9397
rect 24682 9325 24688 9359
rect 24722 9325 24728 9359
rect 24682 9287 24728 9325
rect 24682 9253 24688 9287
rect 24722 9253 24728 9287
rect 24682 9215 24728 9253
rect 24682 9181 24688 9215
rect 24722 9181 24728 9215
rect 24682 9134 24728 9181
rect 25810 10079 25856 10126
rect 25810 10045 25816 10079
rect 25850 10045 25856 10079
rect 25810 10007 25856 10045
rect 25810 9973 25816 10007
rect 25850 9973 25856 10007
rect 25810 9935 25856 9973
rect 25810 9901 25816 9935
rect 25850 9901 25856 9935
rect 25810 9863 25856 9901
rect 25810 9829 25816 9863
rect 25850 9829 25856 9863
rect 25810 9791 25856 9829
rect 25810 9757 25816 9791
rect 25850 9757 25856 9791
rect 25810 9719 25856 9757
rect 25810 9685 25816 9719
rect 25850 9685 25856 9719
rect 25810 9647 25856 9685
rect 25810 9613 25816 9647
rect 25850 9613 25856 9647
rect 25810 9575 25856 9613
rect 25810 9541 25816 9575
rect 25850 9541 25856 9575
rect 25810 9503 25856 9541
rect 25810 9469 25816 9503
rect 25850 9469 25856 9503
rect 25810 9431 25856 9469
rect 25810 9397 25816 9431
rect 25850 9397 25856 9431
rect 25810 9359 25856 9397
rect 25810 9325 25816 9359
rect 25850 9325 25856 9359
rect 25810 9287 25856 9325
rect 25810 9253 25816 9287
rect 25850 9253 25856 9287
rect 25810 9215 25856 9253
rect 25810 9181 25816 9215
rect 25850 9181 25856 9215
rect 24792 9138 24912 9162
rect 24792 9124 24826 9138
rect 24769 9118 24826 9124
rect 24878 9124 24912 9138
rect 25810 9134 25856 9181
rect 37730 10102 37852 10140
rect 37730 10068 37812 10102
rect 37846 10068 37852 10102
rect 37730 10030 37852 10068
rect 37730 9996 37812 10030
rect 37846 9996 37852 10030
rect 37730 9958 37852 9996
rect 37730 9924 37812 9958
rect 37846 9924 37852 9958
rect 37730 9886 37852 9924
rect 37730 9852 37812 9886
rect 37846 9852 37852 9886
rect 37730 9814 37852 9852
rect 37730 9780 37812 9814
rect 37846 9780 37852 9814
rect 37730 9742 37852 9780
rect 37730 9708 37812 9742
rect 37846 9708 37852 9742
rect 37730 9670 37852 9708
rect 37730 9636 37812 9670
rect 37846 9636 37852 9670
rect 37730 9598 37852 9636
rect 37730 9564 37812 9598
rect 37846 9564 37852 9598
rect 37730 9549 37852 9564
rect 38064 10534 38110 10581
rect 38064 10500 38070 10534
rect 38104 10500 38110 10534
rect 38064 10462 38110 10500
rect 38064 10428 38070 10462
rect 38104 10428 38110 10462
rect 38064 10390 38110 10428
rect 38064 10356 38070 10390
rect 38104 10356 38110 10390
rect 38064 10318 38110 10356
rect 38064 10284 38070 10318
rect 38104 10284 38110 10318
rect 38064 10246 38110 10284
rect 38064 10212 38070 10246
rect 38104 10212 38110 10246
rect 38064 10174 38110 10212
rect 38064 10140 38070 10174
rect 38104 10140 38110 10174
rect 38064 10102 38110 10140
rect 38064 10068 38070 10102
rect 38104 10068 38110 10102
rect 38064 10030 38110 10068
rect 38064 9996 38070 10030
rect 38104 9996 38110 10030
rect 38064 9958 38110 9996
rect 38064 9924 38070 9958
rect 38104 9924 38110 9958
rect 38064 9886 38110 9924
rect 38272 10534 38318 10549
rect 38272 10500 38278 10534
rect 38312 10500 38318 10534
rect 38272 10462 38318 10500
rect 38272 10428 38278 10462
rect 38312 10428 38318 10462
rect 38272 10390 38318 10428
rect 38272 10356 38278 10390
rect 38312 10356 38318 10390
rect 38272 10318 38318 10356
rect 38272 10284 38278 10318
rect 38312 10284 38318 10318
rect 38272 10246 38318 10284
rect 38272 10212 38278 10246
rect 38312 10212 38318 10246
rect 38530 10534 38576 10549
rect 38530 10500 38536 10534
rect 38570 10500 38576 10534
rect 38530 10462 38576 10500
rect 38530 10428 38536 10462
rect 38570 10428 38576 10462
rect 38530 10390 38576 10428
rect 38530 10356 38536 10390
rect 38570 10356 38576 10390
rect 38530 10318 38576 10356
rect 38530 10284 38536 10318
rect 38570 10284 38576 10318
rect 38530 10246 38576 10284
rect 38530 10245 38536 10246
rect 38272 10174 38318 10212
rect 38272 10140 38278 10174
rect 38312 10140 38318 10174
rect 38272 10102 38318 10140
rect 38272 10068 38278 10102
rect 38312 10068 38318 10102
rect 38504 10228 38536 10245
rect 38570 10245 38576 10246
rect 38788 10534 38834 10549
rect 38788 10500 38794 10534
rect 38828 10500 38834 10534
rect 38788 10462 38834 10500
rect 38788 10428 38794 10462
rect 38828 10428 38834 10462
rect 38788 10390 38834 10428
rect 38788 10356 38794 10390
rect 38828 10356 38834 10390
rect 38788 10318 38834 10356
rect 38788 10284 38794 10318
rect 38828 10284 38834 10318
rect 38788 10246 38834 10284
rect 38570 10228 38601 10245
rect 38504 10176 38527 10228
rect 38579 10176 38601 10228
rect 38504 10174 38601 10176
rect 38504 10164 38536 10174
rect 38570 10164 38601 10174
rect 38504 10112 38527 10164
rect 38579 10112 38601 10164
rect 38504 10102 38601 10112
rect 38504 10093 38536 10102
rect 38272 10030 38318 10068
rect 38272 9996 38278 10030
rect 38312 9996 38318 10030
rect 38272 9958 38318 9996
rect 38272 9924 38278 9958
rect 38312 9924 38318 9958
rect 38272 9914 38318 9924
rect 38530 10068 38536 10093
rect 38570 10093 38601 10102
rect 38788 10212 38794 10246
rect 38828 10212 38834 10246
rect 39046 10534 39092 10549
rect 39046 10500 39052 10534
rect 39086 10500 39092 10534
rect 39046 10462 39092 10500
rect 39046 10428 39052 10462
rect 39086 10428 39092 10462
rect 39046 10390 39092 10428
rect 39046 10356 39052 10390
rect 39086 10356 39092 10390
rect 39046 10318 39092 10356
rect 39046 10284 39052 10318
rect 39086 10284 39092 10318
rect 39046 10246 39092 10284
rect 39046 10245 39052 10246
rect 38788 10174 38834 10212
rect 38788 10140 38794 10174
rect 38828 10140 38834 10174
rect 38788 10102 38834 10140
rect 38570 10068 38576 10093
rect 38530 10030 38576 10068
rect 38530 9996 38536 10030
rect 38570 9996 38576 10030
rect 38530 9958 38576 9996
rect 38530 9924 38536 9958
rect 38570 9924 38576 9958
rect 38064 9852 38070 9886
rect 38104 9852 38110 9886
rect 38064 9814 38110 9852
rect 38064 9780 38070 9814
rect 38104 9780 38110 9814
rect 38064 9742 38110 9780
rect 38064 9708 38070 9742
rect 38104 9708 38110 9742
rect 38257 9886 38335 9914
rect 38257 9878 38278 9886
rect 38312 9878 38335 9886
rect 38257 9826 38270 9878
rect 38322 9826 38335 9878
rect 38257 9814 38335 9826
rect 38257 9762 38270 9814
rect 38322 9762 38335 9814
rect 38257 9742 38335 9762
rect 38257 9729 38278 9742
rect 38064 9670 38110 9708
rect 38064 9636 38070 9670
rect 38104 9636 38110 9670
rect 38064 9598 38110 9636
rect 38064 9564 38070 9598
rect 38104 9564 38110 9598
rect 24878 9118 25769 9124
rect 24769 9084 24784 9118
rect 24818 9086 24826 9118
rect 24818 9084 24856 9086
rect 24890 9084 24928 9118
rect 24962 9084 25000 9118
rect 25034 9084 25072 9118
rect 25106 9084 25144 9118
rect 25178 9084 25216 9118
rect 25250 9084 25288 9118
rect 25322 9084 25360 9118
rect 25394 9084 25432 9118
rect 25466 9084 25504 9118
rect 25538 9084 25576 9118
rect 25610 9084 25648 9118
rect 25682 9084 25720 9118
rect 25754 9084 25769 9118
rect 24769 9078 25769 9084
rect 24792 9072 24912 9078
rect 25402 8427 26382 8462
rect 25402 8162 26222 8427
rect 25142 7886 25302 7892
rect 23610 7880 24610 7886
rect 23610 7846 23625 7880
rect 23659 7873 23697 7880
rect 23731 7873 23769 7880
rect 23659 7846 23664 7873
rect 23803 7846 23841 7880
rect 23875 7846 23913 7880
rect 23947 7846 23985 7880
rect 24019 7846 24057 7880
rect 24091 7846 24129 7880
rect 24163 7846 24201 7880
rect 24235 7846 24273 7880
rect 24307 7846 24345 7880
rect 24379 7846 24417 7880
rect 24451 7846 24489 7880
rect 24523 7846 24561 7880
rect 24595 7846 24610 7880
rect 23610 7840 23664 7846
rect 17052 7633 19932 7660
rect 16832 7620 19932 7633
rect 16832 7586 17531 7620
rect 17565 7586 17603 7620
rect 17637 7586 17675 7620
rect 17709 7586 17747 7620
rect 17781 7586 17819 7620
rect 17853 7586 17891 7620
rect 17925 7586 17963 7620
rect 17997 7586 18035 7620
rect 18069 7586 18107 7620
rect 18141 7586 18179 7620
rect 18213 7586 18251 7620
rect 18285 7586 18323 7620
rect 18357 7586 18395 7620
rect 18429 7590 18981 7620
rect 18429 7586 18532 7590
rect 16832 7580 18532 7586
rect 18934 7586 18981 7590
rect 19015 7586 19053 7620
rect 19087 7586 19125 7620
rect 19159 7586 19197 7620
rect 19231 7586 19269 7620
rect 19303 7586 19341 7620
rect 19375 7586 19413 7620
rect 19447 7586 19485 7620
rect 19519 7586 19557 7620
rect 19591 7586 19629 7620
rect 19663 7586 19701 7620
rect 19735 7586 19773 7620
rect 19807 7586 19845 7620
rect 19879 7590 19932 7620
rect 19879 7586 19926 7590
rect 18934 7580 19926 7586
rect 13676 7516 13746 7530
rect -3618 6809 -3596 6811
rect -3675 6798 -3596 6809
rect -3675 6746 -3662 6798
rect -3610 6746 -3596 6798
rect -3675 6737 -3652 6746
rect -3618 6737 -3596 6746
rect -3675 6734 -3596 6737
rect -3675 6682 -3662 6734
rect -3610 6682 -3596 6734
rect -3675 6670 -3652 6682
rect -3618 6670 -3596 6682
rect -3675 6618 -3662 6670
rect -3610 6618 -3596 6670
rect -3675 6606 -3652 6618
rect -3916 6555 -3870 6593
rect -3916 6521 -3910 6555
rect -3876 6521 -3870 6555
rect -3916 6483 -3870 6521
rect -3916 6449 -3910 6483
rect -3876 6449 -3870 6483
rect -3916 6411 -3870 6449
rect -3916 6377 -3910 6411
rect -3876 6377 -3870 6411
rect -3916 6339 -3870 6377
rect -3916 6305 -3910 6339
rect -3876 6305 -3870 6339
rect -3916 6267 -3870 6305
rect -3916 6233 -3910 6267
rect -3876 6233 -3870 6267
rect -3916 6195 -3870 6233
rect -3916 6161 -3910 6195
rect -3876 6161 -3870 6195
rect -3916 6123 -3870 6161
rect -3916 6089 -3910 6123
rect -3876 6089 -3870 6123
rect -3916 6051 -3870 6089
rect -3916 6017 -3910 6051
rect -3876 6017 -3870 6051
rect -3916 5979 -3870 6017
rect -3916 5945 -3910 5979
rect -3876 5945 -3870 5979
rect -3916 5907 -3870 5945
rect -3916 5901 -3910 5907
rect -4174 5835 -4128 5873
rect -4174 5801 -4168 5835
rect -4134 5801 -4128 5835
rect -4174 5763 -4128 5801
rect -4174 5729 -4168 5763
rect -4134 5729 -4128 5763
rect -4690 5657 -4684 5691
rect -4650 5657 -4644 5691
rect -4690 5619 -4644 5657
rect -4690 5585 -4684 5619
rect -4650 5585 -4644 5619
rect -4690 5538 -4644 5585
rect -4432 5691 -4386 5693
rect -4432 5657 -4426 5691
rect -4392 5657 -4386 5691
rect -4432 5619 -4386 5657
rect -4432 5585 -4426 5619
rect -4392 5585 -4386 5619
rect -4432 5538 -4386 5585
rect -4174 5691 -4128 5729
rect -3932 5887 -3910 5901
rect -3876 5901 -3870 5907
rect -3658 6593 -3652 6606
rect -3618 6606 -3596 6618
rect 13066 6700 13746 7516
rect 16412 7452 16662 7560
rect 16402 7176 16662 7452
rect 17428 7505 17474 7548
rect 17428 7471 17434 7505
rect 17468 7471 17474 7505
rect 18462 7505 18532 7580
rect 18462 7480 18492 7505
rect 17428 7433 17474 7471
rect 17428 7399 17434 7433
rect 17468 7399 17474 7433
rect 17428 7361 17474 7399
rect 17428 7327 17434 7361
rect 17468 7327 17474 7361
rect 17428 7289 17474 7327
rect 17428 7255 17434 7289
rect 17468 7255 17474 7289
rect 17428 7240 17474 7255
rect 18486 7471 18492 7480
rect 18526 7471 18532 7505
rect 18486 7433 18532 7471
rect 18486 7399 18492 7433
rect 18526 7399 18532 7433
rect 18486 7361 18532 7399
rect 18486 7327 18492 7361
rect 18526 7327 18532 7361
rect 18486 7289 18532 7327
rect 18486 7255 18492 7289
rect 18526 7255 18532 7289
rect 16220 7090 16270 7104
rect 16220 7056 16228 7090
rect 16262 7056 16270 7090
rect 16220 7018 16270 7056
rect 16220 6984 16228 7018
rect 16262 6984 16270 7018
rect 16220 6946 16270 6984
rect 16220 6912 16228 6946
rect 16262 6912 16270 6946
rect 16220 6874 16270 6912
rect 16220 6840 16228 6874
rect 16262 6840 16270 6874
rect 16220 6802 16270 6840
rect 13066 6666 13142 6700
rect 13176 6666 13242 6700
rect 13276 6666 13342 6700
rect 13376 6666 13442 6700
rect 13476 6666 13542 6700
rect 13576 6666 13642 6700
rect 13676 6666 13746 6700
rect -3618 6593 -3612 6606
rect -3658 6555 -3612 6593
rect 13066 6600 13746 6666
rect 13066 6570 13142 6600
rect -3658 6521 -3652 6555
rect -3618 6521 -3612 6555
rect -3658 6483 -3612 6521
rect -3658 6449 -3652 6483
rect -3618 6449 -3612 6483
rect -3658 6411 -3612 6449
rect -3658 6377 -3652 6411
rect -3618 6377 -3612 6411
rect -3658 6339 -3612 6377
rect -3658 6305 -3652 6339
rect -3618 6305 -3612 6339
rect -3658 6267 -3612 6305
rect -3658 6233 -3652 6267
rect -3618 6233 -3612 6267
rect -3658 6195 -3612 6233
rect -3658 6161 -3652 6195
rect -3618 6161 -3612 6195
rect 13111 6566 13142 6570
rect 13176 6566 13242 6600
rect 13276 6566 13342 6600
rect 13376 6566 13442 6600
rect 13476 6566 13542 6600
rect 13576 6566 13642 6600
rect 13676 6570 13746 6600
rect 14761 6730 15371 6775
rect 14761 6696 14792 6730
rect 14826 6696 14892 6730
rect 14926 6696 14992 6730
rect 15026 6696 15092 6730
rect 15126 6696 15192 6730
rect 15226 6696 15292 6730
rect 15326 6696 15371 6730
rect 14761 6630 15371 6696
rect 16220 6768 16228 6802
rect 16262 6768 16270 6802
rect 16220 6730 16270 6768
rect 16220 6696 16228 6730
rect 16262 6696 16270 6730
rect 16220 6683 16270 6696
rect 16422 7090 16662 7176
rect 17422 7217 17742 7240
rect 17422 7183 17434 7217
rect 17468 7183 17742 7217
rect 17422 7180 17742 7183
rect 17422 7145 17455 7180
rect 17422 7111 17434 7145
rect 16422 7056 16546 7090
rect 16580 7056 16662 7090
rect 16422 7018 16662 7056
rect 16422 6984 16546 7018
rect 16580 6984 16662 7018
rect 16422 6946 16662 6984
rect 16422 6912 16546 6946
rect 16580 6912 16662 6946
rect 16422 6874 16662 6912
rect 16422 6840 16546 6874
rect 16580 6840 16662 6874
rect 16422 6802 16662 6840
rect 16422 6768 16546 6802
rect 16580 6768 16662 6802
rect 16422 6730 16662 6768
rect 16422 6696 16546 6730
rect 16580 6696 16662 6730
rect 14761 6596 14792 6630
rect 14826 6596 14892 6630
rect 14926 6596 14992 6630
rect 15026 6596 15092 6630
rect 15126 6596 15192 6630
rect 15226 6596 15292 6630
rect 15326 6596 15371 6630
rect 13676 6566 13721 6570
rect 13111 6500 13721 6566
rect 13111 6466 13142 6500
rect 13176 6466 13242 6500
rect 13276 6466 13342 6500
rect 13376 6466 13442 6500
rect 13476 6466 13542 6500
rect 13576 6466 13642 6500
rect 13676 6466 13721 6500
rect 13111 6400 13721 6466
rect 13111 6366 13142 6400
rect 13176 6366 13242 6400
rect 13276 6366 13342 6400
rect 13376 6366 13442 6400
rect 13476 6366 13542 6400
rect 13576 6366 13642 6400
rect 13676 6366 13721 6400
rect 13111 6300 13721 6366
rect 13111 6266 13142 6300
rect 13176 6266 13242 6300
rect 13276 6266 13342 6300
rect 13376 6266 13442 6300
rect 13476 6266 13542 6300
rect 13576 6266 13642 6300
rect 13676 6266 13721 6300
rect 13111 6200 13721 6266
rect 13111 6170 13142 6200
rect -3658 6123 -3612 6161
rect -3658 6089 -3652 6123
rect -3618 6089 -3612 6123
rect -3658 6051 -3612 6089
rect -3658 6017 -3652 6051
rect -3618 6017 -3612 6051
rect -3658 5979 -3612 6017
rect -3658 5945 -3652 5979
rect -3618 5945 -3612 5979
rect -3658 5907 -3612 5945
rect -3876 5887 -3852 5901
rect -3932 5835 -3919 5887
rect -3867 5835 -3852 5887
rect -3932 5823 -3910 5835
rect -3876 5823 -3852 5835
rect -3932 5771 -3919 5823
rect -3867 5771 -3852 5823
rect -3932 5763 -3852 5771
rect -3932 5759 -3910 5763
rect -3876 5759 -3852 5763
rect -3932 5707 -3919 5759
rect -3867 5707 -3852 5759
rect -3932 5693 -3852 5707
rect -3658 5873 -3652 5907
rect -3618 5873 -3612 5907
rect 13066 6166 13142 6170
rect 13176 6166 13242 6200
rect 13276 6166 13342 6200
rect 13376 6166 13442 6200
rect 13476 6166 13542 6200
rect 13576 6166 13642 6200
rect 13676 6170 13721 6200
rect 14761 6530 15371 6596
rect 14761 6496 14792 6530
rect 14826 6496 14892 6530
rect 14926 6496 14992 6530
rect 15026 6496 15092 6530
rect 15126 6496 15192 6530
rect 15226 6496 15292 6530
rect 15326 6496 15371 6530
rect 14761 6430 15371 6496
rect 14761 6396 14792 6430
rect 14826 6396 14892 6430
rect 14926 6396 14992 6430
rect 15026 6396 15092 6430
rect 15126 6396 15192 6430
rect 15226 6396 15292 6430
rect 15326 6396 15371 6430
rect 14761 6330 15371 6396
rect 14761 6296 14792 6330
rect 14826 6296 14892 6330
rect 14926 6296 14992 6330
rect 15026 6296 15092 6330
rect 15126 6296 15192 6330
rect 15226 6296 15292 6330
rect 15326 6296 15371 6330
rect 16422 6539 16662 6696
rect 16856 7090 16906 7104
rect 16856 7056 16864 7090
rect 16898 7056 16906 7090
rect 16856 7018 16906 7056
rect 16856 6984 16864 7018
rect 16898 6984 16906 7018
rect 16856 6946 16906 6984
rect 16856 6912 16864 6946
rect 16898 6912 16906 6946
rect 17422 7073 17455 7111
rect 17422 7039 17434 7073
rect 17422 7001 17455 7039
rect 17422 6967 17434 7001
rect 17699 7000 17742 7180
rect 17468 6967 17742 7000
rect 17422 6940 17742 6967
rect 18486 7217 18532 7255
rect 18486 7183 18492 7217
rect 18526 7183 18532 7217
rect 18486 7145 18532 7183
rect 18486 7111 18492 7145
rect 18526 7111 18532 7145
rect 18486 7073 18532 7111
rect 18486 7039 18492 7073
rect 18526 7039 18532 7073
rect 18486 7001 18532 7039
rect 18486 6967 18492 7001
rect 18526 6967 18532 7001
rect 16856 6874 16906 6912
rect 16856 6840 16864 6874
rect 16898 6840 16906 6874
rect 16856 6802 16906 6840
rect 16856 6768 16864 6802
rect 16898 6768 16906 6802
rect 16856 6730 16906 6768
rect 16856 6696 16864 6730
rect 16898 6696 16906 6730
rect 16856 6683 16906 6696
rect 17428 6929 17474 6940
rect 17428 6895 17434 6929
rect 17468 6895 17474 6929
rect 17428 6857 17474 6895
rect 17428 6823 17434 6857
rect 17468 6823 17474 6857
rect 17428 6785 17474 6823
rect 17428 6751 17434 6785
rect 17468 6751 17474 6785
rect 17428 6713 17474 6751
rect 16422 6359 16436 6539
rect 16616 6359 16662 6539
rect 16422 6302 16662 6359
rect 17428 6679 17434 6713
rect 17468 6679 17474 6713
rect 17428 6641 17474 6679
rect 17428 6607 17434 6641
rect 17468 6607 17474 6641
rect 17428 6569 17474 6607
rect 17428 6535 17434 6569
rect 17468 6535 17474 6569
rect 17428 6497 17474 6535
rect 17428 6463 17434 6497
rect 17468 6463 17474 6497
rect 17428 6425 17474 6463
rect 17428 6391 17434 6425
rect 17468 6391 17474 6425
rect 17428 6353 17474 6391
rect 17428 6319 17434 6353
rect 17468 6319 17474 6353
rect 14761 6230 15371 6296
rect 14761 6196 14792 6230
rect 14826 6196 14892 6230
rect 14926 6196 14992 6230
rect 15026 6196 15092 6230
rect 15126 6196 15192 6230
rect 15226 6196 15292 6230
rect 15326 6196 15371 6230
rect 14761 6180 15371 6196
rect 17428 6281 17474 6319
rect 17428 6247 17434 6281
rect 17468 6247 17474 6281
rect 17428 6209 17474 6247
rect 13676 6166 13746 6170
rect -3658 5835 -3612 5873
rect -3658 5801 -3652 5835
rect -3618 5801 -3612 5835
rect -3658 5763 -3612 5801
rect -3658 5729 -3652 5763
rect -3618 5729 -3612 5763
rect -4174 5657 -4168 5691
rect -4134 5657 -4128 5691
rect -4174 5619 -4128 5657
rect -4174 5585 -4168 5619
rect -4134 5585 -4128 5619
rect -4174 5538 -4128 5585
rect -3916 5691 -3870 5693
rect -3916 5657 -3910 5691
rect -3876 5657 -3870 5691
rect -3916 5619 -3870 5657
rect -3916 5585 -3910 5619
rect -3876 5585 -3870 5619
rect -3916 5538 -3870 5585
rect -3658 5691 -3612 5729
rect -3488 5885 -3384 5901
rect -3488 5833 -3465 5885
rect -3413 5833 -3384 5885
rect -3488 5821 -3384 5833
rect -3488 5769 -3465 5821
rect -3413 5769 -3384 5821
rect -3488 5757 -3384 5769
rect -3488 5705 -3465 5757
rect -3413 5705 -3384 5757
rect -3488 5692 -3384 5705
rect -3658 5657 -3652 5691
rect -3618 5657 -3612 5691
rect -3658 5619 -3612 5657
rect -3658 5585 -3652 5619
rect -3618 5585 -3612 5619
rect -3658 5538 -3612 5585
rect -7786 5500 -7538 5506
rect -7786 5466 -7687 5500
rect -7653 5466 -7615 5500
rect -7581 5466 -7538 5500
rect -7786 5460 -7538 5466
rect -7472 5500 -7280 5506
rect -7472 5466 -7429 5500
rect -7395 5466 -7357 5500
rect -7323 5466 -7280 5500
rect -7472 5460 -7280 5466
rect -7214 5500 -7022 5506
rect -7214 5466 -7171 5500
rect -7137 5466 -7099 5500
rect -7065 5466 -7022 5500
rect -7214 5460 -7022 5466
rect -7786 5450 -7022 5460
rect -6956 5500 -6764 5506
rect -6956 5466 -6913 5500
rect -6879 5466 -6841 5500
rect -6807 5466 -6764 5500
rect -6956 5460 -6764 5466
rect -6698 5500 -6506 5506
rect -6698 5466 -6655 5500
rect -6621 5466 -6583 5500
rect -6549 5466 -6506 5500
rect -6698 5460 -6506 5466
rect -6440 5500 -6248 5506
rect -6440 5466 -6397 5500
rect -6363 5466 -6325 5500
rect -6291 5466 -6248 5500
rect -6440 5460 -6248 5466
rect -6182 5500 -5990 5506
rect -6182 5466 -6139 5500
rect -6105 5466 -6067 5500
rect -6033 5466 -5990 5500
rect -6182 5460 -5990 5466
rect -5924 5500 -5732 5506
rect -5924 5466 -5881 5500
rect -5847 5466 -5809 5500
rect -5775 5466 -5732 5500
rect -5924 5460 -5732 5466
rect -5666 5500 -5474 5506
rect -5666 5466 -5623 5500
rect -5589 5466 -5551 5500
rect -5517 5466 -5474 5500
rect -5666 5460 -5474 5466
rect -5408 5500 -5216 5506
rect -5408 5466 -5365 5500
rect -5331 5466 -5293 5500
rect -5259 5466 -5216 5500
rect -5408 5460 -5216 5466
rect -5150 5500 -4958 5506
rect -5150 5466 -5107 5500
rect -5073 5466 -5035 5500
rect -5001 5466 -4958 5500
rect -5150 5460 -4958 5466
rect -4892 5500 -4700 5506
rect -4892 5466 -4849 5500
rect -4815 5466 -4777 5500
rect -4743 5466 -4700 5500
rect -4892 5460 -4700 5466
rect -4634 5500 -4442 5506
rect -4634 5466 -4591 5500
rect -4557 5466 -4519 5500
rect -4485 5466 -4442 5500
rect -4634 5460 -4442 5466
rect -6956 5450 -4442 5460
rect -4376 5500 -4184 5506
rect -4376 5466 -4333 5500
rect -4299 5466 -4261 5500
rect -4227 5466 -4184 5500
rect -4376 5460 -4184 5466
rect -4118 5500 -3926 5506
rect -4118 5466 -4075 5500
rect -4041 5466 -4003 5500
rect -3969 5466 -3926 5500
rect -4118 5460 -3926 5466
rect -3860 5500 -3668 5506
rect -3860 5466 -3817 5500
rect -3783 5466 -3745 5500
rect -3711 5466 -3668 5500
rect -3860 5460 -3668 5466
rect -4376 5450 -3668 5460
rect -7786 5396 -3668 5450
rect 13066 5440 13746 6166
rect 14736 5562 15416 6180
rect 17428 6175 17434 6209
rect 17468 6175 17474 6209
rect 17428 6137 17474 6175
rect 17428 6103 17434 6137
rect 17468 6103 17474 6137
rect 17428 6065 17474 6103
rect 17428 6031 17434 6065
rect 17468 6031 17474 6065
rect 17428 5993 17474 6031
rect 17428 5959 17434 5993
rect 17468 5959 17474 5993
rect 17428 5921 17474 5959
rect 17428 5887 17434 5921
rect 17468 5887 17474 5921
rect 17428 5849 17474 5887
rect 17428 5815 17434 5849
rect 17468 5815 17474 5849
rect 17428 5777 17474 5815
rect 17428 5743 17434 5777
rect 17468 5743 17474 5777
rect 17428 5705 17474 5743
rect 17428 5671 17434 5705
rect 17468 5671 17474 5705
rect 17428 5633 17474 5671
rect 17428 5599 17434 5633
rect 17468 5599 17474 5633
rect 16482 5562 16658 5570
rect 14736 5440 16664 5562
rect 13066 5370 16664 5440
rect 13066 5350 14792 5370
rect 13066 5316 13142 5350
rect 13176 5316 13242 5350
rect 13276 5316 13342 5350
rect 13376 5316 13442 5350
rect 13476 5316 13542 5350
rect 13576 5316 13642 5350
rect 13676 5336 14792 5350
rect 14826 5336 14892 5370
rect 14926 5336 14992 5370
rect 15026 5336 15092 5370
rect 15126 5336 15192 5370
rect 15226 5336 15292 5370
rect 15326 5336 16664 5370
rect 13676 5316 16664 5336
rect 13066 5270 16664 5316
rect 13066 5250 14792 5270
rect 13066 5216 13142 5250
rect 13176 5216 13242 5250
rect 13276 5216 13342 5250
rect 13376 5216 13442 5250
rect 13476 5216 13542 5250
rect 13576 5216 13642 5250
rect 13676 5236 14792 5250
rect 14826 5236 14892 5270
rect 14926 5236 14992 5270
rect 15026 5236 15092 5270
rect 15126 5236 15192 5270
rect 15226 5236 15292 5270
rect 15326 5236 16664 5270
rect 13676 5216 16664 5236
rect 13066 5210 16664 5216
rect 13111 5208 16664 5210
rect 17428 5561 17474 5599
rect 17428 5527 17434 5561
rect 17468 5527 17474 5561
rect 17428 5489 17474 5527
rect 17428 5455 17434 5489
rect 17468 5455 17474 5489
rect 17428 5417 17474 5455
rect 17428 5383 17434 5417
rect 17468 5383 17474 5417
rect 17428 5345 17474 5383
rect 17428 5311 17434 5345
rect 17468 5311 17474 5345
rect 17428 5273 17474 5311
rect 17428 5239 17434 5273
rect 17468 5239 17474 5273
rect 13111 5170 15371 5208
rect 13111 5150 14792 5170
rect 13111 5116 13142 5150
rect 13176 5116 13242 5150
rect 13276 5116 13342 5150
rect 13376 5116 13442 5150
rect 13476 5116 13542 5150
rect 13576 5116 13642 5150
rect 13676 5136 14792 5150
rect 14826 5136 14892 5170
rect 14926 5136 14992 5170
rect 15026 5136 15092 5170
rect 15126 5136 15192 5170
rect 15226 5136 15292 5170
rect 15326 5136 15371 5170
rect 13676 5116 15371 5136
rect 13111 5070 15371 5116
rect 13111 5050 14792 5070
rect 13111 5016 13142 5050
rect 13176 5016 13242 5050
rect 13276 5016 13342 5050
rect 13376 5016 13442 5050
rect 13476 5016 13542 5050
rect 13576 5016 13642 5050
rect 13676 5036 14792 5050
rect 14826 5036 14892 5070
rect 14926 5036 14992 5070
rect 15026 5036 15092 5070
rect 15126 5036 15192 5070
rect 15226 5036 15292 5070
rect 15326 5036 15371 5070
rect 13676 5016 15371 5036
rect 13111 4970 15371 5016
rect 13111 4950 14792 4970
rect 13111 4916 13142 4950
rect 13176 4916 13242 4950
rect 13276 4916 13342 4950
rect 13376 4916 13442 4950
rect 13476 4916 13542 4950
rect 13576 4916 13642 4950
rect 13676 4936 14792 4950
rect 14826 4936 14892 4970
rect 14926 4936 14992 4970
rect 15026 4936 15092 4970
rect 15126 4936 15192 4970
rect 15226 4936 15292 4970
rect 15326 4936 15371 4970
rect 13676 4916 15371 4936
rect 13111 4870 15371 4916
rect 13111 4850 14792 4870
rect 13111 4816 13142 4850
rect 13176 4816 13242 4850
rect 13276 4816 13342 4850
rect 13376 4816 13442 4850
rect 13476 4816 13542 4850
rect 13576 4816 13642 4850
rect 13676 4836 14792 4850
rect 14826 4836 14892 4870
rect 14926 4836 14992 4870
rect 15026 4836 15092 4870
rect 15126 4836 15192 4870
rect 15226 4836 15292 4870
rect 15326 4836 15371 4870
rect 13676 4816 15371 4836
rect 13111 4805 15371 4816
rect 16220 5059 16270 5073
rect 16220 5025 16228 5059
rect 16262 5025 16270 5059
rect 16220 4987 16270 5025
rect 16220 4953 16228 4987
rect 16262 4953 16270 4987
rect 16220 4915 16270 4953
rect 16220 4881 16228 4915
rect 16262 4881 16270 4915
rect 16220 4843 16270 4881
rect 16220 4809 16228 4843
rect 16262 4809 16270 4843
rect 13111 4785 14816 4805
rect 13586 4750 14816 4785
rect 16220 4771 16270 4809
rect 16220 4737 16228 4771
rect 16262 4737 16270 4771
rect 16220 4699 16270 4737
rect 16220 4665 16228 4699
rect 16262 4665 16270 4699
rect 16220 4652 16270 4665
rect 16482 5066 16658 5208
rect 17428 5201 17474 5239
rect 17428 5167 17434 5201
rect 17468 5167 17474 5201
rect 17428 5129 17474 5167
rect 17428 5095 17434 5129
rect 17468 5095 17474 5129
rect 16482 5059 16778 5066
rect 16482 5025 16546 5059
rect 16580 5025 16778 5059
rect 16482 4987 16778 5025
rect 16482 4953 16546 4987
rect 16580 4953 16778 4987
rect 16482 4915 16778 4953
rect 16482 4881 16546 4915
rect 16580 4881 16778 4915
rect 16482 4843 16778 4881
rect 16482 4809 16546 4843
rect 16580 4809 16778 4843
rect 16482 4771 16778 4809
rect 16482 4737 16546 4771
rect 16580 4737 16778 4771
rect 16482 4699 16778 4737
rect 16482 4665 16546 4699
rect 16580 4665 16778 4699
rect 16482 4642 16778 4665
rect 16856 5059 16906 5073
rect 16856 5025 16864 5059
rect 16898 5025 16906 5059
rect 16856 4987 16906 5025
rect 16856 4953 16864 4987
rect 16898 4953 16906 4987
rect 16856 4915 16906 4953
rect 16856 4881 16864 4915
rect 16898 4881 16906 4915
rect 16856 4843 16906 4881
rect 16856 4809 16864 4843
rect 16898 4809 16906 4843
rect 16856 4771 16906 4809
rect 16856 4737 16864 4771
rect 16898 4737 16906 4771
rect 16856 4699 16906 4737
rect 16856 4665 16864 4699
rect 16898 4665 16906 4699
rect 16856 4652 16906 4665
rect 17428 5057 17474 5095
rect 17428 5023 17434 5057
rect 17468 5023 17474 5057
rect 17428 4985 17474 5023
rect 17428 4951 17434 4985
rect 17468 4951 17474 4985
rect 17428 4913 17474 4951
rect 17428 4879 17434 4913
rect 17468 4879 17474 4913
rect 17428 4841 17474 4879
rect 17428 4807 17434 4841
rect 17468 4807 17474 4841
rect 17428 4769 17474 4807
rect 17428 4735 17434 4769
rect 17468 4735 17474 4769
rect 17428 4697 17474 4735
rect 17428 4663 17434 4697
rect 17468 4663 17474 4697
rect 16482 4640 16658 4642
rect 16706 4628 16776 4642
rect 17428 4625 17474 4663
rect 17428 4591 17434 4625
rect 17468 4591 17474 4625
rect 17428 4548 17474 4591
rect 18486 6929 18532 6967
rect 18486 6895 18492 6929
rect 18526 6895 18532 6929
rect 18486 6857 18532 6895
rect 18486 6823 18492 6857
rect 18526 6823 18532 6857
rect 18486 6785 18532 6823
rect 18486 6751 18492 6785
rect 18526 6751 18532 6785
rect 18486 6713 18532 6751
rect 18486 6679 18492 6713
rect 18526 6679 18532 6713
rect 18486 6641 18532 6679
rect 18486 6607 18492 6641
rect 18526 6607 18532 6641
rect 18486 6569 18532 6607
rect 18878 7505 18924 7548
rect 19936 7510 19982 7548
rect 20012 7510 20152 7770
rect 23532 7783 23578 7830
rect 23532 7749 23538 7783
rect 23572 7749 23578 7783
rect 23642 7821 23664 7840
rect 23716 7821 23728 7846
rect 23780 7840 24610 7846
rect 25110 7880 26110 7886
rect 25110 7846 25125 7880
rect 25159 7863 25197 7880
rect 25231 7863 25269 7880
rect 25159 7846 25164 7863
rect 25303 7846 25341 7880
rect 25375 7846 25413 7880
rect 25447 7846 25485 7880
rect 25519 7846 25557 7880
rect 25591 7846 25629 7880
rect 25663 7846 25701 7880
rect 25735 7846 25773 7880
rect 25807 7846 25845 7880
rect 25879 7846 25917 7880
rect 25951 7846 25989 7880
rect 26023 7846 26061 7880
rect 26095 7846 26110 7880
rect 25110 7840 25164 7846
rect 23780 7821 23812 7840
rect 23642 7782 23812 7821
rect 24642 7783 24688 7830
rect 23532 7711 23578 7749
rect 23532 7682 23538 7711
rect 18878 7471 18884 7505
rect 18918 7471 18924 7505
rect 18878 7433 18924 7471
rect 18878 7399 18884 7433
rect 18918 7399 18924 7433
rect 18878 7361 18924 7399
rect 19922 7505 20152 7510
rect 19922 7471 19942 7505
rect 19976 7471 20152 7505
rect 19922 7433 20152 7471
rect 19922 7399 19942 7433
rect 19976 7399 20152 7433
rect 19922 7370 20152 7399
rect 21862 7677 23538 7682
rect 23572 7677 23578 7711
rect 21862 7639 23578 7677
rect 21862 7631 23538 7639
rect 18878 7327 18884 7361
rect 18918 7327 18924 7361
rect 18878 7289 18924 7327
rect 18878 7255 18884 7289
rect 18918 7255 18924 7289
rect 18878 7217 18924 7255
rect 18878 7183 18884 7217
rect 18918 7183 18924 7217
rect 18878 7145 18924 7183
rect 18878 7111 18884 7145
rect 18918 7111 18924 7145
rect 18878 7073 18924 7111
rect 18878 7039 18884 7073
rect 18918 7039 18924 7073
rect 18878 7001 18924 7039
rect 18878 6967 18884 7001
rect 18918 6967 18924 7001
rect 18878 6929 18924 6967
rect 18878 6895 18884 6929
rect 18918 6895 18924 6929
rect 18878 6857 18924 6895
rect 18878 6823 18884 6857
rect 18918 6823 18924 6857
rect 18878 6785 18924 6823
rect 18878 6751 18884 6785
rect 18918 6751 18924 6785
rect 18878 6713 18924 6751
rect 18878 6679 18884 6713
rect 18918 6679 18924 6713
rect 18878 6641 18924 6679
rect 18878 6607 18884 6641
rect 18918 6607 18924 6641
rect 18878 6600 18924 6607
rect 19936 7361 19982 7370
rect 19936 7327 19942 7361
rect 19976 7327 19982 7361
rect 19936 7289 19982 7327
rect 19936 7255 19942 7289
rect 19976 7255 19982 7289
rect 19936 7217 19982 7255
rect 19936 7183 19942 7217
rect 19976 7183 19982 7217
rect 19936 7145 19982 7183
rect 19936 7111 19942 7145
rect 19976 7111 19982 7145
rect 19936 7073 19982 7111
rect 19936 7039 19942 7073
rect 19976 7039 19982 7073
rect 21862 7093 21898 7631
rect 22436 7605 23538 7631
rect 23572 7605 23578 7639
rect 22436 7567 23578 7605
rect 22436 7533 23538 7567
rect 23572 7533 23578 7567
rect 22436 7495 23578 7533
rect 22436 7461 23538 7495
rect 23572 7461 23578 7495
rect 22436 7423 23578 7461
rect 22436 7389 23538 7423
rect 23572 7389 23578 7423
rect 22436 7351 23578 7389
rect 22436 7317 23538 7351
rect 23572 7317 23578 7351
rect 22436 7279 23578 7317
rect 22436 7245 23538 7279
rect 23572 7245 23578 7279
rect 22436 7207 23578 7245
rect 22436 7173 23538 7207
rect 23572 7173 23578 7207
rect 22436 7135 23578 7173
rect 22436 7101 23538 7135
rect 23572 7101 23578 7135
rect 22436 7093 23578 7101
rect 21862 7063 23578 7093
rect 21862 7062 23538 7063
rect 19936 7001 19982 7039
rect 19936 6967 19942 7001
rect 19976 6967 19982 7001
rect 19936 6929 19982 6967
rect 19936 6895 19942 6929
rect 19976 6895 19982 6929
rect 23532 7029 23538 7062
rect 23572 7029 23578 7063
rect 23532 6991 23578 7029
rect 23532 6957 23538 6991
rect 23572 6957 23578 6991
rect 23532 6919 23578 6957
rect 23532 6902 23538 6919
rect 19936 6857 19982 6895
rect 19936 6823 19942 6857
rect 19976 6823 19982 6857
rect 19936 6785 19982 6823
rect 19936 6751 19942 6785
rect 19976 6751 19982 6785
rect 19936 6713 19982 6751
rect 19936 6679 19942 6713
rect 19976 6679 19982 6713
rect 23502 6885 23538 6902
rect 23572 6885 23578 6919
rect 23502 6838 23578 6885
rect 24642 7749 24648 7783
rect 24682 7749 24688 7783
rect 24642 7711 24688 7749
rect 24642 7677 24648 7711
rect 24682 7677 24688 7711
rect 24642 7639 24688 7677
rect 24642 7605 24648 7639
rect 24682 7605 24688 7639
rect 24642 7567 24688 7605
rect 24642 7533 24648 7567
rect 24682 7533 24688 7567
rect 24642 7495 24688 7533
rect 24642 7461 24648 7495
rect 24682 7461 24688 7495
rect 24642 7423 24688 7461
rect 24642 7389 24648 7423
rect 24682 7389 24688 7423
rect 24642 7351 24688 7389
rect 24642 7317 24648 7351
rect 24682 7317 24688 7351
rect 24642 7279 24688 7317
rect 24642 7245 24648 7279
rect 24682 7245 24688 7279
rect 24642 7207 24688 7245
rect 24642 7173 24648 7207
rect 24682 7173 24688 7207
rect 24642 7135 24688 7173
rect 24642 7101 24648 7135
rect 24682 7101 24688 7135
rect 24642 7063 24688 7101
rect 24642 7029 24648 7063
rect 24682 7029 24688 7063
rect 24642 6991 24688 7029
rect 24642 6957 24648 6991
rect 24682 6957 24688 6991
rect 24642 6919 24688 6957
rect 24642 6885 24648 6919
rect 24682 6892 24688 6919
rect 25032 7783 25078 7830
rect 25032 7749 25038 7783
rect 25072 7749 25078 7783
rect 25142 7811 25164 7840
rect 25216 7811 25228 7846
rect 25280 7840 26110 7846
rect 25280 7811 25302 7840
rect 26182 7830 26222 8162
rect 25142 7782 25302 7811
rect 26142 7783 26222 7830
rect 25032 7711 25078 7749
rect 25032 7677 25038 7711
rect 25072 7677 25078 7711
rect 25032 7639 25078 7677
rect 25032 7605 25038 7639
rect 25072 7605 25078 7639
rect 25032 7567 25078 7605
rect 25032 7533 25038 7567
rect 25072 7533 25078 7567
rect 25032 7495 25078 7533
rect 25032 7461 25038 7495
rect 25072 7461 25078 7495
rect 25032 7423 25078 7461
rect 25032 7389 25038 7423
rect 25072 7389 25078 7423
rect 25032 7351 25078 7389
rect 25032 7317 25038 7351
rect 25072 7317 25078 7351
rect 25032 7279 25078 7317
rect 25032 7245 25038 7279
rect 25072 7245 25078 7279
rect 25032 7207 25078 7245
rect 25032 7173 25038 7207
rect 25072 7173 25078 7207
rect 25032 7135 25078 7173
rect 25032 7101 25038 7135
rect 25072 7101 25078 7135
rect 25032 7063 25078 7101
rect 25032 7029 25038 7063
rect 25072 7029 25078 7063
rect 25032 6991 25078 7029
rect 25032 6957 25038 6991
rect 25072 6957 25078 6991
rect 25032 6919 25078 6957
rect 26142 7749 26148 7783
rect 26182 7749 26222 7783
rect 26142 7711 26222 7749
rect 26142 7677 26148 7711
rect 26182 7677 26222 7711
rect 26142 7639 26222 7677
rect 26142 7605 26148 7639
rect 26182 7605 26222 7639
rect 26142 7567 26222 7605
rect 26142 7533 26148 7567
rect 26182 7533 26222 7567
rect 26142 7495 26222 7533
rect 26142 7461 26148 7495
rect 26182 7479 26222 7495
rect 26338 7479 26382 8427
rect 37730 8450 37814 9549
rect 38064 9517 38110 9564
rect 38272 9708 38278 9729
rect 38312 9729 38335 9742
rect 38530 9886 38576 9924
rect 38788 10068 38794 10102
rect 38828 10068 38834 10102
rect 39027 10225 39052 10245
rect 39086 10245 39092 10246
rect 39304 10534 39350 10549
rect 39304 10500 39310 10534
rect 39344 10500 39350 10534
rect 39304 10462 39350 10500
rect 39304 10428 39310 10462
rect 39344 10428 39350 10462
rect 39304 10390 39350 10428
rect 39304 10356 39310 10390
rect 39344 10356 39350 10390
rect 39304 10318 39350 10356
rect 39304 10284 39310 10318
rect 39344 10284 39350 10318
rect 39304 10246 39350 10284
rect 39086 10225 39111 10245
rect 39027 10173 39043 10225
rect 39095 10173 39111 10225
rect 39027 10161 39052 10173
rect 39086 10161 39111 10173
rect 39027 10109 39043 10161
rect 39095 10109 39111 10161
rect 39027 10102 39111 10109
rect 39027 10093 39052 10102
rect 38788 10030 38834 10068
rect 38788 9996 38794 10030
rect 38828 9996 38834 10030
rect 38788 9958 38834 9996
rect 38788 9924 38794 9958
rect 38828 9924 38834 9958
rect 38788 9914 38834 9924
rect 39046 10068 39052 10093
rect 39086 10093 39111 10102
rect 39304 10212 39310 10246
rect 39344 10212 39350 10246
rect 39562 10534 39608 10549
rect 39562 10500 39568 10534
rect 39602 10500 39608 10534
rect 39562 10462 39608 10500
rect 39562 10428 39568 10462
rect 39602 10428 39608 10462
rect 39562 10390 39608 10428
rect 39562 10356 39568 10390
rect 39602 10356 39608 10390
rect 39562 10318 39608 10356
rect 39562 10284 39568 10318
rect 39602 10284 39608 10318
rect 39562 10246 39608 10284
rect 39562 10245 39568 10246
rect 39304 10174 39350 10212
rect 39304 10140 39310 10174
rect 39344 10140 39350 10174
rect 39304 10102 39350 10140
rect 39086 10068 39092 10093
rect 39046 10030 39092 10068
rect 39046 9996 39052 10030
rect 39086 9996 39092 10030
rect 39046 9958 39092 9996
rect 39046 9924 39052 9958
rect 39086 9924 39092 9958
rect 38530 9852 38536 9886
rect 38570 9852 38576 9886
rect 38530 9814 38576 9852
rect 38530 9780 38536 9814
rect 38570 9780 38576 9814
rect 38530 9742 38576 9780
rect 38312 9708 38318 9729
rect 38272 9670 38318 9708
rect 38272 9636 38278 9670
rect 38312 9636 38318 9670
rect 38272 9598 38318 9636
rect 38272 9564 38278 9598
rect 38312 9564 38318 9598
rect 38272 9549 38318 9564
rect 38530 9708 38536 9742
rect 38570 9708 38576 9742
rect 38771 9886 38855 9914
rect 38771 9877 38794 9886
rect 38828 9877 38855 9886
rect 38771 9825 38787 9877
rect 38839 9825 38855 9877
rect 38771 9814 38855 9825
rect 38771 9813 38794 9814
rect 38828 9813 38855 9814
rect 38771 9761 38787 9813
rect 38839 9761 38855 9813
rect 38771 9742 38855 9761
rect 38771 9729 38794 9742
rect 38530 9670 38576 9708
rect 38530 9636 38536 9670
rect 38570 9636 38576 9670
rect 38530 9598 38576 9636
rect 38530 9564 38536 9598
rect 38570 9564 38576 9598
rect 38530 9549 38576 9564
rect 38788 9708 38794 9729
rect 38828 9729 38855 9742
rect 39046 9886 39092 9924
rect 39304 10068 39310 10102
rect 39344 10068 39350 10102
rect 39542 10227 39568 10245
rect 39602 10245 39608 10246
rect 39820 10534 39866 10549
rect 39820 10500 39826 10534
rect 39860 10500 39866 10534
rect 39820 10462 39866 10500
rect 39820 10428 39826 10462
rect 39860 10428 39866 10462
rect 39820 10390 39866 10428
rect 39820 10356 39826 10390
rect 39860 10356 39866 10390
rect 39820 10318 39866 10356
rect 39820 10284 39826 10318
rect 39860 10284 39866 10318
rect 39820 10246 39866 10284
rect 39602 10227 39630 10245
rect 39542 10175 39559 10227
rect 39611 10175 39630 10227
rect 39542 10174 39630 10175
rect 39542 10163 39568 10174
rect 39602 10163 39630 10174
rect 39542 10111 39559 10163
rect 39611 10111 39630 10163
rect 39542 10102 39630 10111
rect 39542 10093 39568 10102
rect 39304 10030 39350 10068
rect 39304 9996 39310 10030
rect 39344 9996 39350 10030
rect 39304 9958 39350 9996
rect 39304 9924 39310 9958
rect 39344 9924 39350 9958
rect 39304 9914 39350 9924
rect 39562 10068 39568 10093
rect 39602 10093 39630 10102
rect 39820 10212 39826 10246
rect 39860 10212 39866 10246
rect 40078 10534 40124 10549
rect 40078 10500 40084 10534
rect 40118 10500 40124 10534
rect 40078 10462 40124 10500
rect 40078 10428 40084 10462
rect 40118 10428 40124 10462
rect 40078 10390 40124 10428
rect 40078 10356 40084 10390
rect 40118 10356 40124 10390
rect 40078 10318 40124 10356
rect 40078 10284 40084 10318
rect 40118 10284 40124 10318
rect 40078 10246 40124 10284
rect 40078 10245 40084 10246
rect 39820 10174 39866 10212
rect 39820 10140 39826 10174
rect 39860 10140 39866 10174
rect 39820 10102 39866 10140
rect 39602 10068 39608 10093
rect 39562 10030 39608 10068
rect 39562 9996 39568 10030
rect 39602 9996 39608 10030
rect 39562 9958 39608 9996
rect 39562 9924 39568 9958
rect 39602 9924 39608 9958
rect 39046 9852 39052 9886
rect 39086 9852 39092 9886
rect 39046 9814 39092 9852
rect 39046 9780 39052 9814
rect 39086 9780 39092 9814
rect 39046 9742 39092 9780
rect 38828 9708 38834 9729
rect 38788 9670 38834 9708
rect 38788 9636 38794 9670
rect 38828 9636 38834 9670
rect 38788 9598 38834 9636
rect 38788 9564 38794 9598
rect 38828 9564 38834 9598
rect 38788 9549 38834 9564
rect 39046 9708 39052 9742
rect 39086 9708 39092 9742
rect 39284 9886 39369 9914
rect 39284 9879 39310 9886
rect 39344 9879 39369 9886
rect 39284 9827 39300 9879
rect 39352 9827 39369 9879
rect 39284 9815 39369 9827
rect 39284 9763 39300 9815
rect 39352 9763 39369 9815
rect 39284 9742 39369 9763
rect 39284 9729 39310 9742
rect 39046 9670 39092 9708
rect 39046 9636 39052 9670
rect 39086 9636 39092 9670
rect 39046 9598 39092 9636
rect 39046 9564 39052 9598
rect 39086 9564 39092 9598
rect 39046 9549 39092 9564
rect 39304 9708 39310 9729
rect 39344 9729 39369 9742
rect 39562 9886 39608 9924
rect 39820 10068 39826 10102
rect 39860 10068 39866 10102
rect 40061 10225 40084 10245
rect 40118 10245 40124 10246
rect 40336 10534 40382 10549
rect 40336 10500 40342 10534
rect 40376 10500 40382 10534
rect 40336 10462 40382 10500
rect 40336 10428 40342 10462
rect 40376 10428 40382 10462
rect 40336 10390 40382 10428
rect 40336 10356 40342 10390
rect 40376 10356 40382 10390
rect 40336 10318 40382 10356
rect 40336 10284 40342 10318
rect 40376 10284 40382 10318
rect 40336 10246 40382 10284
rect 40118 10225 40143 10245
rect 40061 10173 40076 10225
rect 40128 10173 40143 10225
rect 40061 10161 40084 10173
rect 40118 10161 40143 10173
rect 40061 10109 40076 10161
rect 40128 10109 40143 10161
rect 40061 10102 40143 10109
rect 40061 10093 40084 10102
rect 39820 10030 39866 10068
rect 39820 9996 39826 10030
rect 39860 9996 39866 10030
rect 39820 9958 39866 9996
rect 39820 9924 39826 9958
rect 39860 9924 39866 9958
rect 39820 9914 39866 9924
rect 40078 10068 40084 10093
rect 40118 10093 40143 10102
rect 40336 10212 40342 10246
rect 40376 10212 40382 10246
rect 40594 10534 40640 10549
rect 40594 10500 40600 10534
rect 40634 10500 40640 10534
rect 40594 10462 40640 10500
rect 40594 10428 40600 10462
rect 40634 10428 40640 10462
rect 40594 10390 40640 10428
rect 40594 10356 40600 10390
rect 40634 10356 40640 10390
rect 40594 10318 40640 10356
rect 40594 10284 40600 10318
rect 40634 10284 40640 10318
rect 40594 10246 40640 10284
rect 40594 10245 40600 10246
rect 40336 10174 40382 10212
rect 40336 10140 40342 10174
rect 40376 10140 40382 10174
rect 40336 10102 40382 10140
rect 40118 10068 40124 10093
rect 40078 10030 40124 10068
rect 40078 9996 40084 10030
rect 40118 9996 40124 10030
rect 40078 9958 40124 9996
rect 40078 9924 40084 9958
rect 40118 9924 40124 9958
rect 39562 9852 39568 9886
rect 39602 9852 39608 9886
rect 39562 9814 39608 9852
rect 39562 9780 39568 9814
rect 39602 9780 39608 9814
rect 39562 9742 39608 9780
rect 39344 9708 39350 9729
rect 39304 9670 39350 9708
rect 39304 9636 39310 9670
rect 39344 9636 39350 9670
rect 39304 9598 39350 9636
rect 39304 9564 39310 9598
rect 39344 9564 39350 9598
rect 39304 9549 39350 9564
rect 39562 9708 39568 9742
rect 39602 9708 39608 9742
rect 39803 9886 39886 9914
rect 39803 9878 39826 9886
rect 39860 9878 39886 9886
rect 39803 9826 39818 9878
rect 39870 9826 39886 9878
rect 39803 9814 39886 9826
rect 39803 9762 39818 9814
rect 39870 9762 39886 9814
rect 39803 9742 39886 9762
rect 39803 9729 39826 9742
rect 39562 9670 39608 9708
rect 39562 9636 39568 9670
rect 39602 9636 39608 9670
rect 39562 9598 39608 9636
rect 39562 9564 39568 9598
rect 39602 9564 39608 9598
rect 39562 9549 39608 9564
rect 39820 9708 39826 9729
rect 39860 9729 39886 9742
rect 40078 9886 40124 9924
rect 40336 10068 40342 10102
rect 40376 10068 40382 10102
rect 40575 10226 40600 10245
rect 40634 10245 40640 10246
rect 40852 10534 40898 10549
rect 40852 10500 40858 10534
rect 40892 10500 40898 10534
rect 40852 10462 40898 10500
rect 40852 10428 40858 10462
rect 40892 10428 40898 10462
rect 40852 10390 40898 10428
rect 40852 10356 40858 10390
rect 40892 10356 40898 10390
rect 40852 10318 40898 10356
rect 40852 10284 40858 10318
rect 40892 10284 40898 10318
rect 40852 10246 40898 10284
rect 40634 10226 40662 10245
rect 40575 10174 40590 10226
rect 40642 10174 40662 10226
rect 40575 10162 40600 10174
rect 40634 10162 40662 10174
rect 40575 10110 40590 10162
rect 40642 10110 40662 10162
rect 40575 10102 40662 10110
rect 40575 10093 40600 10102
rect 40336 10030 40382 10068
rect 40336 9996 40342 10030
rect 40376 9996 40382 10030
rect 40336 9958 40382 9996
rect 40336 9924 40342 9958
rect 40376 9924 40382 9958
rect 40336 9914 40382 9924
rect 40594 10068 40600 10093
rect 40634 10093 40662 10102
rect 40852 10212 40858 10246
rect 40892 10212 40898 10246
rect 40852 10174 40898 10212
rect 40852 10140 40858 10174
rect 40892 10140 40898 10174
rect 40852 10102 40898 10140
rect 40634 10068 40640 10093
rect 40594 10030 40640 10068
rect 40594 9996 40600 10030
rect 40634 9996 40640 10030
rect 40594 9958 40640 9996
rect 40594 9924 40600 9958
rect 40634 9924 40640 9958
rect 40078 9852 40084 9886
rect 40118 9852 40124 9886
rect 40078 9814 40124 9852
rect 40078 9780 40084 9814
rect 40118 9780 40124 9814
rect 40078 9742 40124 9780
rect 39860 9708 39866 9729
rect 39820 9670 39866 9708
rect 39820 9636 39826 9670
rect 39860 9636 39866 9670
rect 39820 9598 39866 9636
rect 39820 9564 39826 9598
rect 39860 9564 39866 9598
rect 39820 9549 39866 9564
rect 40078 9708 40084 9742
rect 40118 9708 40124 9742
rect 40315 9886 40406 9914
rect 40315 9878 40342 9886
rect 40376 9878 40406 9886
rect 40315 9826 40335 9878
rect 40387 9826 40406 9878
rect 40315 9814 40406 9826
rect 40315 9762 40335 9814
rect 40387 9762 40406 9814
rect 40315 9742 40406 9762
rect 40315 9729 40342 9742
rect 40078 9670 40124 9708
rect 40078 9636 40084 9670
rect 40118 9636 40124 9670
rect 40078 9598 40124 9636
rect 40078 9564 40084 9598
rect 40118 9564 40124 9598
rect 40078 9549 40124 9564
rect 40336 9708 40342 9729
rect 40376 9729 40406 9742
rect 40594 9886 40640 9924
rect 40852 10068 40858 10102
rect 40892 10068 40898 10102
rect 40852 10030 40898 10068
rect 40852 9996 40858 10030
rect 40892 9996 40898 10030
rect 40852 9958 40898 9996
rect 40852 9924 40858 9958
rect 40892 9924 40898 9958
rect 40852 9914 40898 9924
rect 40594 9852 40600 9886
rect 40634 9852 40640 9886
rect 40594 9814 40640 9852
rect 40594 9780 40600 9814
rect 40634 9780 40640 9814
rect 40594 9742 40640 9780
rect 40376 9708 40382 9729
rect 40336 9670 40382 9708
rect 40336 9636 40342 9670
rect 40376 9636 40382 9670
rect 40336 9598 40382 9636
rect 40336 9564 40342 9598
rect 40376 9564 40382 9598
rect 40336 9549 40382 9564
rect 40594 9708 40600 9742
rect 40634 9708 40640 9742
rect 40831 9886 40919 9914
rect 40831 9879 40858 9886
rect 40892 9879 40919 9886
rect 40831 9827 40850 9879
rect 40902 9827 40919 9879
rect 40831 9815 40919 9827
rect 40831 9763 40850 9815
rect 40902 9763 40919 9815
rect 40831 9742 40919 9763
rect 40831 9728 40858 9742
rect 40594 9670 40640 9708
rect 40594 9636 40600 9670
rect 40634 9636 40640 9670
rect 40594 9598 40640 9636
rect 40594 9564 40600 9598
rect 40634 9564 40640 9598
rect 40594 9549 40640 9564
rect 40852 9708 40858 9728
rect 40892 9728 40919 9742
rect 43358 9815 44648 9970
rect 40892 9708 40898 9728
rect 40852 9670 40898 9708
rect 40852 9636 40858 9670
rect 40892 9636 40898 9670
rect 40852 9598 40898 9636
rect 40852 9564 40858 9598
rect 40892 9564 40898 9598
rect 40852 9549 40898 9564
rect 37862 9511 38110 9517
rect 37862 9477 37905 9511
rect 37939 9477 37977 9511
rect 38011 9477 38110 9511
rect 37862 9471 38110 9477
rect 38328 9511 38520 9517
rect 38328 9477 38371 9511
rect 38405 9477 38443 9511
rect 38477 9477 38520 9511
rect 38328 9471 38520 9477
rect 38586 9511 38778 9517
rect 38586 9477 38629 9511
rect 38663 9477 38701 9511
rect 38735 9477 38778 9511
rect 38586 9471 38778 9477
rect 38844 9511 39036 9517
rect 38844 9477 38887 9511
rect 38921 9477 38959 9511
rect 38993 9477 39036 9511
rect 38844 9471 39036 9477
rect 39102 9511 39294 9517
rect 39102 9477 39145 9511
rect 39179 9477 39217 9511
rect 39251 9477 39294 9511
rect 39102 9471 39294 9477
rect 39360 9511 39552 9517
rect 39360 9477 39403 9511
rect 39437 9477 39475 9511
rect 39509 9477 39552 9511
rect 39360 9471 39552 9477
rect 39618 9511 39810 9517
rect 39618 9477 39661 9511
rect 39695 9477 39733 9511
rect 39767 9477 39810 9511
rect 39618 9471 39810 9477
rect 39876 9511 40068 9517
rect 39876 9477 39919 9511
rect 39953 9477 39991 9511
rect 40025 9477 40068 9511
rect 39876 9471 40068 9477
rect 40134 9511 40326 9517
rect 40134 9477 40177 9511
rect 40211 9477 40249 9511
rect 40283 9477 40326 9511
rect 40134 9471 40326 9477
rect 40392 9511 40584 9517
rect 40392 9477 40435 9511
rect 40469 9477 40507 9511
rect 40541 9477 40584 9511
rect 40392 9471 40584 9477
rect 40650 9511 40842 9517
rect 40650 9477 40693 9511
rect 40727 9477 40765 9511
rect 40799 9477 40842 9511
rect 40650 9471 40842 9477
rect 37862 9408 40842 9471
rect 37730 8376 41924 8450
rect 37730 8360 38054 8376
rect 37730 8326 37905 8360
rect 37939 8326 37977 8360
rect 38011 8326 38054 8360
rect 37730 8320 38054 8326
rect 38120 8360 38312 8376
rect 38120 8326 38163 8360
rect 38197 8326 38235 8360
rect 38269 8326 38312 8360
rect 38120 8320 38312 8326
rect 38378 8360 38570 8376
rect 38378 8326 38421 8360
rect 38455 8326 38493 8360
rect 38527 8326 38570 8360
rect 38378 8320 38570 8326
rect 38636 8366 41150 8376
rect 38636 8360 38828 8366
rect 38636 8326 38679 8360
rect 38713 8326 38751 8360
rect 38785 8326 38828 8360
rect 38636 8320 38828 8326
rect 38894 8360 39086 8366
rect 38894 8326 38937 8360
rect 38971 8326 39009 8360
rect 39043 8326 39086 8360
rect 38894 8320 39086 8326
rect 39152 8360 39344 8366
rect 39152 8326 39195 8360
rect 39229 8326 39267 8360
rect 39301 8326 39344 8360
rect 39152 8320 39344 8326
rect 39410 8360 39602 8366
rect 39410 8326 39453 8360
rect 39487 8326 39525 8360
rect 39559 8326 39602 8360
rect 39410 8320 39602 8326
rect 39668 8360 39860 8366
rect 39668 8326 39711 8360
rect 39745 8326 39783 8360
rect 39817 8326 39860 8360
rect 39668 8320 39860 8326
rect 39926 8360 40118 8366
rect 39926 8326 39969 8360
rect 40003 8326 40041 8360
rect 40075 8326 40118 8360
rect 39926 8320 40118 8326
rect 40184 8360 40376 8366
rect 40184 8326 40227 8360
rect 40261 8326 40299 8360
rect 40333 8326 40376 8360
rect 40184 8320 40376 8326
rect 40442 8360 40634 8366
rect 40442 8326 40485 8360
rect 40519 8326 40557 8360
rect 40591 8326 40634 8360
rect 40442 8320 40634 8326
rect 40700 8360 40892 8366
rect 40700 8326 40743 8360
rect 40777 8326 40815 8360
rect 40849 8326 40892 8360
rect 40700 8320 40892 8326
rect 40958 8360 41150 8366
rect 40958 8326 41001 8360
rect 41035 8326 41073 8360
rect 41107 8326 41150 8360
rect 40958 8320 41150 8326
rect 41216 8360 41408 8376
rect 41216 8326 41259 8360
rect 41293 8326 41331 8360
rect 41365 8326 41408 8360
rect 41216 8320 41408 8326
rect 41474 8360 41666 8376
rect 41474 8326 41517 8360
rect 41551 8326 41589 8360
rect 41623 8326 41666 8360
rect 41474 8320 41666 8326
rect 41732 8360 41924 8376
rect 41732 8326 41775 8360
rect 41809 8326 41847 8360
rect 41881 8326 41924 8360
rect 41732 8320 41924 8326
rect 37730 8241 37852 8320
rect 37730 8207 37812 8241
rect 37846 8207 37852 8241
rect 37730 8169 37852 8207
rect 37730 8135 37812 8169
rect 37846 8135 37852 8169
rect 37730 8113 37852 8135
rect 26182 7461 26382 7479
rect 26142 7452 26382 7461
rect 37806 8097 37852 8113
rect 37806 8063 37812 8097
rect 37846 8063 37852 8097
rect 37806 8025 37852 8063
rect 37806 7991 37812 8025
rect 37846 7991 37852 8025
rect 37806 7953 37852 7991
rect 37806 7919 37812 7953
rect 37846 7919 37852 7953
rect 37806 7881 37852 7919
rect 37806 7847 37812 7881
rect 37846 7847 37852 7881
rect 37806 7809 37852 7847
rect 37806 7775 37812 7809
rect 37846 7775 37852 7809
rect 37806 7737 37852 7775
rect 37806 7703 37812 7737
rect 37846 7703 37852 7737
rect 37806 7665 37852 7703
rect 37806 7631 37812 7665
rect 37846 7631 37852 7665
rect 37806 7593 37852 7631
rect 37806 7559 37812 7593
rect 37846 7559 37852 7593
rect 37806 7521 37852 7559
rect 37806 7487 37812 7521
rect 37846 7487 37852 7521
rect 26142 7423 26188 7452
rect 26142 7389 26148 7423
rect 26182 7389 26188 7423
rect 26142 7351 26188 7389
rect 26142 7317 26148 7351
rect 26182 7317 26188 7351
rect 26142 7279 26188 7317
rect 26142 7245 26148 7279
rect 26182 7245 26188 7279
rect 26142 7207 26188 7245
rect 26142 7173 26148 7207
rect 26182 7173 26188 7207
rect 26142 7135 26188 7173
rect 26142 7101 26148 7135
rect 26182 7101 26188 7135
rect 26142 7063 26188 7101
rect 26142 7029 26148 7063
rect 26182 7029 26188 7063
rect 26142 6991 26188 7029
rect 26142 6957 26148 6991
rect 26182 6957 26188 6991
rect 25032 6892 25038 6919
rect 24682 6885 24712 6892
rect 24642 6838 24712 6885
rect 23502 6772 23532 6838
rect 24362 6828 24522 6832
rect 23610 6822 24610 6828
rect 23610 6788 23625 6822
rect 23659 6788 23697 6822
rect 23731 6788 23769 6822
rect 23803 6788 23841 6822
rect 23875 6788 23913 6822
rect 23947 6788 23985 6822
rect 24019 6788 24057 6822
rect 24091 6788 24129 6822
rect 24163 6788 24201 6822
rect 24235 6788 24273 6822
rect 24307 6788 24345 6822
rect 24379 6808 24417 6822
rect 24451 6808 24489 6822
rect 24379 6788 24384 6808
rect 24523 6788 24561 6822
rect 24595 6788 24610 6822
rect 23610 6782 24384 6788
rect 23502 6725 23578 6772
rect 24362 6756 24384 6782
rect 24436 6756 24448 6788
rect 24500 6782 24610 6788
rect 24500 6756 24522 6782
rect 24682 6772 24712 6838
rect 24362 6742 24522 6756
rect 23502 6712 23538 6725
rect 19936 6641 19982 6679
rect 19936 6607 19942 6641
rect 19976 6607 19982 6641
rect 18486 6535 18492 6569
rect 18526 6535 18532 6569
rect 18486 6497 18532 6535
rect 18486 6463 18492 6497
rect 18526 6463 18532 6497
rect 18486 6425 18532 6463
rect 18486 6391 18492 6425
rect 18526 6391 18532 6425
rect 18486 6353 18532 6391
rect 18486 6319 18492 6353
rect 18526 6319 18532 6353
rect 18486 6281 18532 6319
rect 18862 6569 19042 6600
rect 18862 6535 18884 6569
rect 18918 6540 19042 6569
rect 18862 6497 18894 6535
rect 18862 6463 18884 6497
rect 18862 6425 18894 6463
rect 18862 6391 18884 6425
rect 18862 6360 18894 6391
rect 19010 6360 19042 6540
rect 18862 6353 19042 6360
rect 18862 6319 18884 6353
rect 18918 6319 19042 6353
rect 18862 6310 19042 6319
rect 19936 6569 19982 6607
rect 19936 6535 19942 6569
rect 19976 6535 19982 6569
rect 19936 6497 19982 6535
rect 19936 6463 19942 6497
rect 19976 6463 19982 6497
rect 19936 6425 19982 6463
rect 19936 6391 19942 6425
rect 19976 6391 19982 6425
rect 19936 6353 19982 6391
rect 19936 6319 19942 6353
rect 19976 6319 19982 6353
rect 18486 6247 18492 6281
rect 18526 6247 18532 6281
rect 18486 6209 18532 6247
rect 18486 6175 18492 6209
rect 18526 6175 18532 6209
rect 18486 6137 18532 6175
rect 18486 6103 18492 6137
rect 18526 6103 18532 6137
rect 18486 6065 18532 6103
rect 18486 6031 18492 6065
rect 18526 6031 18532 6065
rect 18486 5993 18532 6031
rect 18486 5959 18492 5993
rect 18526 5959 18532 5993
rect 18486 5921 18532 5959
rect 18486 5887 18492 5921
rect 18526 5887 18532 5921
rect 18486 5849 18532 5887
rect 18486 5815 18492 5849
rect 18526 5815 18532 5849
rect 18486 5777 18532 5815
rect 18486 5743 18492 5777
rect 18526 5743 18532 5777
rect 18486 5705 18532 5743
rect 18486 5671 18492 5705
rect 18526 5671 18532 5705
rect 18486 5633 18532 5671
rect 18486 5599 18492 5633
rect 18526 5599 18532 5633
rect 18486 5561 18532 5599
rect 18486 5527 18492 5561
rect 18526 5527 18532 5561
rect 18486 5489 18532 5527
rect 18486 5455 18492 5489
rect 18526 5455 18532 5489
rect 18486 5417 18532 5455
rect 18486 5383 18492 5417
rect 18526 5383 18532 5417
rect 18486 5345 18532 5383
rect 18486 5311 18492 5345
rect 18526 5311 18532 5345
rect 18486 5273 18532 5311
rect 18486 5239 18492 5273
rect 18526 5239 18532 5273
rect 18486 5201 18532 5239
rect 18486 5167 18492 5201
rect 18526 5167 18532 5201
rect 18486 5129 18532 5167
rect 18486 5095 18492 5129
rect 18526 5095 18532 5129
rect 18486 5057 18532 5095
rect 18486 5023 18492 5057
rect 18526 5023 18532 5057
rect 18486 4985 18532 5023
rect 18486 4951 18492 4985
rect 18526 4951 18532 4985
rect 18486 4913 18532 4951
rect 18486 4879 18492 4913
rect 18526 4879 18532 4913
rect 18486 4841 18532 4879
rect 18486 4807 18492 4841
rect 18526 4807 18532 4841
rect 18486 4769 18532 4807
rect 18486 4735 18492 4769
rect 18526 4735 18532 4769
rect 18486 4697 18532 4735
rect 18486 4663 18492 4697
rect 18526 4663 18532 4697
rect 18486 4625 18532 4663
rect 18486 4591 18492 4625
rect 18526 4591 18532 4625
rect 18486 4548 18532 4591
rect 18878 6281 18924 6310
rect 18878 6247 18884 6281
rect 18918 6247 18924 6281
rect 18878 6209 18924 6247
rect 18878 6175 18884 6209
rect 18918 6175 18924 6209
rect 18878 6137 18924 6175
rect 18878 6103 18884 6137
rect 18918 6103 18924 6137
rect 18878 6065 18924 6103
rect 18878 6031 18884 6065
rect 18918 6031 18924 6065
rect 18878 5993 18924 6031
rect 18878 5959 18884 5993
rect 18918 5959 18924 5993
rect 18878 5921 18924 5959
rect 18878 5887 18884 5921
rect 18918 5887 18924 5921
rect 18878 5849 18924 5887
rect 18878 5815 18884 5849
rect 18918 5815 18924 5849
rect 18878 5777 18924 5815
rect 18878 5743 18884 5777
rect 18918 5743 18924 5777
rect 18878 5705 18924 5743
rect 18878 5671 18884 5705
rect 18918 5671 18924 5705
rect 18878 5633 18924 5671
rect 18878 5599 18884 5633
rect 18918 5599 18924 5633
rect 18878 5561 18924 5599
rect 18878 5527 18884 5561
rect 18918 5527 18924 5561
rect 18878 5489 18924 5527
rect 18878 5455 18884 5489
rect 18918 5455 18924 5489
rect 18878 5417 18924 5455
rect 18878 5383 18884 5417
rect 18918 5383 18924 5417
rect 18878 5345 18924 5383
rect 18878 5311 18884 5345
rect 18918 5311 18924 5345
rect 18878 5273 18924 5311
rect 18878 5239 18884 5273
rect 18918 5239 18924 5273
rect 18878 5201 18924 5239
rect 18878 5167 18884 5201
rect 18918 5167 18924 5201
rect 18878 5129 18924 5167
rect 18878 5095 18884 5129
rect 18918 5095 18924 5129
rect 18878 5057 18924 5095
rect 18878 5023 18884 5057
rect 18918 5023 18924 5057
rect 18878 4985 18924 5023
rect 18878 4951 18884 4985
rect 18918 4951 18924 4985
rect 18878 4913 18924 4951
rect 18878 4879 18884 4913
rect 18918 4879 18924 4913
rect 18878 4841 18924 4879
rect 18878 4807 18884 4841
rect 18918 4807 18924 4841
rect 18878 4769 18924 4807
rect 18878 4735 18884 4769
rect 18918 4735 18924 4769
rect 18878 4697 18924 4735
rect 18878 4663 18884 4697
rect 18918 4663 18924 4697
rect 18878 4625 18924 4663
rect 18878 4591 18884 4625
rect 18918 4591 18924 4625
rect 18878 4548 18924 4591
rect 19936 6281 19982 6319
rect 19936 6247 19942 6281
rect 19976 6247 19982 6281
rect 19936 6209 19982 6247
rect 19936 6175 19942 6209
rect 19976 6175 19982 6209
rect 19936 6137 19982 6175
rect 19936 6103 19942 6137
rect 19976 6103 19982 6137
rect 19936 6065 19982 6103
rect 19936 6031 19942 6065
rect 19976 6031 19982 6065
rect 19936 5993 19982 6031
rect 19936 5959 19942 5993
rect 19976 5959 19982 5993
rect 19936 5921 19982 5959
rect 19936 5887 19942 5921
rect 19976 5887 19982 5921
rect 19936 5849 19982 5887
rect 19936 5815 19942 5849
rect 19976 5815 19982 5849
rect 23532 6691 23538 6712
rect 23572 6691 23578 6725
rect 23532 6653 23578 6691
rect 23532 6619 23538 6653
rect 23572 6619 23578 6653
rect 23532 6581 23578 6619
rect 23532 6547 23538 6581
rect 23572 6547 23578 6581
rect 23532 6509 23578 6547
rect 23532 6475 23538 6509
rect 23572 6475 23578 6509
rect 23532 6437 23578 6475
rect 23532 6403 23538 6437
rect 23572 6403 23578 6437
rect 23532 6365 23578 6403
rect 23532 6331 23538 6365
rect 23572 6331 23578 6365
rect 23532 6293 23578 6331
rect 23532 6259 23538 6293
rect 23572 6259 23578 6293
rect 23532 6221 23578 6259
rect 23532 6187 23538 6221
rect 23572 6187 23578 6221
rect 23532 6149 23578 6187
rect 23532 6115 23538 6149
rect 23572 6115 23578 6149
rect 23532 6077 23578 6115
rect 23532 6043 23538 6077
rect 23572 6043 23578 6077
rect 23532 6005 23578 6043
rect 23532 5971 23538 6005
rect 23572 5971 23578 6005
rect 23532 5933 23578 5971
rect 23532 5899 23538 5933
rect 23572 5899 23578 5933
rect 23532 5861 23578 5899
rect 23532 5842 23538 5861
rect 19936 5777 19982 5815
rect 19936 5743 19942 5777
rect 19976 5743 19982 5777
rect 19936 5705 19982 5743
rect 19936 5671 19942 5705
rect 19976 5671 19982 5705
rect 19936 5633 19982 5671
rect 23502 5827 23538 5842
rect 23572 5827 23578 5861
rect 23502 5780 23578 5827
rect 24642 6725 24712 6772
rect 24642 6691 24648 6725
rect 24682 6702 24712 6725
rect 25002 6885 25038 6892
rect 25072 6885 25078 6919
rect 25002 6838 25078 6885
rect 25002 6772 25032 6838
rect 25142 6828 25302 6942
rect 26142 6919 26188 6957
rect 26142 6885 26148 6919
rect 26182 6902 26188 6919
rect 37806 7449 37852 7487
rect 37806 7415 37812 7449
rect 37846 7415 37852 7449
rect 37806 7377 37852 7415
rect 37806 7343 37812 7377
rect 37846 7343 37852 7377
rect 37806 7305 37852 7343
rect 37806 7271 37812 7305
rect 37846 7271 37852 7305
rect 37806 7233 37852 7271
rect 37806 7199 37812 7233
rect 37846 7199 37852 7233
rect 37806 7161 37852 7199
rect 37806 7127 37812 7161
rect 37846 7127 37852 7161
rect 37806 7089 37852 7127
rect 37806 7055 37812 7089
rect 37846 7055 37852 7089
rect 37806 7017 37852 7055
rect 37806 6983 37812 7017
rect 37846 6983 37852 7017
rect 37806 6945 37852 6983
rect 37806 6911 37812 6945
rect 37846 6911 37852 6945
rect 26182 6885 26212 6902
rect 25852 6828 26012 6842
rect 26142 6838 26212 6885
rect 25110 6822 25874 6828
rect 25926 6822 25938 6828
rect 25990 6822 26110 6828
rect 25110 6788 25125 6822
rect 25159 6788 25197 6822
rect 25231 6788 25269 6822
rect 25303 6788 25341 6822
rect 25375 6788 25413 6822
rect 25447 6788 25485 6822
rect 25519 6788 25557 6822
rect 25591 6788 25629 6822
rect 25663 6788 25701 6822
rect 25735 6788 25773 6822
rect 25807 6788 25845 6822
rect 26023 6788 26061 6822
rect 26095 6788 26110 6822
rect 25110 6782 25874 6788
rect 25852 6776 25874 6782
rect 25926 6776 25938 6788
rect 25990 6782 26110 6788
rect 25990 6776 26012 6782
rect 25002 6725 25078 6772
rect 25852 6742 26012 6776
rect 26182 6772 26212 6838
rect 25002 6702 25038 6725
rect 24682 6691 24688 6702
rect 24642 6653 24688 6691
rect 24642 6619 24648 6653
rect 24682 6619 24688 6653
rect 24642 6581 24688 6619
rect 24642 6547 24648 6581
rect 24682 6547 24688 6581
rect 24642 6509 24688 6547
rect 24642 6475 24648 6509
rect 24682 6475 24688 6509
rect 24642 6437 24688 6475
rect 24642 6403 24648 6437
rect 24682 6403 24688 6437
rect 24642 6365 24688 6403
rect 24642 6331 24648 6365
rect 24682 6331 24688 6365
rect 24642 6293 24688 6331
rect 24642 6259 24648 6293
rect 24682 6259 24688 6293
rect 24642 6221 24688 6259
rect 24642 6187 24648 6221
rect 24682 6187 24688 6221
rect 24642 6149 24688 6187
rect 24642 6115 24648 6149
rect 24682 6115 24688 6149
rect 24642 6077 24688 6115
rect 24642 6043 24648 6077
rect 24682 6043 24688 6077
rect 24642 6005 24688 6043
rect 24642 5971 24648 6005
rect 24682 5971 24688 6005
rect 24642 5933 24688 5971
rect 24642 5899 24648 5933
rect 24682 5899 24688 5933
rect 24642 5861 24688 5899
rect 24642 5827 24648 5861
rect 24682 5842 24688 5861
rect 25032 6691 25038 6702
rect 25072 6691 25078 6725
rect 25032 6653 25078 6691
rect 25032 6619 25038 6653
rect 25072 6619 25078 6653
rect 25032 6581 25078 6619
rect 25032 6547 25038 6581
rect 25072 6547 25078 6581
rect 25032 6509 25078 6547
rect 25032 6475 25038 6509
rect 25072 6475 25078 6509
rect 25032 6437 25078 6475
rect 25032 6403 25038 6437
rect 25072 6403 25078 6437
rect 25032 6365 25078 6403
rect 25032 6331 25038 6365
rect 25072 6331 25078 6365
rect 25032 6293 25078 6331
rect 25032 6259 25038 6293
rect 25072 6259 25078 6293
rect 25032 6221 25078 6259
rect 25032 6187 25038 6221
rect 25072 6187 25078 6221
rect 25032 6149 25078 6187
rect 25032 6115 25038 6149
rect 25072 6115 25078 6149
rect 25032 6077 25078 6115
rect 25032 6043 25038 6077
rect 25072 6043 25078 6077
rect 25032 6005 25078 6043
rect 25032 5971 25038 6005
rect 25072 5971 25078 6005
rect 25032 5933 25078 5971
rect 25032 5899 25038 5933
rect 25072 5899 25078 5933
rect 25032 5861 25078 5899
rect 25032 5852 25038 5861
rect 24682 5827 24712 5842
rect 23502 5714 23532 5780
rect 23642 5770 23812 5802
rect 24642 5780 24712 5827
rect 23610 5764 24610 5770
rect 23610 5730 23625 5764
rect 23659 5763 23697 5764
rect 23731 5763 23769 5764
rect 23659 5730 23664 5763
rect 23803 5730 23841 5764
rect 23875 5730 23913 5764
rect 23947 5730 23985 5764
rect 24019 5730 24057 5764
rect 24091 5730 24129 5764
rect 24163 5730 24201 5764
rect 24235 5730 24273 5764
rect 24307 5730 24345 5764
rect 24379 5730 24417 5764
rect 24451 5730 24489 5764
rect 24523 5730 24561 5764
rect 24595 5730 24610 5764
rect 23610 5724 23664 5730
rect 23502 5667 23578 5714
rect 23642 5711 23664 5724
rect 23716 5711 23728 5730
rect 23780 5724 24610 5730
rect 23780 5711 23812 5724
rect 24682 5714 24712 5780
rect 23642 5682 23812 5711
rect 23502 5652 23538 5667
rect 19936 5599 19942 5633
rect 19976 5599 19982 5633
rect 19936 5561 19982 5599
rect 19936 5527 19942 5561
rect 19976 5527 19982 5561
rect 19936 5489 19982 5527
rect 19936 5455 19942 5489
rect 19976 5455 19982 5489
rect 19936 5417 19982 5455
rect 19936 5383 19942 5417
rect 19976 5383 19982 5417
rect 19936 5345 19982 5383
rect 19936 5311 19942 5345
rect 19976 5311 19982 5345
rect 19936 5273 19982 5311
rect 19936 5239 19942 5273
rect 19976 5239 19982 5273
rect 19936 5201 19982 5239
rect 19936 5167 19942 5201
rect 19976 5167 19982 5201
rect 19936 5129 19982 5167
rect 23532 5633 23538 5652
rect 23572 5633 23578 5667
rect 23532 5595 23578 5633
rect 23532 5561 23538 5595
rect 23572 5561 23578 5595
rect 23532 5523 23578 5561
rect 23532 5489 23538 5523
rect 23572 5489 23578 5523
rect 23532 5451 23578 5489
rect 23532 5417 23538 5451
rect 23572 5417 23578 5451
rect 23532 5379 23578 5417
rect 23532 5345 23538 5379
rect 23572 5345 23578 5379
rect 23532 5307 23578 5345
rect 23532 5273 23538 5307
rect 23572 5273 23578 5307
rect 23532 5235 23578 5273
rect 23532 5201 23538 5235
rect 23572 5201 23578 5235
rect 23532 5163 23578 5201
rect 19936 5095 19942 5129
rect 19976 5095 19982 5129
rect 19936 5057 19982 5095
rect 19936 5023 19942 5057
rect 19976 5023 19982 5057
rect 19936 4985 19982 5023
rect 19936 4951 19942 4985
rect 19976 4951 19982 4985
rect 19936 4913 19982 4951
rect 19936 4879 19942 4913
rect 19976 4879 19982 4913
rect 19936 4841 19982 4879
rect 19936 4807 19942 4841
rect 19976 4807 19982 4841
rect 19936 4769 19982 4807
rect 19936 4735 19942 4769
rect 19976 4735 19982 4769
rect 19936 4697 19982 4735
rect 20522 5133 20572 5147
rect 20522 5099 20530 5133
rect 20564 5099 20572 5133
rect 20522 5061 20572 5099
rect 20522 5027 20530 5061
rect 20564 5027 20572 5061
rect 20522 4989 20572 5027
rect 20522 4955 20530 4989
rect 20564 4955 20572 4989
rect 20522 4917 20572 4955
rect 20522 4883 20530 4917
rect 20564 4883 20572 4917
rect 20522 4845 20572 4883
rect 20522 4811 20530 4845
rect 20564 4811 20572 4845
rect 20522 4773 20572 4811
rect 20522 4739 20530 4773
rect 20564 4739 20572 4773
rect 20522 4726 20572 4739
rect 20840 5133 20890 5147
rect 20840 5099 20848 5133
rect 20882 5099 20890 5133
rect 20840 5061 20890 5099
rect 20840 5027 20848 5061
rect 20882 5027 20890 5061
rect 20840 4989 20890 5027
rect 20840 4955 20848 4989
rect 20882 4955 20890 4989
rect 20840 4917 20890 4955
rect 20840 4883 20848 4917
rect 20882 4883 20890 4917
rect 20840 4845 20890 4883
rect 20840 4811 20848 4845
rect 20882 4811 20890 4845
rect 20840 4773 20890 4811
rect 20840 4739 20848 4773
rect 20882 4739 20890 4773
rect 20840 4726 20890 4739
rect 21158 5133 21208 5147
rect 21158 5099 21166 5133
rect 21200 5099 21208 5133
rect 21158 5061 21208 5099
rect 21158 5027 21166 5061
rect 21200 5027 21208 5061
rect 21158 4989 21208 5027
rect 21158 4955 21166 4989
rect 21200 4955 21208 4989
rect 21158 4917 21208 4955
rect 21158 4883 21166 4917
rect 21200 4883 21208 4917
rect 21158 4845 21208 4883
rect 21158 4811 21166 4845
rect 21200 4811 21208 4845
rect 21158 4773 21208 4811
rect 21158 4739 21166 4773
rect 21200 4739 21208 4773
rect 21158 4726 21208 4739
rect 21476 5133 21526 5147
rect 21476 5099 21484 5133
rect 21518 5099 21526 5133
rect 21476 5061 21526 5099
rect 21476 5027 21484 5061
rect 21518 5027 21526 5061
rect 21476 4989 21526 5027
rect 21476 4955 21484 4989
rect 21518 4955 21526 4989
rect 21476 4917 21526 4955
rect 21476 4883 21484 4917
rect 21518 4883 21526 4917
rect 21476 4845 21526 4883
rect 21476 4811 21484 4845
rect 21518 4811 21526 4845
rect 21476 4773 21526 4811
rect 23532 5129 23538 5163
rect 23572 5129 23578 5163
rect 23532 5091 23578 5129
rect 23532 5057 23538 5091
rect 23572 5057 23578 5091
rect 23532 5019 23578 5057
rect 23532 4985 23538 5019
rect 23572 4985 23578 5019
rect 23532 4947 23578 4985
rect 23532 4913 23538 4947
rect 23572 4913 23578 4947
rect 23532 4875 23578 4913
rect 23532 4841 23538 4875
rect 23572 4841 23578 4875
rect 23532 4803 23578 4841
rect 23532 4782 23538 4803
rect 21476 4739 21484 4773
rect 21518 4739 21526 4773
rect 21476 4726 21526 4739
rect 23502 4769 23538 4782
rect 23572 4769 23578 4803
rect 19936 4663 19942 4697
rect 19976 4663 19982 4697
rect 19936 4625 19982 4663
rect 19936 4591 19942 4625
rect 19976 4591 19982 4625
rect 23502 4722 23578 4769
rect 24642 5667 24712 5714
rect 24642 5633 24648 5667
rect 24682 5652 24712 5667
rect 25002 5827 25038 5852
rect 25072 5827 25078 5861
rect 25002 5780 25078 5827
rect 26142 6725 26212 6772
rect 26142 6691 26148 6725
rect 26182 6712 26212 6725
rect 27710 6877 27760 6891
rect 27710 6843 27718 6877
rect 27752 6843 27760 6877
rect 27710 6805 27760 6843
rect 27710 6771 27718 6805
rect 27752 6771 27760 6805
rect 27710 6733 27760 6771
rect 26182 6691 26188 6712
rect 26142 6653 26188 6691
rect 26142 6619 26148 6653
rect 26182 6619 26188 6653
rect 26142 6581 26188 6619
rect 26142 6547 26148 6581
rect 26182 6547 26188 6581
rect 26142 6509 26188 6547
rect 26142 6475 26148 6509
rect 26182 6475 26188 6509
rect 26142 6437 26188 6475
rect 27710 6699 27718 6733
rect 27752 6699 27760 6733
rect 27710 6661 27760 6699
rect 27710 6627 27718 6661
rect 27752 6627 27760 6661
rect 27710 6589 27760 6627
rect 27710 6555 27718 6589
rect 27752 6555 27760 6589
rect 27710 6517 27760 6555
rect 27710 6483 27718 6517
rect 27752 6483 27760 6517
rect 27710 6470 27760 6483
rect 27964 6877 28146 6900
rect 27964 6865 28036 6877
rect 28070 6865 28146 6877
rect 27964 6813 28035 6865
rect 28087 6813 28146 6865
rect 27964 6805 28146 6813
rect 27964 6801 28036 6805
rect 28070 6801 28146 6805
rect 27964 6749 28035 6801
rect 28087 6749 28146 6801
rect 27964 6737 28146 6749
rect 27964 6685 28035 6737
rect 28087 6685 28146 6737
rect 27964 6673 28146 6685
rect 27964 6621 28035 6673
rect 28087 6621 28146 6673
rect 27964 6609 28146 6621
rect 27964 6557 28035 6609
rect 28087 6557 28146 6609
rect 27964 6555 28036 6557
rect 28070 6555 28146 6557
rect 27964 6545 28146 6555
rect 27964 6493 28035 6545
rect 28087 6493 28146 6545
rect 27964 6483 28036 6493
rect 28070 6483 28146 6493
rect 27964 6466 28146 6483
rect 28342 6877 28732 6900
rect 28342 6843 28354 6877
rect 28388 6843 28672 6877
rect 28706 6843 28732 6877
rect 28342 6805 28732 6843
rect 28342 6771 28354 6805
rect 28388 6771 28672 6805
rect 28706 6771 28732 6805
rect 28342 6733 28732 6771
rect 28342 6699 28354 6733
rect 28388 6699 28672 6733
rect 28706 6699 28732 6733
rect 28342 6661 28732 6699
rect 28342 6627 28354 6661
rect 28388 6627 28672 6661
rect 28706 6627 28732 6661
rect 28342 6589 28732 6627
rect 28342 6555 28354 6589
rect 28388 6555 28672 6589
rect 28706 6555 28732 6589
rect 28342 6517 28732 6555
rect 28342 6483 28354 6517
rect 28388 6483 28672 6517
rect 28706 6483 28732 6517
rect 28342 6470 28732 6483
rect 28974 6877 29364 6900
rect 28974 6843 28990 6877
rect 29024 6843 29308 6877
rect 29342 6843 29364 6877
rect 28974 6805 29364 6843
rect 28974 6771 28990 6805
rect 29024 6771 29308 6805
rect 29342 6771 29364 6805
rect 28974 6733 29364 6771
rect 28974 6699 28990 6733
rect 29024 6699 29308 6733
rect 29342 6699 29364 6733
rect 28974 6661 29364 6699
rect 28974 6627 28990 6661
rect 29024 6627 29308 6661
rect 29342 6627 29364 6661
rect 28974 6589 29364 6627
rect 28974 6555 28990 6589
rect 29024 6555 29308 6589
rect 29342 6555 29364 6589
rect 28974 6517 29364 6555
rect 28974 6483 28990 6517
rect 29024 6483 29308 6517
rect 29342 6483 29364 6517
rect 28974 6470 29364 6483
rect 29618 6877 29668 6891
rect 29618 6843 29626 6877
rect 29660 6843 29668 6877
rect 29618 6805 29668 6843
rect 29618 6771 29626 6805
rect 29660 6771 29668 6805
rect 29618 6733 29668 6771
rect 29618 6699 29626 6733
rect 29660 6699 29668 6733
rect 29618 6661 29668 6699
rect 29618 6627 29626 6661
rect 29660 6627 29668 6661
rect 37806 6873 37852 6911
rect 37806 6839 37812 6873
rect 37846 6839 37852 6873
rect 37806 6801 37852 6839
rect 37806 6767 37812 6801
rect 37846 6767 37852 6801
rect 37806 6729 37852 6767
rect 37806 6695 37812 6729
rect 37846 6695 37852 6729
rect 37806 6657 37852 6695
rect 29618 6589 29668 6627
rect 29618 6555 29626 6589
rect 29660 6555 29668 6589
rect 29618 6517 29668 6555
rect 29618 6483 29626 6517
rect 29660 6483 29668 6517
rect 29618 6470 29668 6483
rect 37595 6636 37683 6651
rect 37595 6584 37612 6636
rect 37664 6584 37683 6636
rect 37595 6572 37683 6584
rect 37595 6520 37612 6572
rect 37664 6520 37683 6572
rect 37595 6508 37683 6520
rect 37595 6456 37612 6508
rect 37664 6456 37683 6508
rect 37595 6443 37683 6456
rect 37806 6623 37812 6657
rect 37846 6623 37852 6657
rect 38064 8241 38110 8288
rect 38064 8207 38070 8241
rect 38104 8207 38110 8241
rect 38064 8169 38110 8207
rect 38064 8135 38070 8169
rect 38104 8135 38110 8169
rect 38064 8097 38110 8135
rect 38064 8063 38070 8097
rect 38104 8063 38110 8097
rect 38064 8025 38110 8063
rect 38064 7991 38070 8025
rect 38104 7991 38110 8025
rect 38064 7953 38110 7991
rect 38064 7919 38070 7953
rect 38104 7919 38110 7953
rect 38064 7881 38110 7919
rect 38064 7847 38070 7881
rect 38104 7847 38110 7881
rect 38064 7809 38110 7847
rect 38064 7775 38070 7809
rect 38104 7775 38110 7809
rect 38064 7737 38110 7775
rect 38064 7703 38070 7737
rect 38104 7703 38110 7737
rect 38064 7665 38110 7703
rect 38064 7631 38070 7665
rect 38104 7631 38110 7665
rect 38064 7593 38110 7631
rect 38064 7559 38070 7593
rect 38104 7559 38110 7593
rect 38322 8241 38368 8288
rect 38322 8207 38328 8241
rect 38362 8207 38368 8241
rect 38322 8169 38368 8207
rect 38322 8135 38328 8169
rect 38362 8135 38368 8169
rect 38322 8097 38368 8135
rect 38322 8063 38328 8097
rect 38362 8063 38368 8097
rect 38322 8025 38368 8063
rect 38322 7991 38328 8025
rect 38362 7991 38368 8025
rect 38322 7953 38368 7991
rect 38322 7919 38328 7953
rect 38362 7919 38368 7953
rect 38322 7881 38368 7919
rect 38322 7847 38328 7881
rect 38362 7847 38368 7881
rect 38322 7809 38368 7847
rect 38322 7775 38328 7809
rect 38362 7775 38368 7809
rect 38322 7737 38368 7775
rect 38322 7703 38328 7737
rect 38362 7703 38368 7737
rect 38322 7665 38368 7703
rect 38322 7631 38328 7665
rect 38362 7631 38368 7665
rect 38322 7593 38368 7631
rect 38322 7561 38328 7593
rect 38064 7521 38110 7559
rect 38064 7487 38070 7521
rect 38104 7487 38110 7521
rect 38064 7449 38110 7487
rect 38064 7415 38070 7449
rect 38104 7415 38110 7449
rect 38064 7377 38110 7415
rect 38064 7343 38070 7377
rect 38104 7343 38110 7377
rect 38302 7559 38328 7561
rect 38362 7561 38368 7593
rect 38580 8241 38626 8288
rect 38580 8207 38586 8241
rect 38620 8207 38626 8241
rect 38580 8169 38626 8207
rect 38580 8135 38586 8169
rect 38620 8135 38626 8169
rect 38580 8097 38626 8135
rect 38580 8063 38586 8097
rect 38620 8063 38626 8097
rect 38580 8025 38626 8063
rect 38580 7991 38586 8025
rect 38620 7991 38626 8025
rect 38580 7953 38626 7991
rect 38580 7919 38586 7953
rect 38620 7919 38626 7953
rect 38580 7881 38626 7919
rect 38580 7847 38586 7881
rect 38620 7847 38626 7881
rect 38580 7809 38626 7847
rect 38580 7775 38586 7809
rect 38620 7775 38626 7809
rect 38580 7737 38626 7775
rect 38580 7703 38586 7737
rect 38620 7703 38626 7737
rect 38580 7665 38626 7703
rect 38580 7631 38586 7665
rect 38620 7631 38626 7665
rect 38580 7593 38626 7631
rect 38362 7559 38388 7561
rect 38302 7521 38388 7559
rect 38302 7515 38328 7521
rect 38362 7515 38388 7521
rect 38302 7463 38319 7515
rect 38371 7463 38388 7515
rect 38302 7451 38388 7463
rect 38302 7399 38319 7451
rect 38371 7399 38388 7451
rect 38302 7377 38388 7399
rect 38302 7356 38328 7377
rect 38064 7305 38110 7343
rect 38064 7271 38070 7305
rect 38104 7271 38110 7305
rect 38064 7233 38110 7271
rect 38064 7199 38070 7233
rect 38104 7199 38110 7233
rect 38064 7161 38110 7199
rect 38064 7127 38070 7161
rect 38104 7127 38110 7161
rect 38064 7089 38110 7127
rect 38064 7055 38070 7089
rect 38104 7055 38110 7089
rect 38064 7017 38110 7055
rect 38064 6983 38070 7017
rect 38104 6983 38110 7017
rect 38064 6945 38110 6983
rect 38064 6911 38070 6945
rect 38104 6911 38110 6945
rect 38064 6873 38110 6911
rect 38064 6839 38070 6873
rect 38104 6839 38110 6873
rect 38064 6801 38110 6839
rect 38064 6767 38070 6801
rect 38104 6767 38110 6801
rect 38064 6729 38110 6767
rect 38064 6695 38070 6729
rect 38104 6695 38110 6729
rect 38064 6657 38110 6695
rect 38064 6651 38070 6657
rect 37806 6585 37852 6623
rect 37806 6551 37812 6585
rect 37846 6551 37852 6585
rect 37806 6513 37852 6551
rect 37806 6479 37812 6513
rect 37846 6479 37852 6513
rect 26142 6403 26148 6437
rect 26182 6403 26188 6437
rect 26142 6365 26188 6403
rect 26142 6331 26148 6365
rect 26182 6331 26188 6365
rect 26142 6293 26188 6331
rect 26142 6259 26148 6293
rect 26182 6259 26188 6293
rect 26142 6221 26188 6259
rect 26142 6187 26148 6221
rect 26182 6187 26188 6221
rect 26142 6149 26188 6187
rect 26142 6115 26148 6149
rect 26182 6115 26188 6149
rect 37806 6441 37852 6479
rect 38056 6638 38070 6651
rect 38104 6651 38110 6657
rect 38322 7343 38328 7356
rect 38362 7356 38388 7377
rect 38580 7559 38586 7593
rect 38620 7559 38626 7593
rect 38580 7521 38626 7559
rect 38580 7487 38586 7521
rect 38620 7487 38626 7521
rect 38580 7449 38626 7487
rect 38580 7415 38586 7449
rect 38620 7415 38626 7449
rect 38580 7377 38626 7415
rect 38362 7343 38368 7356
rect 38322 7305 38368 7343
rect 38322 7271 38328 7305
rect 38362 7271 38368 7305
rect 38322 7233 38368 7271
rect 38322 7199 38328 7233
rect 38362 7199 38368 7233
rect 38322 7161 38368 7199
rect 38322 7127 38328 7161
rect 38362 7127 38368 7161
rect 38322 7089 38368 7127
rect 38322 7055 38328 7089
rect 38362 7055 38368 7089
rect 38322 7017 38368 7055
rect 38322 6983 38328 7017
rect 38362 6983 38368 7017
rect 38322 6945 38368 6983
rect 38322 6911 38328 6945
rect 38362 6911 38368 6945
rect 38322 6873 38368 6911
rect 38322 6839 38328 6873
rect 38362 6839 38368 6873
rect 38322 6801 38368 6839
rect 38322 6767 38328 6801
rect 38362 6767 38368 6801
rect 38322 6729 38368 6767
rect 38322 6695 38328 6729
rect 38362 6695 38368 6729
rect 38322 6657 38368 6695
rect 38104 6638 38118 6651
rect 38056 6586 38060 6638
rect 38112 6586 38118 6638
rect 38056 6585 38118 6586
rect 38056 6574 38070 6585
rect 38104 6574 38118 6585
rect 38056 6522 38060 6574
rect 38112 6522 38118 6574
rect 38056 6513 38118 6522
rect 38056 6510 38070 6513
rect 38104 6510 38118 6513
rect 38056 6458 38060 6510
rect 38112 6458 38118 6510
rect 38056 6443 38118 6458
rect 38322 6623 38328 6657
rect 38362 6623 38368 6657
rect 38580 7343 38586 7377
rect 38620 7343 38626 7377
rect 38580 7305 38626 7343
rect 38580 7271 38586 7305
rect 38620 7271 38626 7305
rect 38580 7233 38626 7271
rect 38580 7199 38586 7233
rect 38620 7199 38626 7233
rect 38580 7161 38626 7199
rect 38580 7127 38586 7161
rect 38620 7127 38626 7161
rect 38580 7089 38626 7127
rect 38838 8241 38884 8288
rect 38838 8207 38844 8241
rect 38878 8207 38884 8241
rect 38838 8169 38884 8207
rect 38838 8135 38844 8169
rect 38878 8135 38884 8169
rect 38838 8097 38884 8135
rect 38838 8063 38844 8097
rect 38878 8063 38884 8097
rect 38838 8025 38884 8063
rect 38838 7991 38844 8025
rect 38878 7991 38884 8025
rect 38838 7953 38884 7991
rect 38838 7919 38844 7953
rect 38878 7919 38884 7953
rect 38838 7881 38884 7919
rect 38838 7847 38844 7881
rect 38878 7847 38884 7881
rect 38838 7809 38884 7847
rect 38838 7775 38844 7809
rect 38878 7775 38884 7809
rect 38838 7737 38884 7775
rect 38838 7703 38844 7737
rect 38878 7703 38884 7737
rect 38838 7665 38884 7703
rect 38838 7631 38844 7665
rect 38878 7631 38884 7665
rect 38838 7593 38884 7631
rect 38838 7559 38844 7593
rect 38878 7559 38884 7593
rect 38838 7521 38884 7559
rect 38838 7487 38844 7521
rect 38878 7487 38884 7521
rect 38838 7449 38884 7487
rect 38838 7415 38844 7449
rect 38878 7415 38884 7449
rect 38838 7377 38884 7415
rect 38838 7343 38844 7377
rect 38878 7343 38884 7377
rect 38838 7305 38884 7343
rect 38838 7271 38844 7305
rect 38878 7271 38884 7305
rect 38838 7233 38884 7271
rect 38838 7199 38844 7233
rect 38878 7199 38884 7233
rect 38838 7161 38884 7199
rect 38838 7127 38844 7161
rect 38878 7127 38884 7161
rect 38838 7125 38884 7127
rect 39096 8241 39142 8288
rect 39096 8207 39102 8241
rect 39136 8207 39142 8241
rect 39096 8169 39142 8207
rect 39096 8135 39102 8169
rect 39136 8135 39142 8169
rect 39096 8097 39142 8135
rect 39096 8063 39102 8097
rect 39136 8063 39142 8097
rect 39096 8025 39142 8063
rect 39096 7991 39102 8025
rect 39136 7991 39142 8025
rect 39096 7953 39142 7991
rect 39096 7919 39102 7953
rect 39136 7919 39142 7953
rect 39096 7881 39142 7919
rect 39096 7847 39102 7881
rect 39136 7847 39142 7881
rect 39096 7809 39142 7847
rect 39096 7775 39102 7809
rect 39136 7775 39142 7809
rect 39096 7737 39142 7775
rect 39096 7703 39102 7737
rect 39136 7703 39142 7737
rect 39096 7665 39142 7703
rect 39096 7631 39102 7665
rect 39136 7631 39142 7665
rect 39096 7593 39142 7631
rect 39096 7559 39102 7593
rect 39136 7559 39142 7593
rect 39096 7521 39142 7559
rect 39096 7487 39102 7521
rect 39136 7487 39142 7521
rect 39096 7449 39142 7487
rect 39096 7415 39102 7449
rect 39136 7415 39142 7449
rect 39096 7377 39142 7415
rect 39096 7343 39102 7377
rect 39136 7343 39142 7377
rect 39096 7305 39142 7343
rect 39096 7271 39102 7305
rect 39136 7271 39142 7305
rect 39096 7233 39142 7271
rect 39096 7199 39102 7233
rect 39136 7199 39142 7233
rect 39096 7161 39142 7199
rect 39096 7127 39102 7161
rect 39136 7127 39142 7161
rect 38580 7055 38586 7089
rect 38620 7055 38626 7089
rect 38580 7017 38626 7055
rect 38580 6983 38586 7017
rect 38620 6983 38626 7017
rect 38580 6945 38626 6983
rect 38580 6911 38586 6945
rect 38620 6911 38626 6945
rect 38802 7112 38915 7125
rect 38802 7060 38835 7112
rect 38887 7060 38915 7112
rect 38802 7055 38844 7060
rect 38878 7055 38915 7060
rect 38802 7048 38915 7055
rect 38802 6996 38835 7048
rect 38887 6996 38915 7048
rect 38802 6984 38844 6996
rect 38878 6984 38915 6996
rect 38802 6932 38835 6984
rect 38887 6932 38915 6984
rect 38802 6918 38844 6932
rect 38580 6873 38626 6911
rect 38580 6839 38586 6873
rect 38620 6839 38626 6873
rect 38580 6801 38626 6839
rect 38580 6767 38586 6801
rect 38620 6767 38626 6801
rect 38580 6729 38626 6767
rect 38580 6695 38586 6729
rect 38620 6695 38626 6729
rect 38580 6657 38626 6695
rect 38580 6652 38586 6657
rect 38322 6585 38368 6623
rect 38322 6551 38328 6585
rect 38362 6551 38368 6585
rect 38322 6513 38368 6551
rect 38322 6479 38328 6513
rect 38362 6479 38368 6513
rect 37806 6407 37812 6441
rect 37846 6407 37852 6441
rect 37806 6369 37852 6407
rect 37806 6335 37812 6369
rect 37846 6335 37852 6369
rect 37806 6256 37852 6335
rect 38064 6441 38110 6443
rect 38064 6407 38070 6441
rect 38104 6407 38110 6441
rect 38064 6369 38110 6407
rect 38064 6335 38070 6369
rect 38104 6335 38110 6369
rect 38064 6288 38110 6335
rect 38322 6441 38368 6479
rect 38567 6637 38586 6652
rect 38620 6652 38626 6657
rect 38838 6911 38844 6918
rect 38878 6918 38915 6932
rect 39096 7089 39142 7127
rect 39354 8241 39400 8288
rect 39354 8207 39360 8241
rect 39394 8207 39400 8241
rect 39354 8169 39400 8207
rect 39354 8135 39360 8169
rect 39394 8135 39400 8169
rect 39354 8097 39400 8135
rect 39354 8063 39360 8097
rect 39394 8063 39400 8097
rect 39354 8025 39400 8063
rect 39354 7991 39360 8025
rect 39394 7991 39400 8025
rect 39354 7953 39400 7991
rect 39354 7919 39360 7953
rect 39394 7919 39400 7953
rect 39354 7881 39400 7919
rect 39354 7847 39360 7881
rect 39394 7847 39400 7881
rect 39354 7809 39400 7847
rect 39354 7775 39360 7809
rect 39394 7775 39400 7809
rect 39354 7737 39400 7775
rect 39354 7703 39360 7737
rect 39394 7703 39400 7737
rect 39354 7665 39400 7703
rect 39354 7631 39360 7665
rect 39394 7631 39400 7665
rect 39354 7593 39400 7631
rect 39354 7559 39360 7593
rect 39394 7559 39400 7593
rect 39354 7521 39400 7559
rect 39354 7487 39360 7521
rect 39394 7487 39400 7521
rect 39354 7449 39400 7487
rect 39354 7415 39360 7449
rect 39394 7415 39400 7449
rect 39354 7377 39400 7415
rect 39354 7343 39360 7377
rect 39394 7343 39400 7377
rect 39354 7305 39400 7343
rect 39354 7271 39360 7305
rect 39394 7271 39400 7305
rect 39354 7233 39400 7271
rect 39354 7199 39360 7233
rect 39394 7199 39400 7233
rect 39354 7161 39400 7199
rect 39354 7127 39360 7161
rect 39394 7127 39400 7161
rect 39354 7125 39400 7127
rect 39612 8241 39658 8288
rect 39612 8207 39618 8241
rect 39652 8207 39658 8241
rect 39612 8169 39658 8207
rect 39612 8135 39618 8169
rect 39652 8135 39658 8169
rect 39612 8097 39658 8135
rect 39612 8063 39618 8097
rect 39652 8063 39658 8097
rect 39612 8025 39658 8063
rect 39612 7991 39618 8025
rect 39652 7991 39658 8025
rect 39612 7953 39658 7991
rect 39612 7919 39618 7953
rect 39652 7919 39658 7953
rect 39612 7881 39658 7919
rect 39612 7847 39618 7881
rect 39652 7847 39658 7881
rect 39612 7809 39658 7847
rect 39612 7775 39618 7809
rect 39652 7775 39658 7809
rect 39612 7737 39658 7775
rect 39612 7703 39618 7737
rect 39652 7703 39658 7737
rect 39612 7665 39658 7703
rect 39612 7631 39618 7665
rect 39652 7631 39658 7665
rect 39612 7593 39658 7631
rect 39612 7559 39618 7593
rect 39652 7559 39658 7593
rect 39612 7521 39658 7559
rect 39612 7487 39618 7521
rect 39652 7487 39658 7521
rect 39612 7449 39658 7487
rect 39612 7415 39618 7449
rect 39652 7415 39658 7449
rect 39612 7377 39658 7415
rect 39612 7343 39618 7377
rect 39652 7343 39658 7377
rect 39612 7305 39658 7343
rect 39612 7271 39618 7305
rect 39652 7271 39658 7305
rect 39612 7233 39658 7271
rect 39612 7199 39618 7233
rect 39652 7199 39658 7233
rect 39612 7161 39658 7199
rect 39612 7127 39618 7161
rect 39652 7127 39658 7161
rect 39096 7055 39102 7089
rect 39136 7055 39142 7089
rect 39096 7017 39142 7055
rect 39096 6983 39102 7017
rect 39136 6983 39142 7017
rect 39096 6945 39142 6983
rect 38878 6911 38884 6918
rect 38838 6873 38884 6911
rect 38838 6839 38844 6873
rect 38878 6839 38884 6873
rect 38838 6801 38884 6839
rect 38838 6767 38844 6801
rect 38878 6767 38884 6801
rect 38838 6729 38884 6767
rect 38838 6695 38844 6729
rect 38878 6695 38884 6729
rect 38838 6657 38884 6695
rect 38620 6637 38638 6652
rect 38567 6585 38577 6637
rect 38629 6585 38638 6637
rect 38567 6573 38586 6585
rect 38620 6573 38638 6585
rect 38567 6521 38577 6573
rect 38629 6521 38638 6573
rect 38567 6513 38638 6521
rect 38567 6509 38586 6513
rect 38620 6509 38638 6513
rect 38567 6457 38577 6509
rect 38629 6457 38638 6509
rect 38567 6444 38638 6457
rect 38838 6623 38844 6657
rect 38878 6623 38884 6657
rect 39096 6911 39102 6945
rect 39136 6911 39142 6945
rect 39332 7110 39421 7125
rect 39332 7058 39351 7110
rect 39403 7058 39421 7110
rect 39332 7055 39360 7058
rect 39394 7055 39421 7058
rect 39332 7046 39421 7055
rect 39332 6994 39351 7046
rect 39403 6994 39421 7046
rect 39332 6983 39360 6994
rect 39394 6983 39421 6994
rect 39332 6982 39421 6983
rect 39332 6930 39351 6982
rect 39403 6930 39421 6982
rect 39332 6918 39360 6930
rect 39096 6873 39142 6911
rect 39096 6839 39102 6873
rect 39136 6839 39142 6873
rect 39096 6801 39142 6839
rect 39096 6767 39102 6801
rect 39136 6767 39142 6801
rect 39096 6729 39142 6767
rect 39096 6695 39102 6729
rect 39136 6695 39142 6729
rect 39096 6657 39142 6695
rect 39096 6651 39102 6657
rect 38838 6585 38884 6623
rect 38838 6551 38844 6585
rect 38878 6551 38884 6585
rect 38838 6513 38884 6551
rect 38838 6479 38844 6513
rect 38878 6479 38884 6513
rect 38322 6407 38328 6441
rect 38362 6407 38368 6441
rect 38322 6369 38368 6407
rect 38322 6335 38328 6369
rect 38362 6335 38368 6369
rect 38322 6288 38368 6335
rect 38580 6441 38626 6444
rect 38580 6407 38586 6441
rect 38620 6407 38626 6441
rect 38580 6369 38626 6407
rect 38580 6335 38586 6369
rect 38620 6335 38626 6369
rect 38580 6288 38626 6335
rect 38838 6441 38884 6479
rect 39081 6636 39102 6651
rect 39136 6651 39142 6657
rect 39354 6911 39360 6918
rect 39394 6918 39421 6930
rect 39612 7089 39658 7127
rect 39870 8241 39916 8288
rect 39870 8207 39876 8241
rect 39910 8207 39916 8241
rect 39870 8169 39916 8207
rect 39870 8135 39876 8169
rect 39910 8135 39916 8169
rect 39870 8097 39916 8135
rect 39870 8063 39876 8097
rect 39910 8063 39916 8097
rect 39870 8025 39916 8063
rect 39870 7991 39876 8025
rect 39910 7991 39916 8025
rect 39870 7953 39916 7991
rect 39870 7919 39876 7953
rect 39910 7919 39916 7953
rect 39870 7881 39916 7919
rect 39870 7847 39876 7881
rect 39910 7847 39916 7881
rect 39870 7809 39916 7847
rect 39870 7775 39876 7809
rect 39910 7775 39916 7809
rect 39870 7737 39916 7775
rect 39870 7703 39876 7737
rect 39910 7703 39916 7737
rect 39870 7665 39916 7703
rect 39870 7631 39876 7665
rect 39910 7631 39916 7665
rect 39870 7593 39916 7631
rect 39870 7559 39876 7593
rect 39910 7559 39916 7593
rect 39870 7521 39916 7559
rect 39870 7487 39876 7521
rect 39910 7487 39916 7521
rect 39870 7449 39916 7487
rect 39870 7415 39876 7449
rect 39910 7415 39916 7449
rect 39870 7377 39916 7415
rect 39870 7343 39876 7377
rect 39910 7343 39916 7377
rect 39870 7305 39916 7343
rect 39870 7271 39876 7305
rect 39910 7271 39916 7305
rect 39870 7233 39916 7271
rect 39870 7199 39876 7233
rect 39910 7199 39916 7233
rect 39870 7161 39916 7199
rect 39870 7127 39876 7161
rect 39910 7127 39916 7161
rect 39870 7125 39916 7127
rect 40128 8241 40174 8288
rect 40128 8207 40134 8241
rect 40168 8207 40174 8241
rect 40128 8169 40174 8207
rect 40128 8135 40134 8169
rect 40168 8135 40174 8169
rect 40128 8097 40174 8135
rect 40128 8063 40134 8097
rect 40168 8063 40174 8097
rect 40128 8025 40174 8063
rect 40128 7991 40134 8025
rect 40168 7991 40174 8025
rect 40128 7953 40174 7991
rect 40128 7919 40134 7953
rect 40168 7919 40174 7953
rect 40128 7881 40174 7919
rect 40128 7847 40134 7881
rect 40168 7847 40174 7881
rect 40128 7809 40174 7847
rect 40128 7775 40134 7809
rect 40168 7775 40174 7809
rect 40128 7737 40174 7775
rect 40128 7703 40134 7737
rect 40168 7703 40174 7737
rect 40128 7665 40174 7703
rect 40128 7631 40134 7665
rect 40168 7631 40174 7665
rect 40128 7593 40174 7631
rect 40128 7559 40134 7593
rect 40168 7559 40174 7593
rect 40128 7521 40174 7559
rect 40128 7487 40134 7521
rect 40168 7487 40174 7521
rect 40128 7449 40174 7487
rect 40128 7415 40134 7449
rect 40168 7415 40174 7449
rect 40128 7377 40174 7415
rect 40128 7343 40134 7377
rect 40168 7343 40174 7377
rect 40128 7305 40174 7343
rect 40128 7271 40134 7305
rect 40168 7271 40174 7305
rect 40128 7233 40174 7271
rect 40128 7199 40134 7233
rect 40168 7199 40174 7233
rect 40128 7161 40174 7199
rect 40128 7127 40134 7161
rect 40168 7127 40174 7161
rect 39612 7055 39618 7089
rect 39652 7055 39658 7089
rect 39612 7017 39658 7055
rect 39612 6983 39618 7017
rect 39652 6983 39658 7017
rect 39612 6945 39658 6983
rect 39394 6911 39400 6918
rect 39354 6873 39400 6911
rect 39354 6839 39360 6873
rect 39394 6839 39400 6873
rect 39354 6801 39400 6839
rect 39354 6767 39360 6801
rect 39394 6767 39400 6801
rect 39354 6729 39400 6767
rect 39354 6695 39360 6729
rect 39394 6695 39400 6729
rect 39354 6657 39400 6695
rect 39136 6636 39157 6651
rect 39081 6584 39093 6636
rect 39145 6584 39157 6636
rect 39081 6572 39102 6584
rect 39136 6572 39157 6584
rect 39081 6520 39093 6572
rect 39145 6520 39157 6572
rect 39081 6513 39157 6520
rect 39081 6508 39102 6513
rect 39136 6508 39157 6513
rect 39081 6456 39093 6508
rect 39145 6456 39157 6508
rect 39081 6444 39157 6456
rect 39354 6623 39360 6657
rect 39394 6623 39400 6657
rect 39612 6911 39618 6945
rect 39652 6911 39658 6945
rect 39846 7089 39936 7125
rect 39846 7078 39876 7089
rect 39910 7078 39936 7089
rect 39846 7026 39866 7078
rect 39918 7026 39936 7078
rect 39846 7017 39936 7026
rect 39846 7014 39876 7017
rect 39910 7014 39936 7017
rect 39846 6962 39866 7014
rect 39918 6962 39936 7014
rect 39846 6945 39936 6962
rect 39846 6918 39876 6945
rect 39612 6873 39658 6911
rect 39612 6839 39618 6873
rect 39652 6839 39658 6873
rect 39612 6801 39658 6839
rect 39612 6767 39618 6801
rect 39652 6767 39658 6801
rect 39612 6729 39658 6767
rect 39612 6695 39618 6729
rect 39652 6695 39658 6729
rect 39612 6657 39658 6695
rect 39612 6651 39618 6657
rect 39354 6585 39400 6623
rect 39354 6551 39360 6585
rect 39394 6551 39400 6585
rect 39354 6513 39400 6551
rect 39354 6479 39360 6513
rect 39394 6479 39400 6513
rect 38838 6407 38844 6441
rect 38878 6407 38884 6441
rect 38838 6369 38884 6407
rect 38838 6335 38844 6369
rect 38878 6335 38884 6369
rect 38838 6288 38884 6335
rect 39096 6441 39142 6444
rect 39096 6407 39102 6441
rect 39136 6407 39142 6441
rect 39096 6369 39142 6407
rect 39096 6335 39102 6369
rect 39136 6335 39142 6369
rect 39096 6288 39142 6335
rect 39354 6441 39400 6479
rect 39595 6637 39618 6651
rect 39652 6651 39658 6657
rect 39870 6911 39876 6918
rect 39910 6918 39936 6945
rect 40128 7089 40174 7127
rect 40386 8241 40432 8288
rect 40386 8207 40392 8241
rect 40426 8207 40432 8241
rect 40386 8169 40432 8207
rect 40386 8135 40392 8169
rect 40426 8135 40432 8169
rect 40386 8097 40432 8135
rect 40386 8063 40392 8097
rect 40426 8063 40432 8097
rect 40386 8025 40432 8063
rect 40386 7991 40392 8025
rect 40426 7991 40432 8025
rect 40386 7953 40432 7991
rect 40386 7919 40392 7953
rect 40426 7919 40432 7953
rect 40386 7881 40432 7919
rect 40386 7847 40392 7881
rect 40426 7847 40432 7881
rect 40386 7809 40432 7847
rect 40386 7775 40392 7809
rect 40426 7775 40432 7809
rect 40386 7737 40432 7775
rect 40386 7703 40392 7737
rect 40426 7703 40432 7737
rect 40386 7665 40432 7703
rect 40386 7631 40392 7665
rect 40426 7631 40432 7665
rect 40386 7593 40432 7631
rect 40386 7559 40392 7593
rect 40426 7559 40432 7593
rect 40386 7521 40432 7559
rect 40386 7487 40392 7521
rect 40426 7487 40432 7521
rect 40386 7449 40432 7487
rect 40386 7415 40392 7449
rect 40426 7415 40432 7449
rect 40386 7377 40432 7415
rect 40386 7343 40392 7377
rect 40426 7343 40432 7377
rect 40386 7305 40432 7343
rect 40386 7271 40392 7305
rect 40426 7271 40432 7305
rect 40386 7233 40432 7271
rect 40386 7199 40392 7233
rect 40426 7199 40432 7233
rect 40386 7161 40432 7199
rect 40386 7127 40392 7161
rect 40426 7127 40432 7161
rect 40386 7125 40432 7127
rect 40644 8241 40690 8288
rect 40644 8207 40650 8241
rect 40684 8207 40690 8241
rect 40644 8169 40690 8207
rect 40644 8135 40650 8169
rect 40684 8135 40690 8169
rect 40644 8097 40690 8135
rect 40644 8063 40650 8097
rect 40684 8063 40690 8097
rect 40644 8025 40690 8063
rect 40644 7991 40650 8025
rect 40684 7991 40690 8025
rect 40644 7953 40690 7991
rect 40644 7919 40650 7953
rect 40684 7919 40690 7953
rect 40644 7881 40690 7919
rect 40644 7847 40650 7881
rect 40684 7847 40690 7881
rect 40644 7809 40690 7847
rect 40644 7775 40650 7809
rect 40684 7775 40690 7809
rect 40644 7737 40690 7775
rect 40644 7703 40650 7737
rect 40684 7703 40690 7737
rect 40644 7665 40690 7703
rect 40644 7631 40650 7665
rect 40684 7631 40690 7665
rect 40644 7593 40690 7631
rect 40644 7559 40650 7593
rect 40684 7559 40690 7593
rect 40644 7521 40690 7559
rect 40644 7487 40650 7521
rect 40684 7487 40690 7521
rect 40644 7449 40690 7487
rect 40644 7415 40650 7449
rect 40684 7415 40690 7449
rect 40644 7377 40690 7415
rect 40644 7343 40650 7377
rect 40684 7343 40690 7377
rect 40644 7305 40690 7343
rect 40644 7271 40650 7305
rect 40684 7271 40690 7305
rect 40644 7233 40690 7271
rect 40644 7199 40650 7233
rect 40684 7199 40690 7233
rect 40644 7161 40690 7199
rect 40644 7127 40650 7161
rect 40684 7127 40690 7161
rect 40128 7055 40134 7089
rect 40168 7055 40174 7089
rect 40128 7017 40174 7055
rect 40128 6983 40134 7017
rect 40168 6983 40174 7017
rect 40128 6945 40174 6983
rect 39910 6911 39916 6918
rect 39870 6873 39916 6911
rect 39870 6839 39876 6873
rect 39910 6839 39916 6873
rect 39870 6801 39916 6839
rect 39870 6767 39876 6801
rect 39910 6767 39916 6801
rect 39870 6729 39916 6767
rect 39870 6695 39876 6729
rect 39910 6695 39916 6729
rect 39870 6657 39916 6695
rect 39652 6637 39672 6651
rect 39595 6585 39607 6637
rect 39659 6585 39672 6637
rect 39595 6573 39618 6585
rect 39652 6573 39672 6585
rect 39595 6521 39607 6573
rect 39659 6521 39672 6573
rect 39595 6513 39672 6521
rect 39595 6509 39618 6513
rect 39652 6509 39672 6513
rect 39595 6457 39607 6509
rect 39659 6457 39672 6509
rect 39595 6443 39672 6457
rect 39870 6623 39876 6657
rect 39910 6623 39916 6657
rect 40128 6911 40134 6945
rect 40168 6911 40174 6945
rect 40365 7111 40455 7125
rect 40365 7059 40383 7111
rect 40435 7059 40455 7111
rect 40365 7055 40392 7059
rect 40426 7055 40455 7059
rect 40365 7047 40455 7055
rect 40365 6995 40383 7047
rect 40435 6995 40455 7047
rect 40365 6983 40392 6995
rect 40426 6983 40455 6995
rect 40365 6931 40383 6983
rect 40435 6931 40455 6983
rect 40365 6918 40392 6931
rect 40128 6873 40174 6911
rect 40128 6839 40134 6873
rect 40168 6839 40174 6873
rect 40128 6801 40174 6839
rect 40128 6767 40134 6801
rect 40168 6767 40174 6801
rect 40128 6729 40174 6767
rect 40128 6695 40134 6729
rect 40168 6695 40174 6729
rect 40128 6657 40174 6695
rect 40128 6651 40134 6657
rect 39870 6585 39916 6623
rect 39870 6551 39876 6585
rect 39910 6551 39916 6585
rect 39870 6513 39916 6551
rect 39870 6479 39876 6513
rect 39910 6479 39916 6513
rect 39354 6407 39360 6441
rect 39394 6407 39400 6441
rect 39354 6369 39400 6407
rect 39354 6335 39360 6369
rect 39394 6335 39400 6369
rect 39354 6288 39400 6335
rect 39612 6441 39658 6443
rect 39612 6407 39618 6441
rect 39652 6407 39658 6441
rect 39612 6369 39658 6407
rect 39612 6335 39618 6369
rect 39652 6335 39658 6369
rect 39612 6288 39658 6335
rect 39870 6441 39916 6479
rect 40109 6636 40134 6651
rect 40168 6651 40174 6657
rect 40386 6911 40392 6918
rect 40426 6918 40455 6931
rect 40644 7089 40690 7127
rect 40902 8241 40948 8288
rect 40902 8207 40908 8241
rect 40942 8207 40948 8241
rect 40902 8169 40948 8207
rect 40902 8135 40908 8169
rect 40942 8135 40948 8169
rect 40902 8097 40948 8135
rect 40902 8063 40908 8097
rect 40942 8063 40948 8097
rect 40902 8025 40948 8063
rect 40902 7991 40908 8025
rect 40942 7991 40948 8025
rect 40902 7953 40948 7991
rect 40902 7919 40908 7953
rect 40942 7919 40948 7953
rect 40902 7881 40948 7919
rect 40902 7847 40908 7881
rect 40942 7847 40948 7881
rect 40902 7809 40948 7847
rect 40902 7775 40908 7809
rect 40942 7775 40948 7809
rect 40902 7737 40948 7775
rect 40902 7703 40908 7737
rect 40942 7703 40948 7737
rect 40902 7665 40948 7703
rect 40902 7631 40908 7665
rect 40942 7631 40948 7665
rect 40902 7593 40948 7631
rect 40902 7559 40908 7593
rect 40942 7559 40948 7593
rect 40902 7521 40948 7559
rect 40902 7487 40908 7521
rect 40942 7487 40948 7521
rect 40902 7449 40948 7487
rect 40902 7415 40908 7449
rect 40942 7415 40948 7449
rect 40902 7377 40948 7415
rect 40902 7343 40908 7377
rect 40942 7343 40948 7377
rect 40902 7305 40948 7343
rect 40902 7271 40908 7305
rect 40942 7271 40948 7305
rect 40902 7233 40948 7271
rect 40902 7199 40908 7233
rect 40942 7199 40948 7233
rect 40902 7161 40948 7199
rect 40902 7127 40908 7161
rect 40942 7127 40948 7161
rect 40902 7125 40948 7127
rect 41160 8241 41206 8288
rect 41160 8207 41166 8241
rect 41200 8207 41206 8241
rect 41160 8169 41206 8207
rect 41160 8135 41166 8169
rect 41200 8135 41206 8169
rect 41160 8097 41206 8135
rect 41160 8063 41166 8097
rect 41200 8063 41206 8097
rect 41160 8025 41206 8063
rect 41160 7991 41166 8025
rect 41200 7991 41206 8025
rect 41160 7953 41206 7991
rect 41160 7919 41166 7953
rect 41200 7919 41206 7953
rect 41160 7881 41206 7919
rect 41160 7847 41166 7881
rect 41200 7847 41206 7881
rect 41160 7809 41206 7847
rect 41160 7775 41166 7809
rect 41200 7775 41206 7809
rect 41160 7737 41206 7775
rect 41160 7703 41166 7737
rect 41200 7703 41206 7737
rect 41160 7665 41206 7703
rect 41160 7631 41166 7665
rect 41200 7631 41206 7665
rect 41160 7593 41206 7631
rect 41160 7559 41166 7593
rect 41200 7559 41206 7593
rect 41418 8241 41464 8288
rect 41418 8207 41424 8241
rect 41458 8207 41464 8241
rect 41418 8169 41464 8207
rect 41418 8135 41424 8169
rect 41458 8135 41464 8169
rect 41418 8097 41464 8135
rect 41418 8063 41424 8097
rect 41458 8063 41464 8097
rect 41418 8025 41464 8063
rect 41418 7991 41424 8025
rect 41458 7991 41464 8025
rect 41418 7953 41464 7991
rect 41418 7919 41424 7953
rect 41458 7919 41464 7953
rect 41418 7881 41464 7919
rect 41418 7847 41424 7881
rect 41458 7847 41464 7881
rect 41418 7809 41464 7847
rect 41418 7775 41424 7809
rect 41458 7775 41464 7809
rect 41418 7737 41464 7775
rect 41418 7703 41424 7737
rect 41458 7703 41464 7737
rect 41418 7665 41464 7703
rect 41418 7631 41424 7665
rect 41458 7631 41464 7665
rect 41418 7593 41464 7631
rect 41418 7561 41424 7593
rect 41160 7521 41206 7559
rect 41160 7487 41166 7521
rect 41200 7487 41206 7521
rect 41160 7449 41206 7487
rect 41160 7415 41166 7449
rect 41200 7415 41206 7449
rect 41160 7377 41206 7415
rect 41160 7343 41166 7377
rect 41200 7343 41206 7377
rect 41398 7559 41424 7561
rect 41458 7561 41464 7593
rect 41676 8241 41722 8288
rect 41676 8207 41682 8241
rect 41716 8207 41722 8241
rect 41676 8169 41722 8207
rect 41676 8135 41682 8169
rect 41716 8135 41722 8169
rect 41676 8097 41722 8135
rect 41676 8063 41682 8097
rect 41716 8063 41722 8097
rect 41676 8025 41722 8063
rect 41676 7991 41682 8025
rect 41716 7991 41722 8025
rect 41676 7953 41722 7991
rect 41676 7919 41682 7953
rect 41716 7919 41722 7953
rect 41676 7881 41722 7919
rect 41676 7847 41682 7881
rect 41716 7847 41722 7881
rect 41676 7809 41722 7847
rect 41676 7775 41682 7809
rect 41716 7775 41722 7809
rect 41676 7737 41722 7775
rect 41676 7703 41682 7737
rect 41716 7703 41722 7737
rect 41676 7665 41722 7703
rect 41676 7631 41682 7665
rect 41716 7631 41722 7665
rect 41676 7593 41722 7631
rect 41458 7559 41488 7561
rect 41398 7521 41488 7559
rect 41398 7514 41424 7521
rect 41458 7514 41488 7521
rect 41398 7462 41417 7514
rect 41469 7462 41488 7514
rect 41398 7450 41488 7462
rect 41398 7398 41417 7450
rect 41469 7398 41488 7450
rect 41398 7377 41488 7398
rect 41398 7356 41424 7377
rect 41160 7305 41206 7343
rect 41160 7271 41166 7305
rect 41200 7271 41206 7305
rect 41160 7233 41206 7271
rect 41160 7199 41166 7233
rect 41200 7199 41206 7233
rect 41160 7161 41206 7199
rect 41160 7127 41166 7161
rect 41200 7127 41206 7161
rect 40644 7055 40650 7089
rect 40684 7055 40690 7089
rect 40644 7017 40690 7055
rect 40644 6983 40650 7017
rect 40684 6983 40690 7017
rect 40644 6945 40690 6983
rect 40426 6911 40432 6918
rect 40386 6873 40432 6911
rect 40386 6839 40392 6873
rect 40426 6839 40432 6873
rect 40386 6801 40432 6839
rect 40386 6767 40392 6801
rect 40426 6767 40432 6801
rect 40386 6729 40432 6767
rect 40386 6695 40392 6729
rect 40426 6695 40432 6729
rect 40386 6657 40432 6695
rect 40168 6636 40193 6651
rect 40109 6584 40125 6636
rect 40177 6584 40193 6636
rect 40109 6572 40134 6584
rect 40168 6572 40193 6584
rect 40109 6520 40125 6572
rect 40177 6520 40193 6572
rect 40109 6513 40193 6520
rect 40109 6508 40134 6513
rect 40168 6508 40193 6513
rect 40109 6456 40125 6508
rect 40177 6456 40193 6508
rect 40109 6443 40193 6456
rect 40386 6623 40392 6657
rect 40426 6623 40432 6657
rect 40644 6911 40650 6945
rect 40684 6911 40690 6945
rect 40884 7109 40967 7125
rect 40884 7057 40898 7109
rect 40950 7057 40967 7109
rect 40884 7055 40908 7057
rect 40942 7055 40967 7057
rect 40884 7045 40967 7055
rect 40884 6993 40898 7045
rect 40950 6993 40967 7045
rect 40884 6983 40908 6993
rect 40942 6983 40967 6993
rect 40884 6981 40967 6983
rect 40884 6929 40898 6981
rect 40950 6929 40967 6981
rect 40884 6918 40908 6929
rect 40644 6873 40690 6911
rect 40644 6839 40650 6873
rect 40684 6839 40690 6873
rect 40644 6801 40690 6839
rect 40644 6767 40650 6801
rect 40684 6767 40690 6801
rect 40644 6729 40690 6767
rect 40644 6695 40650 6729
rect 40684 6695 40690 6729
rect 40644 6657 40690 6695
rect 40644 6651 40650 6657
rect 40386 6585 40432 6623
rect 40386 6551 40392 6585
rect 40426 6551 40432 6585
rect 40386 6513 40432 6551
rect 40386 6479 40392 6513
rect 40426 6479 40432 6513
rect 39870 6407 39876 6441
rect 39910 6407 39916 6441
rect 39870 6369 39916 6407
rect 39870 6335 39876 6369
rect 39910 6335 39916 6369
rect 39870 6288 39916 6335
rect 40128 6441 40174 6443
rect 40128 6407 40134 6441
rect 40168 6407 40174 6441
rect 40128 6369 40174 6407
rect 40128 6335 40134 6369
rect 40168 6335 40174 6369
rect 40128 6288 40174 6335
rect 40386 6441 40432 6479
rect 40627 6637 40650 6651
rect 40684 6651 40690 6657
rect 40902 6911 40908 6918
rect 40942 6918 40967 6929
rect 41160 7089 41206 7127
rect 41160 7055 41166 7089
rect 41200 7055 41206 7089
rect 41160 7017 41206 7055
rect 41160 6983 41166 7017
rect 41200 6983 41206 7017
rect 41160 6945 41206 6983
rect 40942 6911 40948 6918
rect 40902 6873 40948 6911
rect 40902 6839 40908 6873
rect 40942 6839 40948 6873
rect 40902 6801 40948 6839
rect 40902 6767 40908 6801
rect 40942 6767 40948 6801
rect 40902 6729 40948 6767
rect 40902 6695 40908 6729
rect 40942 6695 40948 6729
rect 40902 6657 40948 6695
rect 40684 6637 40707 6651
rect 40627 6585 40640 6637
rect 40692 6585 40707 6637
rect 40627 6573 40650 6585
rect 40684 6573 40707 6585
rect 40627 6521 40640 6573
rect 40692 6521 40707 6573
rect 40627 6513 40707 6521
rect 40627 6509 40650 6513
rect 40684 6509 40707 6513
rect 40627 6457 40640 6509
rect 40692 6457 40707 6509
rect 40627 6443 40707 6457
rect 40902 6623 40908 6657
rect 40942 6623 40948 6657
rect 41160 6911 41166 6945
rect 41200 6911 41206 6945
rect 41160 6873 41206 6911
rect 41160 6839 41166 6873
rect 41200 6839 41206 6873
rect 41160 6801 41206 6839
rect 41160 6767 41166 6801
rect 41200 6767 41206 6801
rect 41160 6729 41206 6767
rect 41160 6695 41166 6729
rect 41200 6695 41206 6729
rect 41160 6657 41206 6695
rect 41160 6651 41166 6657
rect 40902 6585 40948 6623
rect 40902 6551 40908 6585
rect 40942 6551 40948 6585
rect 40902 6513 40948 6551
rect 40902 6479 40908 6513
rect 40942 6479 40948 6513
rect 40386 6407 40392 6441
rect 40426 6407 40432 6441
rect 40386 6369 40432 6407
rect 40386 6335 40392 6369
rect 40426 6335 40432 6369
rect 40386 6288 40432 6335
rect 40644 6441 40690 6443
rect 40644 6407 40650 6441
rect 40684 6407 40690 6441
rect 40644 6369 40690 6407
rect 40644 6335 40650 6369
rect 40684 6335 40690 6369
rect 40644 6288 40690 6335
rect 40902 6441 40948 6479
rect 41143 6637 41166 6651
rect 41200 6651 41206 6657
rect 41418 7343 41424 7356
rect 41458 7356 41488 7377
rect 41676 7559 41682 7593
rect 41716 7559 41722 7593
rect 41934 8241 41980 8288
rect 41934 8207 41940 8241
rect 41974 8207 41980 8241
rect 41934 8169 41980 8207
rect 41934 8135 41940 8169
rect 41974 8135 41980 8169
rect 41934 8097 41980 8135
rect 41934 8063 41940 8097
rect 41974 8063 41980 8097
rect 41934 8025 41980 8063
rect 41934 7991 41940 8025
rect 41974 7991 41980 8025
rect 41934 7953 41980 7991
rect 41934 7919 41940 7953
rect 41974 7919 41980 7953
rect 41934 7881 41980 7919
rect 41934 7847 41940 7881
rect 41974 7847 41980 7881
rect 41934 7809 41980 7847
rect 41934 7775 41940 7809
rect 41974 7775 41980 7809
rect 41934 7737 41980 7775
rect 41934 7703 41940 7737
rect 41974 7703 41980 7737
rect 41934 7665 41980 7703
rect 43358 7779 43495 9815
rect 44507 7779 44648 9815
rect 43358 7672 44648 7779
rect 41934 7631 41940 7665
rect 41974 7631 41980 7665
rect 41934 7593 41980 7631
rect 41934 7561 41940 7593
rect 41676 7521 41722 7559
rect 41676 7487 41682 7521
rect 41716 7487 41722 7521
rect 41676 7449 41722 7487
rect 41676 7415 41682 7449
rect 41716 7415 41722 7449
rect 41676 7377 41722 7415
rect 41458 7343 41464 7356
rect 41418 7305 41464 7343
rect 41418 7271 41424 7305
rect 41458 7271 41464 7305
rect 41418 7233 41464 7271
rect 41418 7199 41424 7233
rect 41458 7199 41464 7233
rect 41418 7161 41464 7199
rect 41418 7127 41424 7161
rect 41458 7127 41464 7161
rect 41418 7089 41464 7127
rect 41418 7055 41424 7089
rect 41458 7055 41464 7089
rect 41418 7017 41464 7055
rect 41418 6983 41424 7017
rect 41458 6983 41464 7017
rect 41418 6945 41464 6983
rect 41418 6911 41424 6945
rect 41458 6911 41464 6945
rect 41418 6873 41464 6911
rect 41418 6839 41424 6873
rect 41458 6839 41464 6873
rect 41418 6801 41464 6839
rect 41418 6767 41424 6801
rect 41458 6767 41464 6801
rect 41418 6729 41464 6767
rect 41418 6695 41424 6729
rect 41458 6695 41464 6729
rect 41418 6657 41464 6695
rect 41200 6637 41222 6651
rect 41143 6585 41157 6637
rect 41209 6585 41222 6637
rect 41143 6573 41166 6585
rect 41200 6573 41222 6585
rect 41143 6521 41157 6573
rect 41209 6521 41222 6573
rect 41143 6513 41222 6521
rect 41143 6509 41166 6513
rect 41200 6509 41222 6513
rect 41143 6457 41157 6509
rect 41209 6457 41222 6509
rect 41143 6443 41222 6457
rect 41418 6623 41424 6657
rect 41458 6623 41464 6657
rect 41676 7343 41682 7377
rect 41716 7343 41722 7377
rect 41917 7559 41940 7561
rect 41974 7561 41980 7593
rect 41974 7559 41996 7561
rect 41917 7548 41996 7559
rect 41917 7496 41930 7548
rect 41982 7496 41996 7548
rect 41917 7487 41940 7496
rect 41974 7487 41996 7496
rect 41917 7484 41996 7487
rect 41917 7432 41930 7484
rect 41982 7432 41996 7484
rect 41917 7420 41940 7432
rect 41974 7420 41996 7432
rect 41917 7368 41930 7420
rect 41982 7368 41996 7420
rect 41917 7356 41940 7368
rect 41676 7305 41722 7343
rect 41676 7271 41682 7305
rect 41716 7271 41722 7305
rect 41676 7233 41722 7271
rect 41676 7199 41682 7233
rect 41716 7199 41722 7233
rect 41676 7161 41722 7199
rect 41676 7127 41682 7161
rect 41716 7127 41722 7161
rect 41676 7089 41722 7127
rect 41676 7055 41682 7089
rect 41716 7055 41722 7089
rect 41676 7017 41722 7055
rect 41676 6983 41682 7017
rect 41716 6983 41722 7017
rect 41676 6945 41722 6983
rect 41676 6911 41682 6945
rect 41716 6911 41722 6945
rect 41676 6873 41722 6911
rect 41676 6839 41682 6873
rect 41716 6839 41722 6873
rect 41676 6801 41722 6839
rect 41676 6767 41682 6801
rect 41716 6767 41722 6801
rect 41676 6729 41722 6767
rect 41676 6695 41682 6729
rect 41716 6695 41722 6729
rect 41676 6657 41722 6695
rect 41676 6651 41682 6657
rect 41418 6585 41464 6623
rect 41418 6551 41424 6585
rect 41458 6551 41464 6585
rect 41418 6513 41464 6551
rect 41418 6479 41424 6513
rect 41458 6479 41464 6513
rect 40902 6407 40908 6441
rect 40942 6407 40948 6441
rect 40902 6369 40948 6407
rect 40902 6335 40908 6369
rect 40942 6335 40948 6369
rect 40902 6288 40948 6335
rect 41160 6441 41206 6443
rect 41160 6407 41166 6441
rect 41200 6407 41206 6441
rect 41160 6369 41206 6407
rect 41160 6335 41166 6369
rect 41200 6335 41206 6369
rect 41160 6288 41206 6335
rect 41418 6441 41464 6479
rect 41660 6637 41682 6651
rect 41716 6651 41722 6657
rect 41934 7343 41940 7356
rect 41974 7356 41996 7368
rect 41974 7343 41980 7356
rect 41934 7305 41980 7343
rect 41934 7271 41940 7305
rect 41974 7271 41980 7305
rect 41934 7233 41980 7271
rect 41934 7199 41940 7233
rect 41974 7199 41980 7233
rect 41934 7161 41980 7199
rect 41934 7127 41940 7161
rect 41974 7127 41980 7161
rect 41934 7089 41980 7127
rect 41934 7055 41940 7089
rect 41974 7055 41980 7089
rect 41934 7017 41980 7055
rect 41934 6983 41940 7017
rect 41974 6983 41980 7017
rect 41934 6945 41980 6983
rect 41934 6911 41940 6945
rect 41974 6911 41980 6945
rect 41934 6873 41980 6911
rect 41934 6839 41940 6873
rect 41974 6839 41980 6873
rect 41934 6801 41980 6839
rect 41934 6767 41940 6801
rect 41974 6767 41980 6801
rect 41934 6729 41980 6767
rect 41934 6695 41940 6729
rect 41974 6695 41980 6729
rect 41934 6657 41980 6695
rect 41716 6637 41740 6651
rect 41660 6585 41673 6637
rect 41725 6585 41740 6637
rect 41660 6573 41682 6585
rect 41716 6573 41740 6585
rect 41660 6521 41673 6573
rect 41725 6521 41740 6573
rect 41660 6513 41740 6521
rect 41660 6509 41682 6513
rect 41716 6509 41740 6513
rect 41660 6457 41673 6509
rect 41725 6457 41740 6509
rect 41660 6443 41740 6457
rect 41934 6623 41940 6657
rect 41974 6623 41980 6657
rect 41934 6585 41980 6623
rect 41934 6551 41940 6585
rect 41974 6551 41980 6585
rect 41934 6513 41980 6551
rect 41934 6479 41940 6513
rect 41974 6479 41980 6513
rect 41418 6407 41424 6441
rect 41458 6407 41464 6441
rect 41418 6369 41464 6407
rect 41418 6335 41424 6369
rect 41458 6335 41464 6369
rect 41418 6288 41464 6335
rect 41676 6441 41722 6443
rect 41676 6407 41682 6441
rect 41716 6407 41722 6441
rect 41676 6369 41722 6407
rect 41676 6335 41682 6369
rect 41716 6335 41722 6369
rect 41676 6288 41722 6335
rect 41934 6441 41980 6479
rect 42104 6635 42208 6651
rect 42104 6583 42127 6635
rect 42179 6583 42208 6635
rect 42104 6571 42208 6583
rect 42104 6519 42127 6571
rect 42179 6519 42208 6571
rect 42104 6507 42208 6519
rect 42104 6455 42127 6507
rect 42179 6455 42208 6507
rect 42104 6442 42208 6455
rect 41934 6407 41940 6441
rect 41974 6407 41980 6441
rect 41934 6369 41980 6407
rect 41934 6335 41940 6369
rect 41974 6335 41980 6369
rect 41934 6288 41980 6335
rect 37806 6250 38054 6256
rect 37806 6216 37905 6250
rect 37939 6216 37977 6250
rect 38011 6216 38054 6250
rect 37806 6210 38054 6216
rect 38120 6250 38312 6256
rect 38120 6216 38163 6250
rect 38197 6216 38235 6250
rect 38269 6216 38312 6250
rect 38120 6210 38312 6216
rect 38378 6250 38570 6256
rect 38378 6216 38421 6250
rect 38455 6216 38493 6250
rect 38527 6216 38570 6250
rect 38378 6210 38570 6216
rect 37806 6200 38570 6210
rect 38636 6250 38828 6256
rect 38636 6216 38679 6250
rect 38713 6216 38751 6250
rect 38785 6216 38828 6250
rect 38636 6210 38828 6216
rect 38894 6250 39086 6256
rect 38894 6216 38937 6250
rect 38971 6216 39009 6250
rect 39043 6216 39086 6250
rect 38894 6210 39086 6216
rect 39152 6250 39344 6256
rect 39152 6216 39195 6250
rect 39229 6216 39267 6250
rect 39301 6216 39344 6250
rect 39152 6210 39344 6216
rect 39410 6250 39602 6256
rect 39410 6216 39453 6250
rect 39487 6216 39525 6250
rect 39559 6216 39602 6250
rect 39410 6210 39602 6216
rect 39668 6250 39860 6256
rect 39668 6216 39711 6250
rect 39745 6216 39783 6250
rect 39817 6216 39860 6250
rect 39668 6210 39860 6216
rect 39926 6250 40118 6256
rect 39926 6216 39969 6250
rect 40003 6216 40041 6250
rect 40075 6216 40118 6250
rect 39926 6210 40118 6216
rect 40184 6250 40376 6256
rect 40184 6216 40227 6250
rect 40261 6216 40299 6250
rect 40333 6216 40376 6250
rect 40184 6210 40376 6216
rect 40442 6250 40634 6256
rect 40442 6216 40485 6250
rect 40519 6216 40557 6250
rect 40591 6216 40634 6250
rect 40442 6210 40634 6216
rect 40700 6250 40892 6256
rect 40700 6216 40743 6250
rect 40777 6216 40815 6250
rect 40849 6216 40892 6250
rect 40700 6210 40892 6216
rect 40958 6250 41150 6256
rect 40958 6216 41001 6250
rect 41035 6216 41073 6250
rect 41107 6216 41150 6250
rect 40958 6210 41150 6216
rect 38636 6200 41150 6210
rect 41216 6250 41408 6256
rect 41216 6216 41259 6250
rect 41293 6216 41331 6250
rect 41365 6216 41408 6250
rect 41216 6210 41408 6216
rect 41474 6250 41666 6256
rect 41474 6216 41517 6250
rect 41551 6216 41589 6250
rect 41623 6216 41666 6250
rect 41474 6210 41666 6216
rect 41732 6250 41924 6256
rect 41732 6216 41775 6250
rect 41809 6216 41847 6250
rect 41881 6216 41924 6250
rect 41732 6210 41924 6216
rect 41216 6200 41924 6210
rect 37806 6146 41924 6200
rect 26142 6077 26188 6115
rect 26142 6043 26148 6077
rect 26182 6043 26188 6077
rect 26142 6005 26188 6043
rect 26142 5971 26148 6005
rect 26182 5971 26188 6005
rect 26142 5933 26188 5971
rect 26142 5899 26148 5933
rect 26182 5899 26188 5933
rect 26142 5861 26188 5899
rect 26142 5827 26148 5861
rect 26182 5852 26188 5861
rect 26182 5827 26222 5852
rect 25002 5714 25032 5780
rect 25142 5770 25302 5792
rect 26142 5780 26222 5827
rect 25110 5764 26110 5770
rect 25110 5730 25125 5764
rect 25159 5758 25197 5764
rect 25231 5758 25269 5764
rect 25303 5730 25341 5764
rect 25375 5730 25413 5764
rect 25447 5730 25485 5764
rect 25519 5730 25557 5764
rect 25591 5730 25629 5764
rect 25663 5730 25701 5764
rect 25735 5730 25773 5764
rect 25807 5730 25845 5764
rect 25879 5730 25917 5764
rect 25951 5730 25989 5764
rect 26023 5730 26061 5764
rect 26095 5730 26110 5764
rect 25110 5724 25159 5730
rect 25002 5667 25078 5714
rect 25142 5706 25159 5724
rect 25211 5706 25223 5730
rect 25275 5724 26110 5730
rect 25275 5706 25302 5724
rect 26182 5714 26222 5780
rect 25142 5682 25302 5706
rect 25002 5662 25038 5667
rect 24682 5633 24688 5652
rect 24642 5595 24688 5633
rect 24642 5561 24648 5595
rect 24682 5561 24688 5595
rect 24642 5523 24688 5561
rect 24642 5489 24648 5523
rect 24682 5489 24688 5523
rect 24642 5451 24688 5489
rect 24642 5417 24648 5451
rect 24682 5417 24688 5451
rect 24642 5379 24688 5417
rect 24642 5345 24648 5379
rect 24682 5345 24688 5379
rect 24642 5307 24688 5345
rect 24642 5273 24648 5307
rect 24682 5273 24688 5307
rect 24642 5235 24688 5273
rect 24642 5201 24648 5235
rect 24682 5201 24688 5235
rect 24642 5163 24688 5201
rect 24642 5129 24648 5163
rect 24682 5129 24688 5163
rect 24642 5091 24688 5129
rect 24642 5057 24648 5091
rect 24682 5057 24688 5091
rect 24642 5019 24688 5057
rect 24642 4985 24648 5019
rect 24682 4985 24688 5019
rect 24642 4947 24688 4985
rect 24642 4913 24648 4947
rect 24682 4913 24688 4947
rect 24642 4875 24688 4913
rect 24642 4841 24648 4875
rect 24682 4841 24688 4875
rect 24642 4803 24688 4841
rect 24642 4769 24648 4803
rect 24682 4772 24688 4803
rect 25032 5633 25038 5662
rect 25072 5633 25078 5667
rect 25032 5595 25078 5633
rect 25032 5561 25038 5595
rect 25072 5561 25078 5595
rect 25032 5523 25078 5561
rect 25032 5489 25038 5523
rect 25072 5489 25078 5523
rect 25032 5451 25078 5489
rect 25032 5417 25038 5451
rect 25072 5417 25078 5451
rect 25032 5379 25078 5417
rect 25032 5345 25038 5379
rect 25072 5345 25078 5379
rect 25032 5307 25078 5345
rect 25032 5273 25038 5307
rect 25072 5273 25078 5307
rect 25032 5235 25078 5273
rect 25032 5201 25038 5235
rect 25072 5201 25078 5235
rect 25032 5163 25078 5201
rect 25032 5129 25038 5163
rect 25072 5129 25078 5163
rect 25032 5091 25078 5129
rect 25032 5057 25038 5091
rect 25072 5057 25078 5091
rect 25032 5019 25078 5057
rect 25032 4985 25038 5019
rect 25072 4985 25078 5019
rect 25032 4947 25078 4985
rect 25032 4913 25038 4947
rect 25072 4913 25078 4947
rect 25032 4875 25078 4913
rect 25032 4841 25038 4875
rect 25072 4841 25078 4875
rect 25032 4803 25078 4841
rect 25032 4782 25038 4803
rect 24682 4769 24712 4772
rect 24362 4743 24522 4762
rect 23502 4656 23532 4722
rect 24362 4712 24379 4743
rect 23610 4706 24379 4712
rect 24431 4706 24443 4743
rect 24495 4712 24522 4743
rect 24642 4722 24712 4769
rect 24495 4706 24610 4712
rect 23610 4672 23625 4706
rect 23659 4672 23697 4706
rect 23731 4672 23769 4706
rect 23803 4672 23841 4706
rect 23875 4672 23913 4706
rect 23947 4672 23985 4706
rect 24019 4672 24057 4706
rect 24091 4672 24129 4706
rect 24163 4672 24201 4706
rect 24235 4672 24273 4706
rect 24307 4672 24345 4706
rect 24379 4672 24417 4691
rect 24451 4672 24489 4691
rect 24523 4672 24561 4706
rect 24595 4672 24610 4706
rect 23610 4666 24610 4672
rect 24682 4656 24712 4722
rect 23502 4609 23578 4656
rect 23502 4592 23538 4609
rect 19936 4548 19982 4591
rect 23532 4575 23538 4592
rect 23572 4575 23578 4609
rect 23532 4537 23578 4575
rect 17484 4510 18476 4516
rect 18934 4510 19926 4516
rect 17484 4476 17531 4510
rect 17565 4476 17603 4510
rect 17637 4476 17675 4510
rect 17709 4476 17747 4510
rect 17781 4476 17819 4510
rect 17853 4476 17891 4510
rect 17925 4476 17963 4510
rect 17997 4476 18035 4510
rect 18069 4476 18107 4510
rect 18141 4476 18179 4510
rect 18213 4476 18251 4510
rect 18285 4476 18323 4510
rect 18357 4476 18395 4510
rect 18429 4476 18981 4510
rect 19015 4476 19053 4510
rect 19087 4476 19125 4510
rect 19159 4476 19197 4510
rect 19231 4476 19269 4510
rect 19303 4476 19341 4510
rect 19375 4476 19413 4510
rect 19447 4476 19485 4510
rect 19519 4476 19557 4510
rect 19591 4476 19629 4510
rect 19663 4476 19701 4510
rect 19735 4476 19773 4510
rect 19807 4476 19845 4510
rect 19879 4476 19926 4510
rect 17484 4470 19926 4476
rect 23532 4503 23538 4537
rect 23572 4503 23578 4537
rect 18392 4440 19012 4470
rect 23532 4465 23578 4503
rect 23532 4431 23538 4465
rect 23572 4431 23578 4465
rect 23532 4393 23578 4431
rect 23532 4359 23538 4393
rect 23572 4359 23578 4393
rect 23532 4321 23578 4359
rect 12752 4230 22752 4306
rect 12752 4209 12847 4230
rect 22627 4209 22752 4230
rect 12752 3815 12824 4209
rect 22650 3815 22752 4209
rect 12752 3794 12847 3815
rect 22627 3794 22752 3815
rect 12752 3730 22752 3794
rect 23532 4287 23538 4321
rect 23572 4287 23578 4321
rect 23532 4249 23578 4287
rect 23532 4215 23538 4249
rect 23572 4215 23578 4249
rect 23532 4177 23578 4215
rect 23532 4143 23538 4177
rect 23572 4143 23578 4177
rect 23532 4105 23578 4143
rect 23532 4071 23538 4105
rect 23572 4071 23578 4105
rect 23532 4033 23578 4071
rect 23532 3999 23538 4033
rect 23572 3999 23578 4033
rect 23532 3961 23578 3999
rect 23532 3927 23538 3961
rect 23572 3927 23578 3961
rect 23532 3889 23578 3927
rect 23532 3855 23538 3889
rect 23572 3855 23578 3889
rect 23532 3817 23578 3855
rect 23532 3783 23538 3817
rect 23572 3783 23578 3817
rect 23532 3745 23578 3783
rect 23532 3711 23538 3745
rect 23572 3711 23578 3745
rect 23532 3664 23578 3711
rect 24642 4609 24712 4656
rect 24642 4575 24648 4609
rect 24682 4582 24712 4609
rect 25002 4769 25038 4782
rect 25072 4769 25078 4803
rect 26142 5667 26222 5714
rect 26142 5633 26148 5667
rect 26182 5662 26222 5667
rect 26182 5633 26188 5662
rect 26142 5595 26188 5633
rect 26142 5561 26148 5595
rect 26182 5561 26188 5595
rect 26142 5523 26188 5561
rect 26142 5489 26148 5523
rect 26182 5489 26188 5523
rect 26142 5451 26188 5489
rect 26142 5417 26148 5451
rect 26182 5417 26188 5451
rect 26142 5379 26188 5417
rect 26142 5345 26148 5379
rect 26182 5345 26188 5379
rect 26142 5307 26188 5345
rect 26142 5273 26148 5307
rect 26182 5273 26188 5307
rect 26142 5235 26188 5273
rect 26142 5201 26148 5235
rect 26182 5201 26188 5235
rect 26142 5163 26188 5201
rect 26142 5129 26148 5163
rect 26182 5129 26188 5163
rect 26142 5091 26188 5129
rect 26142 5057 26148 5091
rect 26182 5057 26188 5091
rect 26142 5019 26188 5057
rect 26142 4985 26148 5019
rect 26182 4985 26188 5019
rect 26142 4947 26188 4985
rect 26142 4913 26148 4947
rect 26182 4913 26188 4947
rect 26142 4875 26188 4913
rect 26142 4841 26148 4875
rect 26182 4841 26188 4875
rect 26142 4803 26188 4841
rect 25002 4722 25078 4769
rect 25852 4753 26012 4802
rect 25002 4656 25042 4722
rect 25852 4712 25869 4753
rect 25110 4706 25869 4712
rect 25921 4706 25933 4753
rect 25985 4712 26012 4753
rect 26142 4769 26148 4803
rect 26182 4792 26188 4803
rect 26182 4769 26212 4792
rect 26142 4722 26212 4769
rect 25985 4706 26110 4712
rect 25110 4672 25125 4706
rect 25159 4672 25197 4706
rect 25231 4672 25269 4706
rect 25303 4672 25341 4706
rect 25375 4672 25413 4706
rect 25447 4672 25485 4706
rect 25519 4672 25557 4706
rect 25591 4672 25629 4706
rect 25663 4672 25701 4706
rect 25735 4672 25773 4706
rect 25807 4672 25845 4706
rect 25985 4701 25989 4706
rect 25879 4672 25917 4701
rect 25951 4672 25989 4701
rect 26023 4672 26061 4706
rect 26095 4672 26110 4706
rect 25110 4666 26110 4672
rect 26182 4656 26212 4722
rect 25002 4609 25078 4656
rect 25002 4592 25038 4609
rect 24682 4575 24688 4582
rect 24642 4537 24688 4575
rect 24642 4503 24648 4537
rect 24682 4503 24688 4537
rect 24642 4465 24688 4503
rect 24642 4431 24648 4465
rect 24682 4431 24688 4465
rect 24642 4393 24688 4431
rect 24642 4359 24648 4393
rect 24682 4359 24688 4393
rect 24642 4321 24688 4359
rect 24642 4287 24648 4321
rect 24682 4287 24688 4321
rect 24642 4249 24688 4287
rect 24642 4215 24648 4249
rect 24682 4215 24688 4249
rect 24642 4177 24688 4215
rect 24642 4143 24648 4177
rect 24682 4143 24688 4177
rect 24642 4105 24688 4143
rect 24642 4071 24648 4105
rect 24682 4071 24688 4105
rect 24642 4033 24688 4071
rect 24642 3999 24648 4033
rect 24682 3999 24688 4033
rect 24642 3961 24688 3999
rect 24642 3927 24648 3961
rect 24682 3927 24688 3961
rect 24642 3889 24688 3927
rect 24642 3855 24648 3889
rect 24682 3855 24688 3889
rect 24642 3817 24688 3855
rect 24642 3783 24648 3817
rect 24682 3783 24688 3817
rect 24642 3745 24688 3783
rect 24642 3711 24648 3745
rect 24682 3711 24688 3745
rect 23642 3678 23812 3692
rect 23642 3654 23669 3678
rect 23610 3648 23669 3654
rect 23721 3648 23733 3678
rect 23785 3654 23812 3678
rect 24642 3664 24688 3711
rect 25032 4575 25038 4592
rect 25072 4575 25078 4609
rect 25032 4537 25078 4575
rect 25032 4503 25038 4537
rect 25072 4503 25078 4537
rect 25032 4465 25078 4503
rect 25032 4431 25038 4465
rect 25072 4431 25078 4465
rect 25032 4393 25078 4431
rect 25032 4359 25038 4393
rect 25072 4359 25078 4393
rect 25032 4321 25078 4359
rect 25032 4287 25038 4321
rect 25072 4287 25078 4321
rect 25032 4249 25078 4287
rect 25032 4215 25038 4249
rect 25072 4215 25078 4249
rect 25032 4177 25078 4215
rect 25032 4143 25038 4177
rect 25072 4143 25078 4177
rect 25032 4105 25078 4143
rect 25032 4071 25038 4105
rect 25072 4071 25078 4105
rect 25032 4033 25078 4071
rect 25032 3999 25038 4033
rect 25072 3999 25078 4033
rect 25032 3961 25078 3999
rect 25032 3927 25038 3961
rect 25072 3927 25078 3961
rect 25032 3889 25078 3927
rect 25032 3855 25038 3889
rect 25072 3855 25078 3889
rect 25032 3817 25078 3855
rect 25032 3783 25038 3817
rect 25072 3783 25078 3817
rect 25032 3745 25078 3783
rect 25032 3711 25038 3745
rect 25072 3711 25078 3745
rect 26142 4609 26212 4656
rect 26142 4575 26148 4609
rect 26182 4602 26212 4609
rect 26182 4575 26188 4602
rect 26142 4537 26188 4575
rect 26142 4503 26148 4537
rect 26182 4503 26188 4537
rect 26142 4465 26188 4503
rect 26142 4431 26148 4465
rect 26182 4431 26188 4465
rect 26142 4393 26188 4431
rect 26142 4359 26148 4393
rect 26182 4359 26188 4393
rect 26142 4321 26188 4359
rect 26142 4287 26148 4321
rect 26182 4287 26188 4321
rect 26142 4249 26188 4287
rect 26142 4215 26148 4249
rect 26182 4215 26188 4249
rect 26142 4177 26188 4215
rect 26142 4143 26148 4177
rect 26182 4143 26188 4177
rect 26142 4105 26188 4143
rect 26142 4071 26148 4105
rect 26182 4071 26188 4105
rect 26142 4033 26188 4071
rect 26142 3999 26148 4033
rect 26182 3999 26188 4033
rect 26142 3961 26188 3999
rect 26142 3927 26148 3961
rect 26182 3927 26188 3961
rect 26142 3889 26188 3927
rect 26142 3855 26148 3889
rect 26182 3855 26188 3889
rect 26142 3817 26188 3855
rect 26142 3783 26148 3817
rect 26182 3783 26188 3817
rect 26142 3745 26188 3783
rect 25032 3664 25078 3711
rect 25142 3678 25302 3722
rect 25142 3654 25164 3678
rect 23785 3648 24610 3654
rect 23610 3614 23625 3648
rect 23659 3626 23669 3648
rect 23731 3626 23733 3648
rect 23659 3614 23697 3626
rect 23731 3614 23769 3626
rect 23803 3614 23841 3648
rect 23875 3614 23913 3648
rect 23947 3614 23985 3648
rect 24019 3614 24057 3648
rect 24091 3614 24129 3648
rect 24163 3614 24201 3648
rect 24235 3614 24273 3648
rect 24307 3614 24345 3648
rect 24379 3614 24417 3648
rect 24451 3614 24489 3648
rect 24523 3614 24561 3648
rect 24595 3614 24610 3648
rect 23610 3608 24610 3614
rect 25110 3648 25164 3654
rect 25216 3648 25228 3678
rect 25280 3654 25302 3678
rect 26142 3711 26148 3745
rect 26182 3711 26188 3745
rect 26142 3664 26188 3711
rect 28320 3678 50460 3843
rect 25280 3648 26110 3654
rect 25110 3614 25125 3648
rect 25159 3626 25164 3648
rect 25159 3614 25197 3626
rect 25231 3614 25269 3626
rect 25303 3614 25341 3648
rect 25375 3614 25413 3648
rect 25447 3614 25485 3648
rect 25519 3614 25557 3648
rect 25591 3614 25629 3648
rect 25663 3614 25701 3648
rect 25735 3614 25773 3648
rect 25807 3614 25845 3648
rect 25879 3614 25917 3648
rect 25951 3614 25989 3648
rect 26023 3614 26061 3648
rect 26095 3614 26110 3648
rect 25110 3608 26110 3614
rect 24362 3513 24522 3552
rect 24362 3461 24384 3513
rect 24436 3461 24448 3513
rect 24500 3461 24522 3513
rect 24362 3422 24522 3461
rect 26538 3493 26588 3507
rect 26856 3502 26906 3507
rect 26538 3459 26546 3493
rect 26580 3459 26588 3493
rect 26538 3421 26588 3459
rect 26538 3387 26546 3421
rect 26580 3387 26588 3421
rect 26538 3349 26588 3387
rect 26538 3315 26546 3349
rect 26580 3315 26588 3349
rect 26538 3277 26588 3315
rect 26538 3243 26546 3277
rect 26580 3243 26588 3277
rect 26538 3205 26588 3243
rect 26538 3171 26546 3205
rect 26580 3171 26588 3205
rect 26538 3133 26588 3171
rect 26538 3099 26546 3133
rect 26580 3099 26588 3133
rect -13168 2928 11340 3093
rect 26538 3086 26588 3099
rect 26652 3493 27012 3502
rect 26652 3463 26864 3493
rect 26898 3463 27012 3493
rect 26652 3091 26705 3463
rect 26949 3091 27012 3463
rect 26652 3072 27012 3091
rect 27174 3493 27224 3507
rect 27174 3459 27182 3493
rect 27216 3459 27224 3493
rect 27174 3421 27224 3459
rect 27174 3387 27182 3421
rect 27216 3387 27224 3421
rect 27174 3349 27224 3387
rect 27174 3315 27182 3349
rect 27216 3315 27224 3349
rect 27174 3277 27224 3315
rect 27174 3243 27182 3277
rect 27216 3243 27224 3277
rect 27174 3205 27224 3243
rect 27174 3171 27182 3205
rect 27216 3171 27224 3205
rect 27174 3133 27224 3171
rect 27174 3099 27182 3133
rect 27216 3099 27224 3133
rect 27174 3086 27224 3099
rect -13168 2172 -13051 2928
rect -12039 2884 11340 2928
rect -12039 2192 3722 2884
rect 4734 2428 11340 2884
rect 28320 2922 32541 3678
rect 33553 3634 50460 3678
rect 33553 2942 49314 3634
rect 50326 2942 50460 3634
rect 33553 2922 50460 2942
rect 28320 2819 50460 2922
rect 28320 2428 29344 2819
rect 4734 2357 29346 2428
rect 4734 2192 10364 2357
rect -12039 2172 10364 2192
rect -13168 2069 10364 2172
rect 10296 1473 10364 2069
rect 11248 1473 29346 2357
rect 10296 1400 29346 1473
rect 30218 1537 52642 1673
rect 30218 1514 38612 1537
rect -15366 787 8992 923
rect -15366 764 -6980 787
rect -15366 8 -15192 764
rect -14308 8 -6980 764
rect -15366 -39 -6980 8
rect -5434 743 8992 787
rect -5434 51 5895 743
rect 6843 51 8992 743
rect 30218 758 30400 1514
rect 31284 758 38612 1514
rect 30218 711 38612 758
rect 40158 1493 52642 1537
rect 40158 801 51487 1493
rect 52435 801 52642 1493
rect 40158 711 52642 801
rect 30218 649 52642 711
rect -5434 -39 8992 51
rect -15366 -62 8992 -39
rect 30219 -62 31242 649
rect -15366 -96 31242 -62
rect -15366 -101 8106 -96
rect 7968 -1022 8106 -101
rect 8038 -1044 8106 -1022
rect 8990 -172 31242 -96
rect 8990 -992 12843 -172
rect 22623 -992 31242 -172
rect 8990 -1044 31242 -992
rect 8038 -1079 31242 -1044
rect 30219 -1083 31242 -1079
<< via1 >>
rect -15293 23151 -14217 23971
rect 5874 23207 6886 23963
rect 8103 23885 8987 24833
rect 30299 23901 31375 24721
rect 51466 23957 52478 24713
rect -13012 21376 -12000 22132
rect -4266 21362 -4261 22182
rect -4261 21362 -3579 22182
rect -3579 21362 -3574 22182
rect 3696 21378 4772 22198
rect 10363 22054 11247 23002
rect 32580 22126 33592 22882
rect 41326 22112 41331 22932
rect 41331 22112 42013 22932
rect 42013 22112 42018 22932
rect 49288 22128 50364 22948
rect 41523 19215 41767 19216
rect 41523 19037 41767 19215
rect 43599 19199 43715 19204
rect 43599 19093 43604 19199
rect 43604 19093 43710 19199
rect 43710 19093 43715 19199
rect 43599 19088 43715 19093
rect 41523 19036 41767 19037
rect -4069 18465 -3825 18466
rect -4069 18287 -3825 18465
rect -1993 18449 -1877 18454
rect -1993 18343 -1988 18449
rect -1988 18343 -1882 18449
rect -1882 18343 -1877 18449
rect -1993 18338 -1877 18343
rect -4069 18286 -3825 18287
rect -6244 17541 -6192 17550
rect -6244 17507 -6239 17541
rect -6239 17507 -6205 17541
rect -6205 17507 -6192 17541
rect -6244 17498 -6192 17507
rect -6180 17541 -6128 17550
rect -6180 17507 -6167 17541
rect -6167 17507 -6133 17541
rect -6133 17507 -6128 17541
rect -6180 17498 -6128 17507
rect -6207 17137 -6155 17175
rect -6207 17123 -6190 17137
rect -6190 17123 -6156 17137
rect -6156 17123 -6155 17137
rect -5866 16251 -5686 16367
rect -6369 16053 -6317 16105
rect -6305 16053 -6253 16105
rect -2682 18023 -2630 18075
rect -2682 17959 -2630 18011
rect -2682 17895 -2630 17947
rect -2934 16286 -2882 16338
rect -2934 16222 -2882 16274
rect -2934 16158 -2882 16210
rect -2173 18046 -2121 18075
rect -2173 18023 -2172 18046
rect -2172 18023 -2121 18046
rect -2173 17974 -2121 18011
rect -2173 17959 -2172 17974
rect -2172 17959 -2121 17974
rect -2173 17940 -2172 17947
rect -2172 17940 -2121 17947
rect -2173 17902 -2121 17940
rect -2173 17895 -2172 17902
rect -2172 17895 -2121 17902
rect -2434 16318 -2382 16334
rect -2434 16284 -2430 16318
rect -2430 16284 -2382 16318
rect -2434 16282 -2382 16284
rect -2434 16246 -2382 16270
rect -2434 16218 -2430 16246
rect -2430 16218 -2382 16246
rect -2434 16174 -2382 16206
rect -2434 16154 -2430 16174
rect -2430 16154 -2382 16174
rect -1658 18046 -1606 18071
rect -1658 18019 -1656 18046
rect -1656 18019 -1606 18046
rect -1658 17974 -1606 18007
rect -1658 17955 -1656 17974
rect -1656 17955 -1606 17974
rect -1658 17940 -1656 17943
rect -1656 17940 -1606 17943
rect -1658 17902 -1606 17940
rect -1658 17891 -1656 17902
rect -1656 17891 -1606 17902
rect -1920 16318 -1868 16340
rect -1920 16288 -1914 16318
rect -1914 16288 -1868 16318
rect -1920 16246 -1868 16276
rect -1920 16224 -1914 16246
rect -1914 16224 -1868 16246
rect -1920 16174 -1868 16212
rect -1920 16160 -1914 16174
rect -1914 16160 -1868 16174
rect -1139 18011 -1087 18063
rect -1139 17947 -1087 17999
rect -1139 17883 -1087 17935
rect -1404 16318 -1352 16341
rect -1404 16289 -1398 16318
rect -1398 16289 -1352 16318
rect -1404 16246 -1352 16277
rect -1404 16225 -1398 16246
rect -1398 16225 -1352 16246
rect -1404 16212 -1398 16213
rect -1398 16212 -1352 16213
rect -1404 16174 -1352 16212
rect -1404 16161 -1398 16174
rect -1398 16161 -1352 16174
rect -628 18046 -576 18067
rect -628 18015 -624 18046
rect -624 18015 -576 18046
rect -628 17974 -576 18003
rect -628 17951 -624 17974
rect -624 17951 -576 17974
rect -628 17902 -576 17939
rect -628 17887 -624 17902
rect -624 17887 -576 17902
rect -882 16292 -830 16344
rect -882 16228 -830 16280
rect -882 16164 -830 16216
rect 24684 18648 24736 18655
rect 24684 18614 24692 18648
rect 24692 18614 24726 18648
rect 24726 18614 24736 18648
rect 24684 18603 24736 18614
rect 24684 18576 24736 18591
rect 24684 18542 24692 18576
rect 24692 18542 24726 18576
rect 24726 18542 24736 18576
rect 24684 18539 24736 18542
rect 24684 18504 24736 18527
rect 24684 18475 24692 18504
rect 24692 18475 24726 18504
rect 24726 18475 24736 18504
rect 24684 18432 24736 18463
rect 24684 18411 24692 18432
rect 24692 18411 24726 18432
rect 24726 18411 24736 18432
rect 24684 18398 24692 18399
rect 24692 18398 24726 18399
rect 24726 18398 24736 18399
rect 24684 18360 24736 18398
rect 24684 18347 24692 18360
rect 24692 18347 24726 18360
rect 24726 18347 24736 18360
rect -376 16318 -324 16338
rect -376 16286 -366 16318
rect -366 16286 -324 16318
rect -376 16246 -324 16274
rect -376 16222 -366 16246
rect -366 16222 -324 16246
rect -376 16174 -324 16210
rect -376 16158 -366 16174
rect -366 16158 -324 16174
rect 23 16161 203 16341
rect -4214 15020 -4098 15200
rect -5437 14935 -5385 14944
rect -5437 14901 -5436 14935
rect -5436 14901 -5402 14935
rect -5402 14901 -5385 14935
rect -5437 14892 -5385 14901
rect -5373 14935 -5321 14944
rect -5373 14901 -5364 14935
rect -5364 14901 -5330 14935
rect -5330 14901 -5321 14935
rect -5373 14892 -5321 14901
rect -5309 14935 -5257 14944
rect -5309 14901 -5292 14935
rect -5292 14901 -5258 14935
rect -5258 14901 -5257 14935
rect -5309 14892 -5257 14901
rect 10333 15018 10358 17054
rect 10358 15018 11256 17054
rect 11256 15018 11281 17054
rect 26798 18648 26850 18659
rect 26798 18614 26808 18648
rect 26808 18614 26842 18648
rect 26842 18614 26850 18648
rect 26798 18607 26850 18614
rect 26798 18576 26850 18595
rect 26798 18543 26808 18576
rect 26808 18543 26842 18576
rect 26842 18543 26850 18576
rect 26798 18504 26850 18531
rect 26798 18479 26808 18504
rect 26808 18479 26842 18504
rect 26842 18479 26850 18504
rect 26798 18432 26850 18467
rect 26798 18415 26808 18432
rect 26808 18415 26842 18432
rect 26842 18415 26850 18432
rect 26798 18398 26808 18403
rect 26808 18398 26842 18403
rect 26842 18398 26850 18403
rect 26798 18360 26850 18398
rect 26798 18351 26808 18360
rect 26808 18351 26842 18360
rect 26842 18351 26850 18360
rect 25741 17534 25750 17557
rect 25750 17534 25784 17557
rect 25784 17534 25793 17557
rect 25741 17505 25793 17534
rect 25741 17462 25750 17493
rect 25750 17462 25784 17493
rect 25784 17462 25793 17493
rect 25741 17441 25793 17462
rect 25741 17424 25793 17429
rect 25741 17390 25750 17424
rect 25750 17390 25784 17424
rect 25784 17390 25793 17424
rect 25741 17377 25793 17390
rect 25741 17352 25793 17365
rect 25741 17318 25750 17352
rect 25750 17318 25784 17352
rect 25784 17318 25793 17352
rect 25741 17313 25793 17318
rect 25741 17280 25793 17301
rect 25741 17249 25750 17280
rect 25750 17249 25784 17280
rect 25784 17249 25793 17280
rect 39348 18291 39400 18300
rect 39348 18257 39353 18291
rect 39353 18257 39387 18291
rect 39387 18257 39400 18291
rect 39348 18248 39400 18257
rect 39412 18291 39464 18300
rect 39412 18257 39425 18291
rect 39425 18257 39459 18291
rect 39459 18257 39464 18291
rect 39412 18248 39464 18257
rect 39385 17887 39437 17925
rect 39385 17873 39402 17887
rect 39402 17873 39436 17887
rect 39436 17873 39437 17887
rect 27855 17534 27866 17555
rect 27866 17534 27900 17555
rect 27900 17534 27907 17555
rect 27855 17503 27907 17534
rect 27855 17462 27866 17491
rect 27866 17462 27900 17491
rect 27900 17462 27907 17491
rect 27855 17439 27907 17462
rect 27855 17424 27907 17427
rect 27855 17390 27866 17424
rect 27866 17390 27900 17424
rect 27900 17390 27907 17424
rect 27855 17375 27907 17390
rect 27855 17352 27907 17363
rect 27855 17318 27866 17352
rect 27866 17318 27900 17352
rect 27900 17318 27907 17352
rect 27855 17311 27907 17318
rect 27855 17280 27907 17299
rect 27855 17247 27866 17280
rect 27866 17247 27900 17280
rect 27900 17247 27907 17280
rect 39726 17001 39906 17117
rect 22553 15745 22925 16117
rect 27939 16248 28055 16812
rect 39223 16803 39275 16855
rect 39287 16803 39339 16855
rect 42910 18773 42962 18825
rect 42910 18709 42962 18761
rect 42910 18645 42962 18697
rect 42658 17036 42710 17088
rect 42658 16972 42710 17024
rect 42658 16908 42710 16960
rect 43419 18796 43471 18825
rect 43419 18773 43420 18796
rect 43420 18773 43471 18796
rect 43419 18724 43471 18761
rect 43419 18709 43420 18724
rect 43420 18709 43471 18724
rect 43419 18690 43420 18697
rect 43420 18690 43471 18697
rect 43419 18652 43471 18690
rect 43419 18645 43420 18652
rect 43420 18645 43471 18652
rect 43158 17068 43210 17084
rect 43158 17034 43162 17068
rect 43162 17034 43210 17068
rect 43158 17032 43210 17034
rect 43158 16996 43210 17020
rect 43158 16968 43162 16996
rect 43162 16968 43210 16996
rect 43158 16924 43210 16956
rect 43158 16904 43162 16924
rect 43162 16904 43210 16924
rect 43934 18796 43986 18821
rect 43934 18769 43936 18796
rect 43936 18769 43986 18796
rect 43934 18724 43986 18757
rect 43934 18705 43936 18724
rect 43936 18705 43986 18724
rect 43934 18690 43936 18693
rect 43936 18690 43986 18693
rect 43934 18652 43986 18690
rect 43934 18641 43936 18652
rect 43936 18641 43986 18652
rect 43672 17068 43724 17090
rect 43672 17038 43678 17068
rect 43678 17038 43724 17068
rect 43672 16996 43724 17026
rect 43672 16974 43678 16996
rect 43678 16974 43724 16996
rect 43672 16924 43724 16962
rect 43672 16910 43678 16924
rect 43678 16910 43724 16924
rect 44453 18761 44505 18813
rect 44453 18697 44505 18749
rect 44453 18633 44505 18685
rect 44188 17068 44240 17091
rect 44188 17039 44194 17068
rect 44194 17039 44240 17068
rect 44188 16996 44240 17027
rect 44188 16975 44194 16996
rect 44194 16975 44240 16996
rect 44188 16962 44194 16963
rect 44194 16962 44240 16963
rect 44188 16924 44240 16962
rect 44188 16911 44194 16924
rect 44194 16911 44240 16924
rect 44964 18796 45016 18817
rect 44964 18765 44968 18796
rect 44968 18765 45016 18796
rect 44964 18724 45016 18753
rect 44964 18701 44968 18724
rect 44968 18701 45016 18724
rect 44964 18652 45016 18689
rect 44964 18637 44968 18652
rect 44968 18637 45016 18652
rect 44710 17042 44762 17094
rect 44710 16978 44762 17030
rect 44710 16914 44762 16966
rect 45216 17068 45268 17088
rect 45216 17036 45226 17068
rect 45226 17036 45268 17068
rect 45216 16996 45268 17024
rect 45216 16972 45226 16996
rect 45226 16972 45268 16996
rect 45216 16924 45268 16960
rect 45216 16908 45226 16924
rect 45226 16908 45268 16924
rect 45602 16881 46486 18213
rect -6947 14754 -6943 14768
rect -6943 14754 -6909 14768
rect -6909 14754 -6895 14768
rect -6947 14716 -6895 14754
rect -6947 14682 -6943 14704
rect -6943 14682 -6909 14704
rect -6909 14682 -6895 14704
rect -6947 14652 -6895 14682
rect -6947 14610 -6943 14640
rect -6943 14610 -6909 14640
rect -6909 14610 -6895 14640
rect -6947 14588 -6895 14610
rect -7453 13060 -7401 13065
rect -7453 13026 -7425 13060
rect -7425 13026 -7401 13060
rect -7453 13013 -7401 13026
rect -7453 12988 -7401 13001
rect -7453 12954 -7425 12988
rect -7425 12954 -7401 12988
rect -7453 12949 -7401 12954
rect -7453 12916 -7401 12937
rect -7453 12885 -7425 12916
rect -7425 12885 -7401 12916
rect -5936 14754 -5911 14755
rect -5911 14754 -5884 14755
rect -5936 14716 -5884 14754
rect -5936 14703 -5911 14716
rect -5911 14703 -5884 14716
rect -5936 14682 -5911 14691
rect -5911 14682 -5884 14691
rect -5936 14644 -5884 14682
rect -5936 14639 -5911 14644
rect -5911 14639 -5884 14644
rect -5936 14610 -5911 14627
rect -5911 14610 -5884 14627
rect -5936 14575 -5884 14610
rect -6434 13060 -6382 13076
rect -6434 13026 -6427 13060
rect -6427 13026 -6393 13060
rect -6393 13026 -6382 13060
rect -6434 13024 -6382 13026
rect -6434 12988 -6382 13012
rect -6434 12960 -6427 12988
rect -6427 12960 -6393 12988
rect -6393 12960 -6382 12988
rect -6434 12916 -6382 12948
rect -6434 12896 -6427 12916
rect -6427 12896 -6393 12916
rect -6393 12896 -6382 12916
rect -4899 14754 -4879 14755
rect -4879 14754 -4847 14755
rect -4899 14716 -4847 14754
rect -4899 14703 -4879 14716
rect -4879 14703 -4847 14716
rect -4899 14682 -4879 14691
rect -4879 14682 -4847 14691
rect -4899 14644 -4847 14682
rect -4899 14639 -4879 14644
rect -4879 14639 -4847 14644
rect -4899 14610 -4879 14627
rect -4879 14610 -4847 14627
rect -4899 14575 -4847 14610
rect -5404 13060 -5352 13086
rect -5404 13034 -5395 13060
rect -5395 13034 -5361 13060
rect -5361 13034 -5352 13060
rect -5404 12988 -5352 13022
rect -5404 12970 -5395 12988
rect -5395 12970 -5361 12988
rect -5361 12970 -5352 12988
rect -5404 12954 -5395 12958
rect -5395 12954 -5361 12958
rect -5361 12954 -5352 12958
rect -5404 12916 -5352 12954
rect -5404 12906 -5395 12916
rect -5395 12906 -5361 12916
rect -5361 12906 -5352 12916
rect 13982 14508 14162 14509
rect 13982 14474 14052 14508
rect 14052 14474 14086 14508
rect 14086 14474 14162 14508
rect 13982 14436 14162 14474
rect 13982 14402 14052 14436
rect 14052 14402 14086 14436
rect 14086 14402 14162 14436
rect 13982 14364 14162 14402
rect 13982 14330 14052 14364
rect 14052 14330 14086 14364
rect 14086 14330 14162 14364
rect 13982 14292 14162 14330
rect 13982 14258 14052 14292
rect 14052 14258 14086 14292
rect 14086 14258 14162 14292
rect 13982 14220 14162 14258
rect 13982 14201 14052 14220
rect 14052 14201 14086 14220
rect 14086 14201 14162 14220
rect -6845 12758 -6793 12767
rect -6845 12724 -6840 12758
rect -6840 12724 -6806 12758
rect -6806 12724 -6793 12758
rect -6845 12715 -6793 12724
rect -6781 12758 -6729 12767
rect -6781 12724 -6768 12758
rect -6768 12724 -6734 12758
rect -6734 12724 -6729 12758
rect -6781 12715 -6729 12724
rect -5315 12570 -4815 12626
rect -5315 12536 -5262 12570
rect -5262 12536 -5228 12570
rect -5228 12536 -4815 12570
rect -5315 12498 -4815 12536
rect -5315 12464 -5262 12498
rect -5262 12464 -5228 12498
rect -5228 12464 -4815 12498
rect -5315 12446 -4815 12464
rect -3918 12820 -3862 12821
rect -3862 12820 -3828 12821
rect -3828 12820 -3802 12821
rect -3918 12782 -3802 12820
rect -3918 12748 -3862 12782
rect -3862 12748 -3828 12782
rect -3828 12748 -3802 12782
rect -3918 12710 -3802 12748
rect -3918 12676 -3862 12710
rect -3862 12676 -3828 12710
rect -3828 12676 -3802 12710
rect -3918 12638 -3802 12676
rect -3918 12604 -3862 12638
rect -3862 12604 -3828 12638
rect -3828 12604 -3802 12638
rect -3918 12566 -3802 12604
rect -3918 12532 -3862 12566
rect -3862 12532 -3828 12566
rect -3828 12532 -3802 12566
rect -3918 12494 -3802 12532
rect -3918 12460 -3862 12494
rect -3862 12460 -3828 12494
rect -3828 12460 -3802 12494
rect -3918 12449 -3802 12460
rect 13014 12026 13028 12052
rect 13028 12026 13130 12052
rect 13014 11988 13130 12026
rect 13014 11954 13028 11988
rect 13028 11954 13130 11988
rect 13014 11916 13130 11954
rect 13014 11882 13028 11916
rect 13028 11882 13130 11916
rect 13014 11844 13130 11882
rect 13014 11810 13028 11844
rect 13028 11810 13130 11844
rect 13014 11808 13130 11810
rect 14999 12026 15110 12052
rect 15110 12026 15115 12052
rect 14999 11988 15115 12026
rect 14999 11954 15110 11988
rect 15110 11954 15115 11988
rect 14999 11916 15115 11954
rect 14999 11882 15110 11916
rect 15110 11882 15115 11916
rect 14999 11844 15115 11882
rect 14999 11810 15110 11844
rect 15110 11810 15115 11844
rect 14999 11808 15115 11810
rect 15609 14201 15725 14509
rect 17104 12324 17108 12351
rect 17108 12324 17220 12351
rect 17104 12286 17220 12324
rect 17104 12252 17108 12286
rect 17108 12252 17220 12286
rect 17104 12214 17220 12252
rect 17104 12180 17108 12214
rect 17108 12180 17220 12214
rect 17104 12142 17220 12180
rect 17104 12108 17108 12142
rect 17108 12108 17220 12142
rect 17104 12070 17220 12108
rect 17104 12036 17108 12070
rect 17108 12036 17220 12070
rect 17104 11998 17220 12036
rect 17104 11979 17108 11998
rect 17108 11979 17220 11998
rect 29253 15208 29300 15215
rect 29300 15208 29334 15215
rect 29334 15208 29369 15215
rect 29253 15170 29369 15208
rect 29253 15136 29300 15170
rect 29300 15136 29334 15170
rect 29334 15136 29369 15170
rect 29253 15098 29369 15136
rect 29253 15064 29300 15098
rect 29300 15064 29334 15098
rect 29334 15064 29369 15098
rect 29253 15026 29369 15064
rect 29253 14992 29300 15026
rect 29300 14992 29334 15026
rect 29334 14992 29369 15026
rect 29253 14954 29369 14992
rect 29253 14920 29300 14954
rect 29300 14920 29334 14954
rect 29334 14920 29369 14954
rect 29253 14882 29369 14920
rect 29253 14848 29300 14882
rect 29300 14848 29334 14882
rect 29334 14848 29369 14882
rect 29253 14843 29369 14848
rect 19933 13499 20305 13871
rect 18498 12092 18538 12119
rect 18538 12092 18572 12119
rect 18572 12092 18614 12119
rect 18498 12054 18614 12092
rect 18498 12020 18538 12054
rect 18538 12020 18572 12054
rect 18572 12020 18614 12054
rect 18498 11982 18614 12020
rect 18498 11948 18538 11982
rect 18538 11948 18572 11982
rect 18572 11948 18614 11982
rect 18498 11939 18614 11948
rect -8566 10755 -8557 10766
rect -8557 10755 -8523 10766
rect -8523 10755 -8514 10766
rect -8566 10717 -8514 10755
rect -8566 10714 -8557 10717
rect -8557 10714 -8523 10717
rect -8523 10714 -8514 10717
rect -8566 10683 -8557 10702
rect -8557 10683 -8523 10702
rect -8523 10683 -8514 10702
rect -8566 10650 -8514 10683
rect -8051 10717 -7999 10733
rect -8051 10683 -8041 10717
rect -8041 10683 -8007 10717
rect -8007 10683 -7999 10717
rect -8051 10681 -7999 10683
rect -7534 10717 -7482 10732
rect -7534 10683 -7525 10717
rect -7525 10683 -7491 10717
rect -7491 10683 -7482 10717
rect -7534 10680 -7482 10683
rect -7018 10717 -6966 10733
rect -7018 10683 -7009 10717
rect -7009 10683 -6975 10717
rect -6975 10683 -6966 10717
rect -7018 10681 -6966 10683
rect -6502 10717 -6450 10731
rect -6502 10683 -6493 10717
rect -6493 10683 -6459 10717
rect -6459 10683 -6450 10717
rect -6502 10679 -6450 10683
rect -5986 10717 -5934 10732
rect -5986 10683 -5977 10717
rect -5977 10683 -5943 10717
rect -5943 10683 -5934 10717
rect -5986 10680 -5934 10683
rect -5470 10717 -5418 10731
rect -5470 10683 -5461 10717
rect -5461 10683 -5427 10717
rect -5427 10683 -5418 10717
rect -5470 10679 -5418 10683
rect -4954 10717 -4902 10732
rect -4954 10683 -4945 10717
rect -4945 10683 -4911 10717
rect -4911 10683 -4902 10717
rect -4954 10680 -4902 10683
rect -4438 10717 -4386 10732
rect -4438 10683 -4429 10717
rect -4429 10683 -4395 10717
rect -4395 10683 -4386 10717
rect -4438 10680 -4386 10683
rect -3922 10717 -3870 10732
rect -3922 10683 -3913 10717
rect -3913 10683 -3879 10717
rect -3879 10683 -3870 10717
rect -3922 10680 -3870 10683
rect 13276 10850 13584 10863
rect 13276 10816 13286 10850
rect 13286 10816 13352 10850
rect 13352 10816 13386 10850
rect 13386 10816 13452 10850
rect 13452 10816 13486 10850
rect 13486 10816 13552 10850
rect 13552 10816 13584 10850
rect 13276 10750 13584 10816
rect 13276 10716 13286 10750
rect 13286 10716 13352 10750
rect 13352 10716 13386 10750
rect 13386 10716 13452 10750
rect 13452 10716 13486 10750
rect 13486 10716 13552 10750
rect 13552 10716 13584 10750
rect 13276 10650 13584 10716
rect 13276 10616 13286 10650
rect 13286 10616 13352 10650
rect 13352 10616 13386 10650
rect 13386 10616 13452 10650
rect 13452 10616 13486 10650
rect 13486 10616 13552 10650
rect 13552 10616 13584 10650
rect 13276 10555 13584 10616
rect -9976 9928 -9412 10492
rect -8824 10467 -8815 10486
rect -8815 10467 -8781 10486
rect -8781 10467 -8772 10486
rect -8824 10434 -8772 10467
rect -8824 10395 -8815 10422
rect -8815 10395 -8781 10422
rect -8781 10395 -8772 10422
rect -8824 10370 -8772 10395
rect -8308 10467 -8299 10488
rect -8299 10467 -8265 10488
rect -8265 10467 -8256 10488
rect -8308 10436 -8256 10467
rect -8308 10395 -8299 10424
rect -8299 10395 -8265 10424
rect -8265 10395 -8256 10424
rect -8308 10372 -8256 10395
rect -7792 10467 -7783 10488
rect -7783 10467 -7749 10488
rect -7749 10467 -7740 10488
rect -7792 10436 -7740 10467
rect -7792 10395 -7783 10424
rect -7783 10395 -7749 10424
rect -7749 10395 -7740 10424
rect -7792 10372 -7740 10395
rect -7276 10467 -7267 10487
rect -7267 10467 -7233 10487
rect -7233 10467 -7224 10487
rect -7276 10435 -7224 10467
rect -7276 10395 -7267 10423
rect -7267 10395 -7233 10423
rect -7233 10395 -7224 10423
rect -7276 10371 -7224 10395
rect -6760 10467 -6751 10488
rect -6751 10467 -6717 10488
rect -6717 10467 -6708 10488
rect -6760 10436 -6708 10467
rect -6760 10395 -6751 10424
rect -6751 10395 -6717 10424
rect -6717 10395 -6708 10424
rect -6760 10372 -6708 10395
rect -6243 10467 -6235 10489
rect -6235 10467 -6201 10489
rect -6201 10467 -6191 10489
rect -6243 10437 -6191 10467
rect -6243 10395 -6235 10425
rect -6235 10395 -6201 10425
rect -6201 10395 -6191 10425
rect -6243 10373 -6191 10395
rect -5728 10467 -5719 10486
rect -5719 10467 -5685 10486
rect -5685 10467 -5676 10486
rect -5728 10434 -5676 10467
rect -5728 10395 -5719 10422
rect -5719 10395 -5685 10422
rect -5685 10395 -5676 10422
rect -5728 10370 -5676 10395
rect -5213 10467 -5203 10487
rect -5203 10467 -5169 10487
rect -5169 10467 -5161 10487
rect -5213 10435 -5161 10467
rect -5213 10395 -5203 10423
rect -5203 10395 -5169 10423
rect -5169 10395 -5161 10423
rect -5213 10371 -5161 10395
rect -4696 10467 -4687 10488
rect -4687 10467 -4653 10488
rect -4653 10467 -4644 10488
rect -4696 10436 -4644 10467
rect -4696 10395 -4687 10424
rect -4687 10395 -4653 10424
rect -4653 10395 -4644 10424
rect -4696 10372 -4644 10395
rect -4180 10467 -4171 10487
rect -4171 10467 -4137 10487
rect -4137 10467 -4128 10487
rect -4180 10435 -4128 10467
rect -4180 10395 -4171 10423
rect -4171 10395 -4137 10423
rect -4137 10395 -4128 10423
rect -4180 10371 -4128 10395
rect -3664 10467 -3655 10487
rect -3655 10467 -3621 10487
rect -3621 10467 -3612 10487
rect -3664 10435 -3612 10467
rect -3664 10395 -3655 10423
rect -3655 10395 -3621 10423
rect -3621 10395 -3612 10423
rect -3664 10371 -3612 10395
rect -7065 9462 -7056 9478
rect -7056 9462 -7022 9478
rect -7022 9462 -7013 9478
rect -7065 9426 -7013 9462
rect -7065 9390 -7056 9414
rect -7056 9390 -7022 9414
rect -7022 9390 -7013 9414
rect -7065 9362 -7013 9390
rect -7322 9102 -7314 9128
rect -7314 9102 -7280 9128
rect -7280 9102 -7270 9128
rect -7322 9076 -7270 9102
rect -7322 9030 -7314 9064
rect -7314 9030 -7280 9064
rect -7280 9030 -7270 9064
rect -7322 9012 -7270 9030
rect -6549 9462 -6540 9475
rect -6540 9462 -6506 9475
rect -6506 9462 -6497 9475
rect -6549 9424 -6497 9462
rect -6549 9423 -6540 9424
rect -6540 9423 -6506 9424
rect -6506 9423 -6497 9424
rect -6549 9390 -6540 9411
rect -6540 9390 -6506 9411
rect -6506 9390 -6497 9411
rect -6549 9359 -6497 9390
rect -6805 9102 -6798 9127
rect -6798 9102 -6764 9127
rect -6764 9102 -6753 9127
rect -6805 9075 -6753 9102
rect -6805 9030 -6798 9063
rect -6798 9030 -6764 9063
rect -6764 9030 -6753 9063
rect -6805 9011 -6753 9030
rect -6033 9462 -6024 9477
rect -6024 9462 -5990 9477
rect -5990 9462 -5981 9477
rect -6033 9425 -5981 9462
rect -6033 9390 -6024 9413
rect -6024 9390 -5990 9413
rect -5990 9390 -5981 9413
rect -6033 9361 -5981 9390
rect -6292 9102 -6282 9129
rect -6282 9102 -6248 9129
rect -6248 9102 -6240 9129
rect -6292 9077 -6240 9102
rect -6292 9064 -6240 9065
rect -6292 9030 -6282 9064
rect -6282 9030 -6248 9064
rect -6248 9030 -6240 9064
rect -6292 9013 -6240 9030
rect -5516 9462 -5508 9475
rect -5508 9462 -5474 9475
rect -5474 9462 -5464 9475
rect -5516 9424 -5464 9462
rect -5516 9423 -5508 9424
rect -5508 9423 -5474 9424
rect -5474 9423 -5464 9424
rect -5516 9390 -5508 9411
rect -5508 9390 -5474 9411
rect -5474 9390 -5464 9411
rect -5516 9359 -5464 9390
rect -5774 9102 -5766 9128
rect -5766 9102 -5732 9128
rect -5732 9102 -5722 9128
rect -5774 9076 -5722 9102
rect -5774 9030 -5766 9064
rect -5766 9030 -5732 9064
rect -5732 9030 -5722 9064
rect -5774 9012 -5722 9030
rect -5002 9462 -4992 9476
rect -4992 9462 -4958 9476
rect -4958 9462 -4950 9476
rect -5002 9424 -4950 9462
rect -5002 9390 -4992 9412
rect -4992 9390 -4958 9412
rect -4958 9390 -4950 9412
rect -5002 9360 -4950 9390
rect -5257 9102 -5250 9128
rect -5250 9102 -5216 9128
rect -5216 9102 -5205 9128
rect -5257 9076 -5205 9102
rect -5257 9030 -5250 9064
rect -5250 9030 -5216 9064
rect -5216 9030 -5205 9064
rect -5257 9012 -5205 9030
rect 13262 9326 13286 9356
rect 13286 9326 13352 9356
rect 13352 9326 13386 9356
rect 13386 9326 13452 9356
rect 13452 9326 13486 9356
rect 13486 9326 13552 9356
rect 13552 9326 13570 9356
rect 13262 9260 13570 9326
rect 13262 9226 13286 9260
rect 13286 9226 13352 9260
rect 13352 9226 13386 9260
rect 13386 9226 13452 9260
rect 13452 9226 13486 9260
rect 13486 9226 13552 9260
rect 13552 9226 13570 9260
rect -4742 9102 -4734 9129
rect -4734 9102 -4700 9129
rect -4700 9102 -4690 9129
rect -4742 9077 -4690 9102
rect -4742 9064 -4690 9065
rect -4742 9030 -4734 9064
rect -4734 9030 -4700 9064
rect -4700 9030 -4690 9064
rect -4742 9013 -4690 9030
rect 13262 9160 13570 9226
rect 13262 9126 13286 9160
rect 13286 9126 13352 9160
rect 13352 9126 13386 9160
rect 13386 9126 13452 9160
rect 13452 9126 13486 9160
rect 13486 9126 13552 9160
rect 13552 9126 13570 9160
rect 13262 9060 13570 9126
rect 13262 9048 13286 9060
rect 13286 9048 13352 9060
rect 13352 9048 13386 9060
rect 13386 9048 13452 9060
rect 13452 9048 13486 9060
rect 13486 9048 13552 9060
rect 13552 9048 13570 9060
rect 16956 11339 17008 11391
rect 17626 11324 17678 11376
rect 15989 11170 16012 11182
rect 16012 11170 16046 11182
rect 16046 11170 16105 11182
rect 15989 11132 16105 11170
rect 15989 11098 16012 11132
rect 16012 11098 16046 11132
rect 16046 11098 16105 11132
rect 15989 11060 16105 11098
rect 15989 11026 16012 11060
rect 16012 11026 16046 11060
rect 16046 11026 16105 11060
rect 15989 10988 16105 11026
rect 15989 10954 16012 10988
rect 16012 10954 16046 10988
rect 16046 10954 16105 10988
rect 15989 10938 16105 10954
rect 14979 8650 14988 8676
rect 14988 8650 15095 8676
rect 14979 8612 15095 8650
rect 14979 8578 14988 8612
rect 14988 8578 15095 8612
rect 14979 8540 15095 8578
rect 14979 8506 14988 8540
rect 14988 8506 15095 8540
rect 14979 8468 15095 8506
rect 14979 8434 14988 8468
rect 14988 8434 15095 8468
rect 14979 8396 15095 8434
rect 14979 8362 14988 8396
rect 14988 8362 15095 8396
rect 14979 8324 15095 8362
rect 14979 8304 14988 8324
rect 14988 8304 15095 8324
rect 18498 11106 18614 11129
rect 18498 11072 18536 11106
rect 18536 11072 18570 11106
rect 18570 11072 18614 11106
rect 18498 11034 18614 11072
rect 18498 11000 18536 11034
rect 18536 11000 18570 11034
rect 18570 11000 18614 11034
rect 18498 10962 18614 11000
rect 18498 10949 18536 10962
rect 18536 10949 18570 10962
rect 18570 10949 18614 10962
rect 16959 8650 17070 8676
rect 17070 8650 17075 8676
rect 16959 8612 17075 8650
rect 16959 8578 17070 8612
rect 17070 8578 17075 8612
rect 16959 8540 17075 8578
rect 16959 8506 17070 8540
rect 17070 8506 17075 8540
rect 16959 8468 17075 8506
rect 16959 8434 17070 8468
rect 17070 8434 17075 8468
rect 16959 8396 17075 8434
rect 16959 8362 17070 8396
rect 17070 8362 17075 8396
rect 16959 8324 17075 8362
rect 16959 8304 17070 8324
rect 17070 8304 17075 8324
rect 16922 8166 16935 8187
rect 16935 8166 16973 8187
rect 16973 8166 17007 8187
rect 17007 8166 17038 8187
rect 16922 8007 17038 8166
rect -7980 5852 -7969 5886
rect -7969 5852 -7935 5886
rect -7935 5852 -7928 5886
rect -7980 5834 -7928 5852
rect -7980 5814 -7928 5822
rect -7980 5780 -7969 5814
rect -7969 5780 -7935 5814
rect -7935 5780 -7928 5814
rect -7980 5770 -7928 5780
rect -7980 5742 -7928 5758
rect -7980 5708 -7969 5742
rect -7969 5708 -7935 5742
rect -7935 5708 -7928 5742
rect -7980 5706 -7928 5708
rect -7273 6737 -7264 6765
rect -7264 6737 -7230 6765
rect -7230 6737 -7221 6765
rect -7273 6713 -7221 6737
rect -7273 6699 -7221 6701
rect -7273 6665 -7264 6699
rect -7264 6665 -7230 6699
rect -7230 6665 -7221 6699
rect -7273 6649 -7221 6665
rect -7532 5873 -7522 5888
rect -7522 5873 -7488 5888
rect -7488 5873 -7480 5888
rect -7532 5836 -7480 5873
rect -7532 5801 -7522 5824
rect -7522 5801 -7488 5824
rect -7488 5801 -7480 5824
rect -7532 5772 -7480 5801
rect -7532 5729 -7522 5760
rect -7522 5729 -7488 5760
rect -7488 5729 -7480 5760
rect -7532 5708 -7480 5729
rect -6757 6339 -6705 6362
rect -6757 6310 -6748 6339
rect -6748 6310 -6714 6339
rect -6714 6310 -6705 6339
rect -6757 6267 -6705 6298
rect -6757 6246 -6748 6267
rect -6748 6246 -6714 6267
rect -6714 6246 -6705 6267
rect -6757 6233 -6748 6234
rect -6748 6233 -6714 6234
rect -6714 6233 -6705 6234
rect -6757 6195 -6705 6233
rect -6757 6182 -6748 6195
rect -6748 6182 -6714 6195
rect -6714 6182 -6705 6195
rect -7015 5873 -7006 5887
rect -7006 5873 -6972 5887
rect -6972 5873 -6963 5887
rect -7015 5835 -6963 5873
rect -7015 5801 -7006 5823
rect -7006 5801 -6972 5823
rect -6972 5801 -6963 5823
rect -7015 5771 -6963 5801
rect -7015 5729 -7006 5759
rect -7006 5729 -6972 5759
rect -6972 5729 -6963 5759
rect -7015 5707 -6963 5729
rect -6241 6339 -6189 6360
rect -6241 6308 -6232 6339
rect -6232 6308 -6198 6339
rect -6198 6308 -6189 6339
rect -6241 6267 -6189 6296
rect -6241 6244 -6232 6267
rect -6232 6244 -6198 6267
rect -6198 6244 -6189 6267
rect -6241 6195 -6189 6232
rect -6241 6180 -6232 6195
rect -6232 6180 -6198 6195
rect -6198 6180 -6189 6195
rect -6499 5873 -6490 5886
rect -6490 5873 -6456 5886
rect -6456 5873 -6447 5886
rect -6499 5835 -6447 5873
rect -6499 5834 -6490 5835
rect -6490 5834 -6456 5835
rect -6456 5834 -6447 5835
rect -6499 5801 -6490 5822
rect -6490 5801 -6456 5822
rect -6456 5801 -6447 5822
rect -6499 5770 -6447 5801
rect -6499 5729 -6490 5758
rect -6490 5729 -6456 5758
rect -6456 5729 -6447 5758
rect -6499 5706 -6447 5729
rect -5726 6305 -5716 6328
rect -5716 6305 -5682 6328
rect -5682 6305 -5674 6328
rect -5726 6276 -5674 6305
rect -5726 6233 -5716 6264
rect -5716 6233 -5682 6264
rect -5682 6233 -5674 6264
rect -5726 6212 -5674 6233
rect -5985 5873 -5974 5887
rect -5974 5873 -5940 5887
rect -5940 5873 -5933 5887
rect -5985 5835 -5933 5873
rect -5985 5801 -5974 5823
rect -5974 5801 -5940 5823
rect -5940 5801 -5933 5823
rect -5985 5771 -5933 5801
rect -5985 5729 -5974 5759
rect -5974 5729 -5940 5759
rect -5940 5729 -5933 5759
rect -5985 5707 -5933 5729
rect -5209 6339 -5157 6361
rect -5209 6309 -5200 6339
rect -5200 6309 -5166 6339
rect -5166 6309 -5157 6339
rect -5209 6267 -5157 6297
rect -5209 6245 -5200 6267
rect -5200 6245 -5166 6267
rect -5166 6245 -5157 6267
rect -5209 6195 -5157 6233
rect -5209 6181 -5200 6195
rect -5200 6181 -5166 6195
rect -5166 6181 -5157 6195
rect -4175 6737 -4168 6764
rect -4168 6737 -4134 6764
rect -4134 6737 -4123 6764
rect -4175 6712 -4123 6737
rect -4175 6699 -4123 6700
rect -4175 6665 -4168 6699
rect -4168 6665 -4134 6699
rect -4134 6665 -4123 6699
rect -4175 6648 -4123 6665
rect -5467 5873 -5458 5886
rect -5458 5873 -5424 5886
rect -5424 5873 -5415 5886
rect -5467 5835 -5415 5873
rect -5467 5834 -5458 5835
rect -5458 5834 -5424 5835
rect -5424 5834 -5415 5835
rect -5467 5801 -5458 5822
rect -5458 5801 -5424 5822
rect -5424 5801 -5415 5822
rect -5467 5770 -5415 5801
rect -5467 5729 -5458 5758
rect -5458 5729 -5424 5758
rect -5424 5729 -5415 5758
rect -5467 5706 -5415 5729
rect -4694 6339 -4642 6359
rect -4694 6307 -4684 6339
rect -4684 6307 -4650 6339
rect -4650 6307 -4642 6339
rect -4694 6267 -4642 6295
rect -4694 6243 -4684 6267
rect -4684 6243 -4650 6267
rect -4650 6243 -4642 6267
rect -4694 6195 -4642 6231
rect -4694 6179 -4684 6195
rect -4684 6179 -4650 6195
rect -4650 6179 -4642 6195
rect -4952 5873 -4942 5887
rect -4942 5873 -4908 5887
rect -4908 5873 -4900 5887
rect -4952 5835 -4900 5873
rect -4952 5801 -4942 5823
rect -4942 5801 -4908 5823
rect -4908 5801 -4900 5823
rect -4952 5771 -4900 5801
rect -4952 5729 -4942 5759
rect -4942 5729 -4908 5759
rect -4908 5729 -4900 5759
rect -4952 5707 -4900 5729
rect -4435 5873 -4426 5887
rect -4426 5873 -4392 5887
rect -4392 5873 -4383 5887
rect -4435 5835 -4383 5873
rect -4435 5801 -4426 5823
rect -4426 5801 -4392 5823
rect -4392 5801 -4383 5823
rect -4435 5771 -4383 5801
rect -4435 5729 -4426 5759
rect -4426 5729 -4392 5759
rect -4392 5729 -4383 5759
rect -4435 5707 -4383 5729
rect 16872 7633 17052 7877
rect 17468 8624 17478 8638
rect 17478 8624 17512 8638
rect 17512 8624 17584 8638
rect 17468 8586 17584 8624
rect 17468 8552 17478 8586
rect 17478 8552 17512 8586
rect 17512 8552 17584 8586
rect 17468 8514 17584 8552
rect 17468 8480 17478 8514
rect 17478 8480 17512 8514
rect 17512 8480 17584 8514
rect 17468 8442 17584 8480
rect 17468 8408 17478 8442
rect 17478 8408 17512 8442
rect 17512 8408 17584 8442
rect 17468 8370 17584 8408
rect 17468 8336 17478 8370
rect 17478 8336 17512 8370
rect 17512 8336 17584 8370
rect 17468 8330 17584 8336
rect 40155 15685 40207 15694
rect 40155 15651 40156 15685
rect 40156 15651 40190 15685
rect 40190 15651 40207 15685
rect 40155 15642 40207 15651
rect 40219 15685 40271 15694
rect 40219 15651 40228 15685
rect 40228 15651 40262 15685
rect 40262 15651 40271 15685
rect 40219 15642 40271 15651
rect 40283 15685 40335 15694
rect 40283 15651 40300 15685
rect 40300 15651 40334 15685
rect 40334 15651 40335 15685
rect 40283 15642 40335 15651
rect 38645 15504 38649 15518
rect 38649 15504 38683 15518
rect 38683 15504 38697 15518
rect 38645 15466 38697 15504
rect 38645 15432 38649 15454
rect 38649 15432 38683 15454
rect 38683 15432 38697 15454
rect 38645 15402 38697 15432
rect 38645 15360 38649 15390
rect 38649 15360 38683 15390
rect 38683 15360 38697 15390
rect 38645 15338 38697 15360
rect 38139 13810 38191 13815
rect 38139 13776 38167 13810
rect 38167 13776 38191 13810
rect 38139 13763 38191 13776
rect 38139 13738 38191 13751
rect 38139 13704 38167 13738
rect 38167 13704 38191 13738
rect 38139 13699 38191 13704
rect 38139 13666 38191 13687
rect 38139 13635 38167 13666
rect 38167 13635 38191 13666
rect 39656 15504 39681 15505
rect 39681 15504 39708 15505
rect 39656 15466 39708 15504
rect 39656 15453 39681 15466
rect 39681 15453 39708 15466
rect 39656 15432 39681 15441
rect 39681 15432 39708 15441
rect 39656 15394 39708 15432
rect 39656 15389 39681 15394
rect 39681 15389 39708 15394
rect 39656 15360 39681 15377
rect 39681 15360 39708 15377
rect 39656 15325 39708 15360
rect 39158 13810 39210 13826
rect 39158 13776 39165 13810
rect 39165 13776 39199 13810
rect 39199 13776 39210 13810
rect 39158 13774 39210 13776
rect 39158 13738 39210 13762
rect 39158 13710 39165 13738
rect 39165 13710 39199 13738
rect 39199 13710 39210 13738
rect 39158 13666 39210 13698
rect 39158 13646 39165 13666
rect 39165 13646 39199 13666
rect 39199 13646 39210 13666
rect 40693 15504 40713 15505
rect 40713 15504 40745 15505
rect 40693 15466 40745 15504
rect 40693 15453 40713 15466
rect 40713 15453 40745 15466
rect 40693 15432 40713 15441
rect 40713 15432 40745 15441
rect 40693 15394 40745 15432
rect 40693 15389 40713 15394
rect 40713 15389 40745 15394
rect 40693 15360 40713 15377
rect 40713 15360 40745 15377
rect 40693 15325 40745 15360
rect 40188 13810 40240 13836
rect 40188 13784 40197 13810
rect 40197 13784 40231 13810
rect 40231 13784 40240 13810
rect 40188 13738 40240 13772
rect 40188 13720 40197 13738
rect 40197 13720 40231 13738
rect 40231 13720 40240 13738
rect 40188 13704 40197 13708
rect 40197 13704 40231 13708
rect 40231 13704 40240 13708
rect 40188 13666 40240 13704
rect 40188 13656 40197 13666
rect 40197 13656 40231 13666
rect 40231 13656 40240 13666
rect 24826 13316 24856 13348
rect 24856 13316 24878 13348
rect 24826 13296 24878 13316
rect 26697 13290 26864 13298
rect 26864 13290 26877 13298
rect 26697 13252 26877 13290
rect 26697 13218 26864 13252
rect 26864 13218 26877 13252
rect 26697 13180 26877 13218
rect 26697 13146 26864 13180
rect 26864 13146 26877 13180
rect 26697 13108 26877 13146
rect 26697 13074 26864 13108
rect 26864 13074 26877 13108
rect 26697 13036 26877 13074
rect 26697 13002 26864 13036
rect 26864 13002 26877 13036
rect 26697 12964 26877 13002
rect 26697 12930 26864 12964
rect 26864 12930 26877 12964
rect 26697 12926 26877 12930
rect 37145 13175 37645 13547
rect 38747 13508 38799 13517
rect 38747 13474 38752 13508
rect 38752 13474 38786 13508
rect 38786 13474 38799 13508
rect 38747 13465 38799 13474
rect 38811 13508 38863 13517
rect 38811 13474 38824 13508
rect 38824 13474 38858 13508
rect 38858 13474 38863 13508
rect 38811 13465 38863 13474
rect 41674 13570 41730 13571
rect 41730 13570 41764 13571
rect 41764 13570 41790 13571
rect 41674 13532 41790 13570
rect 41674 13498 41730 13532
rect 41730 13498 41764 13532
rect 41764 13498 41790 13532
rect 41674 13460 41790 13498
rect 41674 13426 41730 13460
rect 41730 13426 41764 13460
rect 41764 13426 41790 13460
rect 41674 13388 41790 13426
rect 41674 13354 41730 13388
rect 41730 13354 41764 13388
rect 41764 13354 41790 13388
rect 41674 13316 41790 13354
rect 41674 13282 41730 13316
rect 41730 13282 41764 13316
rect 41764 13282 41790 13316
rect 41674 13244 41790 13282
rect 41674 13210 41730 13244
rect 41730 13210 41764 13244
rect 41764 13210 41790 13244
rect 41674 13199 41790 13210
rect 25666 12292 25718 12298
rect 25666 12258 25682 12292
rect 25682 12258 25718 12292
rect 25666 12246 25718 12258
rect 37026 11505 37035 11516
rect 37035 11505 37069 11516
rect 37069 11505 37078 11516
rect 37026 11467 37078 11505
rect 37026 11464 37035 11467
rect 37035 11464 37069 11467
rect 37069 11464 37078 11467
rect 37026 11433 37035 11452
rect 37035 11433 37069 11452
rect 37069 11433 37078 11452
rect 37026 11400 37078 11433
rect 37541 11467 37593 11483
rect 37541 11433 37551 11467
rect 37551 11433 37585 11467
rect 37585 11433 37593 11467
rect 37541 11431 37593 11433
rect 38058 11467 38110 11482
rect 38058 11433 38067 11467
rect 38067 11433 38101 11467
rect 38101 11433 38110 11467
rect 38058 11430 38110 11433
rect 38574 11467 38626 11483
rect 38574 11433 38583 11467
rect 38583 11433 38617 11467
rect 38617 11433 38626 11467
rect 38574 11431 38626 11433
rect 39090 11467 39142 11481
rect 39090 11433 39099 11467
rect 39099 11433 39133 11467
rect 39133 11433 39142 11467
rect 39090 11429 39142 11433
rect 39606 11467 39658 11482
rect 39606 11433 39615 11467
rect 39615 11433 39649 11467
rect 39649 11433 39658 11467
rect 39606 11430 39658 11433
rect 40122 11467 40174 11481
rect 40122 11433 40131 11467
rect 40131 11433 40165 11467
rect 40165 11433 40174 11467
rect 40122 11429 40174 11433
rect 40638 11467 40690 11482
rect 40638 11433 40647 11467
rect 40647 11433 40681 11467
rect 40681 11433 40690 11467
rect 40638 11430 40690 11433
rect 41154 11467 41206 11482
rect 41154 11433 41163 11467
rect 41163 11433 41197 11467
rect 41197 11433 41206 11467
rect 41154 11430 41206 11433
rect 41670 11467 41722 11482
rect 41670 11433 41679 11467
rect 41679 11433 41713 11467
rect 41713 11433 41722 11467
rect 41670 11430 41722 11433
rect 24826 11234 24878 11243
rect 24826 11200 24856 11234
rect 24856 11200 24878 11234
rect 24826 11191 24878 11200
rect 36768 11217 36777 11236
rect 36777 11217 36811 11236
rect 36811 11217 36820 11236
rect 36768 11184 36820 11217
rect 21137 9038 21253 9346
rect 22655 9251 23027 10391
rect 19478 8330 19594 8638
rect 17885 8140 17897 8166
rect 17897 8140 17935 8166
rect 17935 8140 17937 8166
rect 17949 8140 17969 8166
rect 17969 8140 18001 8166
rect 18013 8140 18041 8166
rect 18041 8140 18065 8166
rect 17885 8114 17937 8140
rect 17949 8114 18001 8140
rect 18013 8114 18065 8140
rect 18077 8140 18079 8166
rect 18079 8140 18113 8166
rect 18113 8140 18129 8166
rect 18077 8114 18129 8140
rect 36768 11145 36777 11172
rect 36777 11145 36811 11172
rect 36811 11145 36820 11172
rect 36768 11120 36820 11145
rect 37284 11217 37293 11238
rect 37293 11217 37327 11238
rect 37327 11217 37336 11238
rect 37284 11186 37336 11217
rect 37284 11145 37293 11174
rect 37293 11145 37327 11174
rect 37327 11145 37336 11174
rect 37284 11122 37336 11145
rect 37800 11217 37809 11238
rect 37809 11217 37843 11238
rect 37843 11217 37852 11238
rect 37800 11186 37852 11217
rect 37800 11145 37809 11174
rect 37809 11145 37843 11174
rect 37843 11145 37852 11174
rect 37800 11122 37852 11145
rect 38316 11217 38325 11237
rect 38325 11217 38359 11237
rect 38359 11217 38368 11237
rect 38316 11185 38368 11217
rect 38316 11145 38325 11173
rect 38325 11145 38359 11173
rect 38359 11145 38368 11173
rect 38316 11121 38368 11145
rect 38832 11217 38841 11238
rect 38841 11217 38875 11238
rect 38875 11217 38884 11238
rect 38832 11186 38884 11217
rect 38832 11145 38841 11174
rect 38841 11145 38875 11174
rect 38875 11145 38884 11174
rect 38832 11122 38884 11145
rect 39349 11217 39357 11239
rect 39357 11217 39391 11239
rect 39391 11217 39401 11239
rect 39349 11187 39401 11217
rect 39349 11145 39357 11175
rect 39357 11145 39391 11175
rect 39391 11145 39401 11175
rect 39349 11123 39401 11145
rect 39864 11217 39873 11236
rect 39873 11217 39907 11236
rect 39907 11217 39916 11236
rect 39864 11184 39916 11217
rect 39864 11145 39873 11172
rect 39873 11145 39907 11172
rect 39907 11145 39916 11172
rect 39864 11120 39916 11145
rect 40379 11217 40389 11237
rect 40389 11217 40423 11237
rect 40423 11217 40431 11237
rect 40379 11185 40431 11217
rect 40379 11145 40389 11173
rect 40389 11145 40423 11173
rect 40423 11145 40431 11173
rect 40379 11121 40431 11145
rect 40896 11217 40905 11238
rect 40905 11217 40939 11238
rect 40939 11217 40948 11238
rect 40896 11186 40948 11217
rect 40896 11145 40905 11174
rect 40905 11145 40939 11174
rect 40939 11145 40948 11174
rect 40896 11122 40948 11145
rect 41412 11217 41421 11237
rect 41421 11217 41455 11237
rect 41455 11217 41464 11237
rect 41412 11185 41464 11217
rect 41412 11145 41421 11173
rect 41421 11145 41455 11173
rect 41455 11145 41464 11173
rect 41412 11121 41464 11145
rect 41928 11217 41937 11237
rect 41937 11217 41971 11237
rect 41971 11217 41980 11237
rect 41928 11185 41980 11217
rect 41928 11145 41937 11173
rect 41937 11145 41971 11173
rect 41971 11145 41980 11173
rect 41928 11121 41980 11145
rect 25671 10176 25723 10198
rect 25671 10146 25682 10176
rect 25682 10146 25720 10176
rect 25720 10146 25723 10176
rect 24826 9118 24878 9138
rect 38527 10212 38536 10228
rect 38536 10212 38570 10228
rect 38570 10212 38579 10228
rect 38527 10176 38579 10212
rect 38527 10140 38536 10164
rect 38536 10140 38570 10164
rect 38570 10140 38579 10164
rect 38527 10112 38579 10140
rect 38270 9852 38278 9878
rect 38278 9852 38312 9878
rect 38312 9852 38322 9878
rect 38270 9826 38322 9852
rect 38270 9780 38278 9814
rect 38278 9780 38312 9814
rect 38312 9780 38322 9814
rect 38270 9762 38322 9780
rect 24826 9086 24856 9118
rect 24856 9086 24878 9118
rect 23664 7846 23697 7873
rect 23697 7846 23716 7873
rect 23728 7846 23731 7873
rect 23731 7846 23769 7873
rect 23769 7846 23780 7873
rect -3662 6771 -3610 6798
rect -3662 6746 -3652 6771
rect -3652 6746 -3618 6771
rect -3618 6746 -3610 6771
rect -3662 6699 -3610 6734
rect -3662 6682 -3652 6699
rect -3652 6682 -3618 6699
rect -3618 6682 -3610 6699
rect -3662 6665 -3652 6670
rect -3652 6665 -3618 6670
rect -3618 6665 -3610 6670
rect -3662 6627 -3610 6665
rect -3662 6618 -3652 6627
rect -3652 6618 -3618 6627
rect -3618 6618 -3610 6627
rect 17455 7145 17699 7180
rect 17455 7111 17468 7145
rect 17468 7111 17699 7145
rect -3919 5873 -3910 5887
rect -3910 5873 -3876 5887
rect -3876 5873 -3867 5887
rect -3919 5835 -3867 5873
rect -3919 5801 -3910 5823
rect -3910 5801 -3876 5823
rect -3876 5801 -3867 5823
rect -3919 5771 -3867 5801
rect -3919 5729 -3910 5759
rect -3910 5729 -3876 5759
rect -3876 5729 -3867 5759
rect -3919 5707 -3867 5729
rect 17455 7073 17699 7111
rect 17455 7039 17468 7073
rect 17468 7039 17699 7073
rect 17455 7001 17699 7039
rect 17455 7000 17468 7001
rect 17468 7000 17699 7001
rect 16436 6359 16616 6539
rect -3465 5851 -3456 5885
rect -3456 5851 -3422 5885
rect -3422 5851 -3413 5885
rect -3465 5833 -3413 5851
rect -3465 5813 -3413 5821
rect -3465 5779 -3456 5813
rect -3456 5779 -3422 5813
rect -3422 5779 -3413 5813
rect -3465 5769 -3413 5779
rect -3465 5741 -3413 5757
rect -3465 5707 -3456 5741
rect -3456 5707 -3422 5741
rect -3422 5707 -3413 5741
rect -3465 5705 -3413 5707
rect 23664 7821 23716 7846
rect 23728 7821 23780 7846
rect 25164 7846 25197 7863
rect 25197 7846 25216 7863
rect 25228 7846 25231 7863
rect 25231 7846 25269 7863
rect 25269 7846 25280 7863
rect 25164 7811 25216 7846
rect 25228 7811 25280 7846
rect 26222 7479 26338 8427
rect 39043 10212 39052 10225
rect 39052 10212 39086 10225
rect 39086 10212 39095 10225
rect 39043 10174 39095 10212
rect 39043 10173 39052 10174
rect 39052 10173 39086 10174
rect 39086 10173 39095 10174
rect 39043 10140 39052 10161
rect 39052 10140 39086 10161
rect 39086 10140 39095 10161
rect 39043 10109 39095 10140
rect 38787 9852 38794 9877
rect 38794 9852 38828 9877
rect 38828 9852 38839 9877
rect 38787 9825 38839 9852
rect 38787 9780 38794 9813
rect 38794 9780 38828 9813
rect 38828 9780 38839 9813
rect 38787 9761 38839 9780
rect 39559 10212 39568 10227
rect 39568 10212 39602 10227
rect 39602 10212 39611 10227
rect 39559 10175 39611 10212
rect 39559 10140 39568 10163
rect 39568 10140 39602 10163
rect 39602 10140 39611 10163
rect 39559 10111 39611 10140
rect 39300 9852 39310 9879
rect 39310 9852 39344 9879
rect 39344 9852 39352 9879
rect 39300 9827 39352 9852
rect 39300 9814 39352 9815
rect 39300 9780 39310 9814
rect 39310 9780 39344 9814
rect 39344 9780 39352 9814
rect 39300 9763 39352 9780
rect 40076 10212 40084 10225
rect 40084 10212 40118 10225
rect 40118 10212 40128 10225
rect 40076 10174 40128 10212
rect 40076 10173 40084 10174
rect 40084 10173 40118 10174
rect 40118 10173 40128 10174
rect 40076 10140 40084 10161
rect 40084 10140 40118 10161
rect 40118 10140 40128 10161
rect 40076 10109 40128 10140
rect 39818 9852 39826 9878
rect 39826 9852 39860 9878
rect 39860 9852 39870 9878
rect 39818 9826 39870 9852
rect 39818 9780 39826 9814
rect 39826 9780 39860 9814
rect 39860 9780 39870 9814
rect 39818 9762 39870 9780
rect 40590 10212 40600 10226
rect 40600 10212 40634 10226
rect 40634 10212 40642 10226
rect 40590 10174 40642 10212
rect 40590 10140 40600 10162
rect 40600 10140 40634 10162
rect 40634 10140 40642 10162
rect 40590 10110 40642 10140
rect 40335 9852 40342 9878
rect 40342 9852 40376 9878
rect 40376 9852 40387 9878
rect 40335 9826 40387 9852
rect 40335 9780 40342 9814
rect 40342 9780 40376 9814
rect 40376 9780 40387 9814
rect 40335 9762 40387 9780
rect 40850 9852 40858 9879
rect 40858 9852 40892 9879
rect 40892 9852 40902 9879
rect 40850 9827 40902 9852
rect 40850 9814 40902 9815
rect 40850 9780 40858 9814
rect 40858 9780 40892 9814
rect 40892 9780 40902 9814
rect 40850 9763 40902 9780
rect 24384 6788 24417 6808
rect 24417 6788 24436 6808
rect 24448 6788 24451 6808
rect 24451 6788 24489 6808
rect 24489 6788 24500 6808
rect 24384 6756 24436 6788
rect 24448 6756 24500 6788
rect 18894 6535 18918 6540
rect 18918 6535 19010 6540
rect 18894 6497 19010 6535
rect 18894 6463 18918 6497
rect 18918 6463 19010 6497
rect 18894 6425 19010 6463
rect 18894 6391 18918 6425
rect 18918 6391 19010 6425
rect 18894 6360 19010 6391
rect 25874 6822 25926 6828
rect 25938 6822 25990 6828
rect 25874 6788 25879 6822
rect 25879 6788 25917 6822
rect 25917 6788 25926 6822
rect 25938 6788 25951 6822
rect 25951 6788 25989 6822
rect 25989 6788 25990 6822
rect 25874 6776 25926 6788
rect 25938 6776 25990 6788
rect 23664 5730 23697 5763
rect 23697 5730 23716 5763
rect 23728 5730 23731 5763
rect 23731 5730 23769 5763
rect 23769 5730 23780 5763
rect 23664 5711 23716 5730
rect 23728 5711 23780 5730
rect 28035 6843 28036 6865
rect 28036 6843 28070 6865
rect 28070 6843 28087 6865
rect 28035 6813 28087 6843
rect 28035 6771 28036 6801
rect 28036 6771 28070 6801
rect 28070 6771 28087 6801
rect 28035 6749 28087 6771
rect 28035 6733 28087 6737
rect 28035 6699 28036 6733
rect 28036 6699 28070 6733
rect 28070 6699 28087 6733
rect 28035 6685 28087 6699
rect 28035 6661 28087 6673
rect 28035 6627 28036 6661
rect 28036 6627 28070 6661
rect 28070 6627 28087 6661
rect 28035 6621 28087 6627
rect 28035 6589 28087 6609
rect 28035 6557 28036 6589
rect 28036 6557 28070 6589
rect 28070 6557 28087 6589
rect 28035 6517 28087 6545
rect 28035 6493 28036 6517
rect 28036 6493 28070 6517
rect 28070 6493 28087 6517
rect 37612 6602 37623 6636
rect 37623 6602 37657 6636
rect 37657 6602 37664 6636
rect 37612 6584 37664 6602
rect 37612 6564 37664 6572
rect 37612 6530 37623 6564
rect 37623 6530 37657 6564
rect 37657 6530 37664 6564
rect 37612 6520 37664 6530
rect 37612 6492 37664 6508
rect 37612 6458 37623 6492
rect 37623 6458 37657 6492
rect 37657 6458 37664 6492
rect 37612 6456 37664 6458
rect 38319 7487 38328 7515
rect 38328 7487 38362 7515
rect 38362 7487 38371 7515
rect 38319 7463 38371 7487
rect 38319 7449 38371 7451
rect 38319 7415 38328 7449
rect 38328 7415 38362 7449
rect 38362 7415 38371 7449
rect 38319 7399 38371 7415
rect 38060 6623 38070 6638
rect 38070 6623 38104 6638
rect 38104 6623 38112 6638
rect 38060 6586 38112 6623
rect 38060 6551 38070 6574
rect 38070 6551 38104 6574
rect 38104 6551 38112 6574
rect 38060 6522 38112 6551
rect 38060 6479 38070 6510
rect 38070 6479 38104 6510
rect 38104 6479 38112 6510
rect 38060 6458 38112 6479
rect 38835 7089 38887 7112
rect 38835 7060 38844 7089
rect 38844 7060 38878 7089
rect 38878 7060 38887 7089
rect 38835 7017 38887 7048
rect 38835 6996 38844 7017
rect 38844 6996 38878 7017
rect 38878 6996 38887 7017
rect 38835 6983 38844 6984
rect 38844 6983 38878 6984
rect 38878 6983 38887 6984
rect 38835 6945 38887 6983
rect 38835 6932 38844 6945
rect 38844 6932 38878 6945
rect 38878 6932 38887 6945
rect 38577 6623 38586 6637
rect 38586 6623 38620 6637
rect 38620 6623 38629 6637
rect 38577 6585 38629 6623
rect 38577 6551 38586 6573
rect 38586 6551 38620 6573
rect 38620 6551 38629 6573
rect 38577 6521 38629 6551
rect 38577 6479 38586 6509
rect 38586 6479 38620 6509
rect 38620 6479 38629 6509
rect 38577 6457 38629 6479
rect 39351 7089 39403 7110
rect 39351 7058 39360 7089
rect 39360 7058 39394 7089
rect 39394 7058 39403 7089
rect 39351 7017 39403 7046
rect 39351 6994 39360 7017
rect 39360 6994 39394 7017
rect 39394 6994 39403 7017
rect 39351 6945 39403 6982
rect 39351 6930 39360 6945
rect 39360 6930 39394 6945
rect 39394 6930 39403 6945
rect 39093 6623 39102 6636
rect 39102 6623 39136 6636
rect 39136 6623 39145 6636
rect 39093 6585 39145 6623
rect 39093 6584 39102 6585
rect 39102 6584 39136 6585
rect 39136 6584 39145 6585
rect 39093 6551 39102 6572
rect 39102 6551 39136 6572
rect 39136 6551 39145 6572
rect 39093 6520 39145 6551
rect 39093 6479 39102 6508
rect 39102 6479 39136 6508
rect 39136 6479 39145 6508
rect 39093 6456 39145 6479
rect 39866 7055 39876 7078
rect 39876 7055 39910 7078
rect 39910 7055 39918 7078
rect 39866 7026 39918 7055
rect 39866 6983 39876 7014
rect 39876 6983 39910 7014
rect 39910 6983 39918 7014
rect 39866 6962 39918 6983
rect 39607 6623 39618 6637
rect 39618 6623 39652 6637
rect 39652 6623 39659 6637
rect 39607 6585 39659 6623
rect 39607 6551 39618 6573
rect 39618 6551 39652 6573
rect 39652 6551 39659 6573
rect 39607 6521 39659 6551
rect 39607 6479 39618 6509
rect 39618 6479 39652 6509
rect 39652 6479 39659 6509
rect 39607 6457 39659 6479
rect 40383 7089 40435 7111
rect 40383 7059 40392 7089
rect 40392 7059 40426 7089
rect 40426 7059 40435 7089
rect 40383 7017 40435 7047
rect 40383 6995 40392 7017
rect 40392 6995 40426 7017
rect 40426 6995 40435 7017
rect 40383 6945 40435 6983
rect 40383 6931 40392 6945
rect 40392 6931 40426 6945
rect 40426 6931 40435 6945
rect 41417 7487 41424 7514
rect 41424 7487 41458 7514
rect 41458 7487 41469 7514
rect 41417 7462 41469 7487
rect 41417 7449 41469 7450
rect 41417 7415 41424 7449
rect 41424 7415 41458 7449
rect 41458 7415 41469 7449
rect 41417 7398 41469 7415
rect 40125 6623 40134 6636
rect 40134 6623 40168 6636
rect 40168 6623 40177 6636
rect 40125 6585 40177 6623
rect 40125 6584 40134 6585
rect 40134 6584 40168 6585
rect 40168 6584 40177 6585
rect 40125 6551 40134 6572
rect 40134 6551 40168 6572
rect 40168 6551 40177 6572
rect 40125 6520 40177 6551
rect 40125 6479 40134 6508
rect 40134 6479 40168 6508
rect 40168 6479 40177 6508
rect 40125 6456 40177 6479
rect 40898 7089 40950 7109
rect 40898 7057 40908 7089
rect 40908 7057 40942 7089
rect 40942 7057 40950 7089
rect 40898 7017 40950 7045
rect 40898 6993 40908 7017
rect 40908 6993 40942 7017
rect 40942 6993 40950 7017
rect 40898 6945 40950 6981
rect 40898 6929 40908 6945
rect 40908 6929 40942 6945
rect 40942 6929 40950 6945
rect 40640 6623 40650 6637
rect 40650 6623 40684 6637
rect 40684 6623 40692 6637
rect 40640 6585 40692 6623
rect 40640 6551 40650 6573
rect 40650 6551 40684 6573
rect 40684 6551 40692 6573
rect 40640 6521 40692 6551
rect 40640 6479 40650 6509
rect 40650 6479 40684 6509
rect 40684 6479 40692 6509
rect 40640 6457 40692 6479
rect 43495 7779 44507 9815
rect 41157 6623 41166 6637
rect 41166 6623 41200 6637
rect 41200 6623 41209 6637
rect 41157 6585 41209 6623
rect 41157 6551 41166 6573
rect 41166 6551 41200 6573
rect 41200 6551 41209 6573
rect 41157 6521 41209 6551
rect 41157 6479 41166 6509
rect 41166 6479 41200 6509
rect 41200 6479 41209 6509
rect 41157 6457 41209 6479
rect 41930 7521 41982 7548
rect 41930 7496 41940 7521
rect 41940 7496 41974 7521
rect 41974 7496 41982 7521
rect 41930 7449 41982 7484
rect 41930 7432 41940 7449
rect 41940 7432 41974 7449
rect 41974 7432 41982 7449
rect 41930 7415 41940 7420
rect 41940 7415 41974 7420
rect 41974 7415 41982 7420
rect 41930 7377 41982 7415
rect 41930 7368 41940 7377
rect 41940 7368 41974 7377
rect 41974 7368 41982 7377
rect 41673 6623 41682 6637
rect 41682 6623 41716 6637
rect 41716 6623 41725 6637
rect 41673 6585 41725 6623
rect 41673 6551 41682 6573
rect 41682 6551 41716 6573
rect 41716 6551 41725 6573
rect 41673 6521 41725 6551
rect 41673 6479 41682 6509
rect 41682 6479 41716 6509
rect 41716 6479 41725 6509
rect 41673 6457 41725 6479
rect 42127 6601 42136 6635
rect 42136 6601 42170 6635
rect 42170 6601 42179 6635
rect 42127 6583 42179 6601
rect 42127 6563 42179 6571
rect 42127 6529 42136 6563
rect 42136 6529 42170 6563
rect 42170 6529 42179 6563
rect 42127 6519 42179 6529
rect 42127 6491 42179 6507
rect 42127 6457 42136 6491
rect 42136 6457 42170 6491
rect 42170 6457 42179 6491
rect 42127 6455 42179 6457
rect 25159 5730 25197 5758
rect 25197 5730 25211 5758
rect 25223 5730 25231 5758
rect 25231 5730 25269 5758
rect 25269 5730 25275 5758
rect 25159 5706 25211 5730
rect 25223 5706 25275 5730
rect 24379 4706 24431 4743
rect 24443 4706 24495 4743
rect 24379 4691 24417 4706
rect 24417 4691 24431 4706
rect 24443 4691 24451 4706
rect 24451 4691 24489 4706
rect 24489 4691 24495 4706
rect 12847 4209 22627 4230
rect 12847 3815 22627 4209
rect 12847 3794 22627 3815
rect 25869 4706 25921 4753
rect 25933 4706 25985 4753
rect 25869 4701 25879 4706
rect 25879 4701 25917 4706
rect 25917 4701 25921 4706
rect 25933 4701 25951 4706
rect 25951 4701 25985 4706
rect 23669 3648 23721 3678
rect 23733 3648 23785 3678
rect 23669 3626 23697 3648
rect 23697 3626 23721 3648
rect 23733 3626 23769 3648
rect 23769 3626 23785 3648
rect 25164 3648 25216 3678
rect 25228 3648 25280 3678
rect 25164 3626 25197 3648
rect 25197 3626 25216 3648
rect 25228 3626 25231 3648
rect 25231 3626 25269 3648
rect 25269 3626 25280 3648
rect 24384 3504 24436 3513
rect 24384 3470 24389 3504
rect 24389 3470 24423 3504
rect 24423 3470 24436 3504
rect 24384 3461 24436 3470
rect 24448 3504 24500 3513
rect 24448 3470 24461 3504
rect 24461 3470 24495 3504
rect 24495 3470 24500 3504
rect 24448 3461 24500 3470
rect 26705 3459 26864 3463
rect 26864 3459 26898 3463
rect 26898 3459 26949 3463
rect 26705 3421 26949 3459
rect 26705 3387 26864 3421
rect 26864 3387 26898 3421
rect 26898 3387 26949 3421
rect 26705 3349 26949 3387
rect 26705 3315 26864 3349
rect 26864 3315 26898 3349
rect 26898 3315 26949 3349
rect 26705 3277 26949 3315
rect 26705 3243 26864 3277
rect 26864 3243 26898 3277
rect 26898 3243 26949 3277
rect 26705 3205 26949 3243
rect 26705 3171 26864 3205
rect 26864 3171 26898 3205
rect 26898 3171 26949 3205
rect 26705 3133 26949 3171
rect 26705 3099 26864 3133
rect 26864 3099 26898 3133
rect 26898 3099 26949 3133
rect 26705 3091 26949 3099
rect -13051 2172 -12039 2928
rect 3722 2192 4734 2884
rect 32541 2922 33553 3678
rect 49314 2942 50326 3634
rect 10364 1473 11248 2357
rect -15192 8 -14308 764
rect 5895 51 6843 743
rect 30400 758 31284 1514
rect 51487 801 52435 1493
rect 8106 -1044 8990 -96
rect 12843 -992 22623 -172
<< metal2 >>
rect -10354 25430 -8968 25616
rect -10354 24654 -10189 25430
rect -9253 24654 -8968 25430
rect -10354 24520 -8968 24654
rect -268 25356 966 25380
rect -268 25216 970 25356
rect -268 24520 -115 25216
rect 821 24520 970 25216
rect -268 24374 970 24520
rect 8036 24833 9060 24867
rect -268 24366 966 24374
rect -15376 23971 -14114 24104
rect -15376 23151 -15293 23971
rect -14217 23151 -14114 23971
rect -15376 764 -14114 23151
rect 5764 23963 7026 24124
rect 5764 23207 5874 23963
rect 6886 23207 7026 23963
rect -13156 22132 -11894 22289
rect -13156 21376 -13012 22132
rect -12000 21376 -11894 22132
rect -13156 2928 -11894 21376
rect -4350 22200 -3490 22289
rect -4350 21344 -4268 22200
rect -3572 21344 -3490 22200
rect -4350 21265 -3490 21344
rect 3606 22198 4868 22290
rect 3606 21378 3696 22198
rect 4772 21378 4868 22198
rect -4092 18466 -3798 18499
rect -4092 18286 -4069 18466
rect -3825 18286 -3798 18466
rect -2036 18454 -1830 18502
rect -2036 18416 -1993 18454
rect -4092 18253 -3798 18286
rect -2038 18338 -1993 18416
rect -1877 18416 -1830 18454
rect -1877 18338 -1828 18416
rect -2038 18258 -1828 18338
rect -2719 18099 -2589 18105
rect -2210 18099 -2080 18105
rect -2036 18099 -1830 18258
rect -1695 18099 -1565 18101
rect -2719 18097 -592 18099
rect -2719 18075 -535 18097
rect -2719 18023 -2682 18075
rect -2630 18023 -2173 18075
rect -2121 18071 -535 18075
rect -2121 18023 -1658 18071
rect -2719 18019 -1658 18023
rect -1606 18067 -535 18071
rect -1606 18063 -628 18067
rect -1606 18019 -1139 18063
rect -2719 18011 -1139 18019
rect -1087 18015 -628 18063
rect -576 18015 -535 18067
rect -1087 18011 -535 18015
rect -2719 17959 -2682 18011
rect -2630 17959 -2173 18011
rect -2121 18007 -535 18011
rect -2121 17959 -1658 18007
rect -2719 17955 -1658 17959
rect -1606 18003 -535 18007
rect -1606 17999 -628 18003
rect -1606 17955 -1139 17999
rect -2719 17947 -1139 17955
rect -1087 17951 -628 17999
rect -576 17951 -535 18003
rect -1087 17947 -535 17951
rect -2719 17895 -2682 17947
rect -2630 17895 -2173 17947
rect -2121 17943 -535 17947
rect -2121 17895 -1658 17943
rect -2719 17891 -1658 17895
rect -1606 17939 -535 17943
rect -1606 17935 -628 17939
rect -1606 17891 -1139 17935
rect -2719 17883 -1139 17891
rect -1087 17887 -628 17935
rect -576 17887 -535 17939
rect -1087 17883 -535 17887
rect -2719 17864 -535 17883
rect -2701 17861 -535 17864
rect -2036 17860 -1830 17861
rect -1695 17860 -1565 17861
rect -1176 17852 -1046 17861
rect -665 17856 -535 17861
rect -6276 17550 -6096 17594
rect -6276 17498 -6244 17550
rect -6192 17498 -6180 17550
rect -6128 17498 -6096 17550
rect -6276 17454 -6096 17498
rect -6246 17175 -6116 17454
rect -6246 17123 -6207 17175
rect -6155 17123 -6116 17175
rect -6246 17084 -6116 17123
rect -5936 16367 -5626 16394
rect -919 16373 -789 16374
rect -15 16373 241 16377
rect -2959 16368 241 16373
rect -5936 16337 -5866 16367
rect -5686 16337 -5626 16367
rect -5936 16281 -5884 16337
rect -5668 16281 -5626 16337
rect -5936 16251 -5866 16281
rect -5686 16251 -5626 16281
rect -5936 16224 -5626 16251
rect -2971 16350 241 16368
rect -2971 16338 -2870 16350
rect -2971 16286 -2934 16338
rect -2882 16294 -2870 16338
rect -2814 16344 241 16350
rect -2814 16341 -882 16344
rect -2814 16340 -1404 16341
rect -2814 16334 -1920 16340
rect -2814 16294 -2434 16334
rect -2882 16286 -2434 16294
rect -2971 16282 -2434 16286
rect -2382 16288 -1920 16334
rect -1868 16289 -1404 16340
rect -1352 16292 -882 16341
rect -830 16341 241 16344
rect -830 16338 23 16341
rect -830 16292 -376 16338
rect -1352 16289 -376 16292
rect -1868 16288 -376 16289
rect -2382 16286 -376 16288
rect -324 16286 23 16338
rect -2382 16282 23 16286
rect -2971 16280 23 16282
rect -2971 16277 -882 16280
rect -2971 16276 -1404 16277
rect -2971 16274 -1920 16276
rect -2971 16222 -2934 16274
rect -2882 16270 -1920 16274
rect -2882 16222 -2870 16270
rect -2971 16214 -2870 16222
rect -2814 16218 -2434 16270
rect -2382 16224 -1920 16270
rect -1868 16225 -1404 16276
rect -1352 16228 -882 16277
rect -830 16274 23 16280
rect -830 16228 -376 16274
rect -1352 16225 -376 16228
rect -1868 16224 -376 16225
rect -2382 16222 -376 16224
rect -324 16222 23 16274
rect -2382 16218 23 16222
rect -2814 16216 23 16218
rect -2814 16214 -882 16216
rect -2971 16213 -882 16214
rect -2971 16212 -1404 16213
rect -2971 16210 -1920 16212
rect -6436 16105 -6196 16184
rect -2971 16158 -2934 16210
rect -2882 16206 -1920 16210
rect -2882 16190 -2434 16206
rect -2882 16158 -2870 16190
rect -2971 16134 -2870 16158
rect -2814 16154 -2434 16190
rect -2382 16160 -1920 16206
rect -1868 16161 -1404 16212
rect -1352 16164 -882 16213
rect -830 16210 23 16216
rect -830 16164 -376 16210
rect -1352 16161 -376 16164
rect -1868 16160 -376 16161
rect -2382 16158 -376 16160
rect -324 16161 23 16210
rect 203 16161 241 16341
rect -324 16158 241 16161
rect -2382 16154 241 16158
rect -2814 16134 241 16154
rect -2971 16128 241 16134
rect -2971 16127 -2756 16128
rect -2918 16113 -2756 16127
rect -2471 16123 -2341 16128
rect -413 16127 -283 16128
rect -15 16127 241 16128
rect -6436 16053 -6369 16105
rect -6317 16053 -6305 16105
rect -6253 16053 -6196 16105
rect -6436 14828 -6196 16053
rect -5466 14944 -5226 15344
rect -4244 15200 -4068 15218
rect -4244 15178 -4214 15200
rect -4098 15178 -4068 15200
rect -4244 15042 -4224 15178
rect -4088 15042 -4068 15178
rect -4244 15020 -4214 15042
rect -4098 15020 -4068 15042
rect -4244 15002 -4068 15020
rect -5466 14892 -5437 14944
rect -5385 14892 -5373 14944
rect -5321 14892 -5309 14944
rect -5257 14892 -5226 14944
rect -5466 14874 -5226 14892
rect -6952 14822 -4835 14828
rect -6994 14809 -4835 14822
rect -6994 14768 -4796 14809
rect -6994 14716 -6947 14768
rect -6895 14755 -4796 14768
rect -6895 14716 -5936 14755
rect -6994 14704 -5936 14716
rect -6994 14652 -6947 14704
rect -6895 14703 -5936 14704
rect -5884 14703 -4899 14755
rect -4847 14703 -4796 14755
rect -6895 14691 -4796 14703
rect -6895 14652 -5936 14691
rect -6994 14640 -5936 14652
rect -6994 14588 -6947 14640
rect -6895 14639 -5936 14640
rect -5884 14639 -4899 14691
rect -4847 14639 -4796 14691
rect -6895 14627 -4796 14639
rect -6895 14588 -5936 14627
rect -6994 14575 -5936 14588
rect -5884 14575 -4899 14627
rect -4847 14575 -4796 14627
rect -6994 14536 -4796 14575
rect -6952 14532 -4796 14536
rect -6436 14524 -6196 14532
rect -5983 14523 -5833 14532
rect -4946 14523 -4796 14532
rect -6481 13127 -6331 13130
rect -5451 13127 -5301 13140
rect -7463 13119 -5301 13127
rect -7500 13097 -5301 13119
rect -7500 13076 -5884 13097
rect -7500 13065 -6434 13076
rect -7500 13013 -7453 13065
rect -7401 13024 -6434 13065
rect -6382 13024 -5884 13076
rect -7401 13013 -5884 13024
rect -7500 13012 -5884 13013
rect -7500 13001 -6434 13012
rect -7500 12949 -7453 13001
rect -7401 12960 -6434 13001
rect -6382 12960 -5884 13012
rect -7401 12949 -5884 12960
rect -7500 12948 -5884 12949
rect -7500 12937 -6434 12948
rect -7500 12885 -7453 12937
rect -7401 12896 -6434 12937
rect -6382 12896 -5884 12948
rect -7401 12885 -5884 12896
rect -7500 12881 -5884 12885
rect -5668 13086 -5301 13097
rect -5668 13034 -5404 13086
rect -5352 13034 -5301 13086
rect -5668 13022 -5301 13034
rect -5668 12970 -5404 13022
rect -5352 12970 -5301 13022
rect -5668 12958 -5301 12970
rect -5668 12906 -5404 12958
rect -5352 12906 -5301 12958
rect -5668 12881 -5301 12906
rect -7500 12854 -5301 12881
rect -7500 12841 -5352 12854
rect -7500 12833 -7350 12841
rect -3939 12823 -3774 12875
rect -3939 12821 -3888 12823
rect -3832 12821 -3774 12823
rect -6872 12769 -6698 12787
rect -6872 12713 -6855 12769
rect -6799 12767 -6775 12769
rect -6793 12715 -6781 12767
rect -6799 12713 -6775 12715
rect -6719 12713 -6698 12769
rect -6872 12701 -6698 12713
rect -5382 12644 -4756 12676
rect -5382 12428 -5333 12644
rect -4797 12428 -4756 12644
rect -5382 12400 -4756 12428
rect -3939 12449 -3918 12821
rect -3802 12449 -3774 12821
rect -3939 12447 -3888 12449
rect -3832 12447 -3774 12449
rect -3939 12404 -3774 12447
rect -8591 10766 -3849 10773
rect -8591 10714 -8566 10766
rect -8514 10734 -3849 10766
rect -8514 10733 -4225 10734
rect -8514 10714 -8051 10733
rect -8591 10702 -8051 10714
rect -8591 10650 -8566 10702
rect -8514 10681 -8051 10702
rect -7999 10732 -7018 10733
rect -7999 10681 -7534 10732
rect -8514 10680 -7534 10681
rect -7482 10681 -7018 10732
rect -6966 10732 -4225 10733
rect -6966 10731 -5986 10732
rect -6966 10681 -6502 10731
rect -7482 10680 -6502 10681
rect -8514 10679 -6502 10680
rect -6450 10680 -5986 10731
rect -5934 10731 -4954 10732
rect -5934 10680 -5470 10731
rect -6450 10679 -5470 10680
rect -5418 10680 -4954 10731
rect -4902 10680 -4438 10732
rect -4386 10680 -4225 10732
rect -5418 10679 -4225 10680
rect -8514 10678 -4225 10679
rect -4169 10678 -4145 10734
rect -4089 10732 -3849 10734
rect -4089 10680 -3922 10732
rect -3870 10680 -3849 10732
rect -4089 10678 -3849 10680
rect -8514 10650 -3849 10678
rect -8591 10640 -3849 10650
rect -10054 10492 -9276 10556
rect -10054 9928 -9976 10492
rect -9412 9928 -9276 10492
rect -8856 10489 -3596 10501
rect -8856 10488 -6243 10489
rect -8856 10486 -8308 10488
rect -8856 10434 -8824 10486
rect -8772 10436 -8308 10486
rect -8256 10436 -7792 10488
rect -7740 10487 -6760 10488
rect -7740 10436 -7276 10487
rect -8772 10435 -7276 10436
rect -7224 10436 -6760 10487
rect -6708 10437 -6243 10488
rect -6191 10488 -3596 10489
rect -6191 10487 -4696 10488
rect -6191 10486 -5213 10487
rect -6191 10456 -5728 10486
rect -6191 10437 -6032 10456
rect -6708 10436 -6032 10437
rect -7224 10435 -6032 10436
rect -8772 10434 -6032 10435
rect -8856 10425 -6032 10434
rect -8856 10424 -6243 10425
rect -8856 10422 -8308 10424
rect -8856 10370 -8824 10422
rect -8772 10372 -8308 10422
rect -8256 10372 -7792 10424
rect -7740 10423 -6760 10424
rect -7740 10372 -7276 10423
rect -8772 10371 -7276 10372
rect -7224 10372 -6760 10423
rect -6708 10373 -6243 10424
rect -6191 10400 -6032 10425
rect -5976 10400 -5952 10456
rect -5896 10434 -5728 10456
rect -5676 10435 -5213 10486
rect -5161 10436 -4696 10487
rect -4644 10487 -3596 10488
rect -4644 10436 -4180 10487
rect -5161 10435 -4180 10436
rect -4128 10435 -3664 10487
rect -3612 10435 -3596 10487
rect -5676 10434 -3596 10435
rect -5896 10424 -3596 10434
rect -5896 10423 -4696 10424
rect -5896 10422 -5213 10423
rect -5896 10400 -5728 10422
rect -6191 10373 -5728 10400
rect -6708 10372 -5728 10373
rect -7224 10371 -5728 10372
rect -8772 10370 -5728 10371
rect -5676 10371 -5213 10422
rect -5161 10372 -4696 10423
rect -4644 10423 -3596 10424
rect -4644 10372 -4180 10423
rect -5161 10371 -4180 10372
rect -4128 10371 -3664 10423
rect -3612 10371 -3596 10423
rect -5676 10370 -3596 10371
rect -8856 10359 -3596 10370
rect -10054 9882 -9276 9928
rect -7088 9478 -4925 9495
rect -7088 9426 -7065 9478
rect -7013 9477 -4925 9478
rect -7013 9475 -6033 9477
rect -7013 9447 -6549 9475
rect -7013 9426 -6850 9447
rect -7088 9414 -6850 9426
rect -7088 9362 -7065 9414
rect -7013 9391 -6850 9414
rect -6794 9391 -6770 9447
rect -6714 9423 -6549 9447
rect -6497 9425 -6033 9475
rect -5981 9476 -4925 9477
rect -5981 9475 -5002 9476
rect -5981 9425 -5516 9475
rect -6497 9423 -5516 9425
rect -5464 9424 -5002 9475
rect -4950 9424 -4925 9476
rect -5464 9423 -4925 9424
rect -6714 9413 -4925 9423
rect -6714 9411 -6033 9413
rect -6714 9391 -6549 9411
rect -7013 9362 -6549 9391
rect -7088 9359 -6549 9362
rect -6497 9361 -6033 9411
rect -5981 9412 -4925 9413
rect -5981 9411 -5002 9412
rect -5981 9361 -5516 9411
rect -6497 9359 -5516 9361
rect -5464 9360 -5002 9411
rect -4950 9360 -4925 9412
rect -5464 9359 -4925 9360
rect -7088 9343 -4925 9359
rect -7335 9138 -4674 9164
rect -7335 9128 -7029 9138
rect -7335 9076 -7322 9128
rect -7270 9082 -7029 9128
rect -6973 9129 -4674 9138
rect -6973 9127 -6292 9129
rect -6973 9082 -6805 9127
rect -7270 9076 -6805 9082
rect -7335 9075 -6805 9076
rect -6753 9077 -6292 9127
rect -6240 9128 -4742 9129
rect -6240 9077 -5774 9128
rect -6753 9076 -5774 9077
rect -5722 9076 -5257 9128
rect -5205 9077 -4742 9128
rect -4690 9077 -4674 9129
rect -5205 9076 -4674 9077
rect -6753 9075 -4674 9076
rect -7335 9065 -4674 9075
rect -7335 9064 -6292 9065
rect -7335 9012 -7322 9064
rect -7270 9063 -6292 9064
rect -7270 9058 -6805 9063
rect -7270 9012 -7029 9058
rect -7335 9002 -7029 9012
rect -6973 9011 -6805 9058
rect -6753 9013 -6292 9063
rect -6240 9064 -4742 9065
rect -6240 9013 -5774 9064
rect -6753 9012 -5774 9013
rect -5722 9012 -5257 9064
rect -5205 9013 -4742 9064
rect -4690 9013 -4674 9065
rect -5205 9012 -4674 9013
rect -6753 9011 -4674 9012
rect -6973 9002 -4674 9011
rect -7335 8979 -4674 9002
rect -7317 6798 -3582 6811
rect -7317 6776 -3662 6798
rect -7317 6765 -7030 6776
rect -7317 6713 -7273 6765
rect -7221 6720 -7030 6765
rect -6974 6764 -3662 6776
rect -6974 6720 -4175 6764
rect -7221 6713 -4175 6720
rect -7317 6712 -4175 6713
rect -4123 6746 -3662 6764
rect -3610 6746 -3582 6798
rect -4123 6734 -3582 6746
rect -4123 6712 -3662 6734
rect -7317 6701 -3662 6712
rect -7317 6649 -7273 6701
rect -7221 6700 -3662 6701
rect -7221 6696 -4175 6700
rect -7221 6649 -7030 6696
rect -7317 6640 -7030 6649
rect -6974 6648 -4175 6696
rect -4123 6682 -3662 6700
rect -3610 6682 -3582 6734
rect -4123 6670 -3582 6682
rect -4123 6648 -3662 6670
rect -6974 6640 -3662 6648
rect -7317 6618 -3662 6640
rect -3610 6618 -3582 6670
rect -7317 6606 -3582 6618
rect -6790 6362 -4598 6375
rect -6790 6310 -6757 6362
rect -6705 6361 -4598 6362
rect -6705 6360 -5209 6361
rect -6705 6310 -6241 6360
rect -6790 6308 -6241 6310
rect -6189 6336 -5209 6360
rect -6189 6308 -6031 6336
rect -6790 6298 -6031 6308
rect -6790 6246 -6757 6298
rect -6705 6296 -6031 6298
rect -6705 6246 -6241 6296
rect -6790 6244 -6241 6246
rect -6189 6244 -6031 6296
rect -6790 6234 -6031 6244
rect -6790 6182 -6757 6234
rect -6705 6232 -6031 6234
rect -6705 6182 -6241 6232
rect -6790 6180 -6241 6182
rect -6189 6200 -6031 6232
rect -5895 6328 -5209 6336
rect -5895 6276 -5726 6328
rect -5674 6309 -5209 6328
rect -5157 6359 -4598 6361
rect -5157 6309 -4694 6359
rect -5674 6307 -4694 6309
rect -4642 6307 -4598 6359
rect -5674 6297 -4598 6307
rect -5674 6276 -5209 6297
rect -5895 6264 -5209 6276
rect -5895 6212 -5726 6264
rect -5674 6245 -5209 6264
rect -5157 6295 -4598 6297
rect -5157 6245 -4694 6295
rect -5674 6243 -4694 6245
rect -4642 6243 -4598 6295
rect -5674 6233 -4598 6243
rect -5674 6212 -5209 6233
rect -5895 6200 -5209 6212
rect -6189 6181 -5209 6200
rect -5157 6231 -4598 6233
rect -5157 6181 -4694 6231
rect -6189 6180 -4694 6181
rect -6790 6179 -4694 6180
rect -4642 6179 -4598 6231
rect -6790 6168 -4598 6179
rect -7997 5888 -3384 5901
rect -7997 5886 -7532 5888
rect -7997 5834 -7980 5886
rect -7928 5836 -7532 5886
rect -7480 5887 -3384 5888
rect -7480 5836 -7015 5887
rect -7928 5835 -7015 5836
rect -6963 5886 -5985 5887
rect -6963 5835 -6499 5886
rect -7928 5834 -6499 5835
rect -6447 5835 -5985 5886
rect -5933 5886 -4952 5887
rect -5933 5835 -5467 5886
rect -6447 5834 -5467 5835
rect -5415 5835 -4952 5886
rect -4900 5835 -4435 5887
rect -4383 5835 -3919 5887
rect -3867 5885 -3384 5887
rect -3867 5835 -3465 5885
rect -5415 5834 -3465 5835
rect -7997 5833 -3465 5834
rect -3413 5833 -3384 5885
rect -7997 5824 -3384 5833
rect -7997 5822 -7532 5824
rect -7997 5770 -7980 5822
rect -7928 5772 -7532 5822
rect -7480 5823 -3384 5824
rect -7480 5772 -7015 5823
rect -7928 5771 -7015 5772
rect -6963 5822 -5985 5823
rect -6963 5771 -6499 5822
rect -7928 5770 -6499 5771
rect -6447 5771 -5985 5822
rect -5933 5822 -4952 5823
rect -5933 5771 -5467 5822
rect -6447 5770 -5467 5771
rect -5415 5771 -4952 5822
rect -4900 5771 -4435 5823
rect -4383 5771 -3919 5823
rect -3867 5821 -3384 5823
rect -3867 5771 -3465 5821
rect -5415 5770 -3465 5771
rect -7997 5769 -3465 5770
rect -3413 5769 -3384 5821
rect -7997 5760 -3384 5769
rect -7997 5758 -7532 5760
rect -7997 5706 -7980 5758
rect -7928 5708 -7532 5758
rect -7480 5759 -3384 5760
rect -7480 5708 -7015 5759
rect -7928 5707 -7015 5708
rect -6963 5758 -5985 5759
rect -6963 5707 -6499 5758
rect -7928 5706 -6499 5707
rect -6447 5707 -5985 5758
rect -5933 5758 -4952 5759
rect -5933 5707 -5467 5758
rect -6447 5706 -5467 5707
rect -5415 5707 -4952 5758
rect -4900 5707 -4435 5759
rect -4383 5707 -3919 5759
rect -3867 5757 -3384 5759
rect -3867 5707 -3465 5757
rect -5415 5706 -3465 5707
rect -7997 5705 -3465 5706
rect -3413 5705 -3384 5757
rect -7997 5693 -3384 5705
rect -3853 5692 -3384 5693
rect -13156 2172 -13051 2928
rect -12039 2172 -11894 2928
rect -13156 2061 -11894 2172
rect 3606 2884 4868 21378
rect 3606 2192 3722 2884
rect 4734 2192 4868 2884
rect 3606 2064 4868 2192
rect -15376 8 -15192 764
rect -14308 8 -14114 764
rect -15376 -106 -14114 8
rect 5764 743 7026 23207
rect 5764 51 5895 743
rect 6843 51 7026 743
rect 8036 23885 8103 24833
rect 8987 23885 9060 24833
rect 8036 742 9060 23885
rect 30216 24721 31478 24854
rect 30216 23901 30299 24721
rect 31375 23901 31478 24721
rect 10298 23002 11322 23039
rect 10298 22054 10363 23002
rect 11247 22054 11322 23002
rect 10298 17054 11322 22054
rect 24680 18659 26854 18698
rect 24680 18655 26798 18659
rect 24680 18603 24684 18655
rect 24736 18607 26798 18655
rect 26850 18607 26854 18659
rect 24736 18603 26854 18607
rect 24680 18595 26854 18603
rect 24680 18591 26798 18595
rect 24680 18539 24684 18591
rect 24736 18543 26798 18591
rect 26850 18543 26854 18595
rect 24736 18539 26854 18543
rect 24680 18531 26854 18539
rect 24680 18527 26798 18531
rect 24680 18475 24684 18527
rect 24736 18479 26798 18527
rect 26850 18479 26854 18531
rect 24736 18475 26854 18479
rect 24680 18467 26854 18475
rect 24680 18463 26798 18467
rect 24680 18411 24684 18463
rect 24736 18415 26798 18463
rect 26850 18415 26854 18467
rect 24736 18411 26854 18415
rect 24680 18403 26854 18411
rect 24680 18399 26798 18403
rect 24680 18347 24684 18399
rect 24736 18351 26798 18399
rect 26850 18351 26854 18403
rect 24736 18347 26854 18351
rect 24680 18306 26854 18347
rect 25738 17557 27912 17596
rect 25738 17505 25741 17557
rect 25793 17555 27912 17557
rect 25793 17505 27855 17555
rect 25738 17503 27855 17505
rect 27907 17503 27912 17555
rect 25738 17493 27912 17503
rect 25738 17441 25741 17493
rect 25793 17491 27912 17493
rect 25793 17441 27855 17491
rect 25738 17439 27855 17441
rect 27907 17439 27912 17491
rect 25738 17429 27912 17439
rect 25738 17377 25741 17429
rect 25793 17427 27912 17429
rect 25793 17377 27855 17427
rect 25738 17375 27855 17377
rect 27907 17375 27912 17427
rect 25738 17365 27912 17375
rect 25738 17313 25741 17365
rect 25793 17363 27912 17365
rect 25793 17313 27855 17363
rect 25738 17311 27855 17313
rect 27907 17311 27912 17363
rect 25738 17301 27912 17311
rect 25738 17249 25741 17301
rect 25793 17299 27912 17301
rect 25793 17249 27855 17299
rect 25738 17247 27855 17249
rect 27907 17247 27912 17299
rect 25738 17208 27912 17247
rect 10298 15018 10333 17054
rect 11281 15018 11322 17054
rect 27888 16812 28098 16828
rect 27888 16798 27939 16812
rect 28055 16798 28098 16812
rect 27888 16262 27929 16798
rect 28065 16262 28098 16798
rect 27888 16248 27939 16262
rect 28055 16248 28098 16262
rect 27888 16222 28098 16248
rect 10298 2357 11322 15018
rect 22522 16117 22962 16152
rect 22522 15745 22553 16117
rect 22925 15745 22962 16117
rect 13932 14509 15772 14530
rect 13932 14201 13982 14509
rect 14162 14201 15609 14509
rect 15725 14201 15772 14509
rect 13932 14180 15772 14201
rect 22522 14168 22962 15745
rect 29188 15217 29438 15286
rect 29188 14841 29243 15217
rect 29379 14841 29438 15217
rect 29188 14748 29438 14841
rect 22522 14099 28190 14168
rect 19900 13882 20312 13910
rect 22522 13882 27809 14099
rect 19890 13871 27809 13882
rect 19890 13499 19933 13871
rect 20305 13803 27809 13871
rect 28105 13803 28190 14099
rect 20305 13728 28190 13803
rect 20305 13499 22962 13728
rect 19890 13442 22962 13499
rect 24792 13348 24912 13352
rect 24792 13296 24826 13348
rect 24878 13296 24912 13348
rect 15942 12351 17262 12400
rect 12982 12052 15142 12100
rect 12982 11808 13014 12052
rect 13130 11808 14999 12052
rect 15115 11808 15142 12052
rect 12982 11770 15142 11808
rect 15942 11979 17104 12351
rect 17220 11979 17262 12351
rect 15942 11930 17262 11979
rect 18466 12119 18646 12154
rect 18466 11939 18498 12119
rect 18614 11939 18646 12119
rect 13198 10863 13662 10942
rect 13198 10555 13276 10863
rect 13584 10555 13662 10863
rect 13198 10496 13662 10555
rect 13194 9356 13644 9424
rect 13194 9048 13262 9356
rect 13570 9048 13644 9356
rect 13194 8988 13644 9048
rect 14157 7930 14507 11770
rect 15942 11182 16162 11930
rect 17510 11462 17962 11498
rect 17510 11430 17545 11462
rect 16922 11391 17545 11430
rect 16922 11339 16956 11391
rect 17008 11339 17545 11391
rect 16922 11326 17545 11339
rect 17921 11326 17962 11462
rect 16922 11324 17626 11326
rect 17678 11324 17962 11326
rect 16922 11290 17962 11324
rect 15942 10938 15989 11182
rect 16105 10938 16162 11182
rect 15942 10890 16162 10938
rect 18466 11129 18646 11939
rect 18466 10949 18498 11129
rect 18614 10949 18646 11129
rect 18466 10904 18646 10949
rect 24792 11243 24912 13296
rect 26152 13314 26912 13322
rect 26152 13298 27004 13314
rect 26152 12926 26697 13298
rect 26877 12926 27004 13298
rect 26152 12902 27004 12926
rect 24792 11191 24826 11243
rect 24878 11191 24912 11243
rect 22632 10391 23060 10446
rect 21088 9346 21302 9398
rect 21088 9340 21137 9346
rect 21253 9340 21302 9346
rect 21088 9044 21127 9340
rect 21263 9044 21302 9340
rect 22632 9251 22655 10391
rect 23027 9251 23060 10391
rect 22632 9202 23060 9251
rect 21088 9038 21137 9044
rect 21253 9038 21302 9044
rect 21088 8994 21302 9038
rect 14932 8676 17122 8700
rect 14932 8304 14979 8676
rect 15095 8304 16959 8676
rect 17075 8304 17122 8676
rect 14932 8270 17122 8304
rect 17446 8638 19636 8674
rect 17446 8330 17468 8638
rect 17584 8636 19478 8638
rect 17584 8340 17726 8636
rect 18182 8340 19478 8636
rect 17584 8330 19478 8340
rect 19594 8330 19636 8638
rect 17446 8294 19636 8330
rect 22785 8208 23011 9202
rect 24792 9138 24912 11191
rect 25632 12298 25762 12312
rect 25632 12246 25666 12298
rect 25718 12246 25762 12298
rect 25632 12241 25762 12246
rect 26154 12241 26571 12902
rect 25632 11824 26571 12241
rect 25632 10198 25762 11824
rect 25632 10146 25671 10198
rect 25723 10146 25762 10198
rect 25632 10132 25762 10146
rect 24792 9086 24826 9138
rect 24878 9086 24912 9138
rect 24792 9072 24912 9086
rect 16902 8187 23011 8208
rect 16902 8007 16922 8187
rect 17038 8166 23011 8187
rect 17038 8114 17885 8166
rect 17937 8114 17949 8166
rect 18001 8114 18013 8166
rect 18065 8114 18077 8166
rect 18129 8114 23011 8166
rect 17038 8007 23011 8114
rect 16902 7982 23011 8007
rect 26182 8427 26382 8462
rect 26182 8421 26222 8427
rect 26338 8421 26382 8427
rect 14157 7877 17082 7930
rect 14157 7633 16872 7877
rect 17052 7633 17082 7877
rect 14157 7580 17082 7633
rect 17862 7240 18152 7982
rect 17422 7180 18152 7240
rect 17422 7000 17455 7180
rect 17699 7000 18152 7180
rect 17422 6940 18152 7000
rect 23642 7873 23812 7912
rect 23642 7821 23664 7873
rect 23716 7821 23728 7873
rect 23780 7821 23812 7873
rect 23642 7772 23812 7821
rect 25142 7863 25302 7892
rect 25142 7811 25164 7863
rect 25216 7811 25228 7863
rect 25280 7811 25302 7863
rect 25142 7772 25302 7811
rect 23642 7492 25302 7772
rect 16423 6600 17064 6606
rect 16423 6540 19042 6600
rect 16423 6539 18894 6540
rect 16423 6359 16436 6539
rect 16616 6360 18894 6539
rect 19010 6360 19042 6540
rect 16616 6359 19042 6360
rect 16423 6316 19042 6359
rect 16759 6310 19042 6316
rect 23642 5763 23812 7492
rect 23642 5711 23664 5763
rect 23716 5711 23728 5763
rect 23780 5711 23812 5763
rect 10298 1473 10364 2357
rect 11248 1473 11322 2357
rect 10298 1402 11322 1473
rect 12752 4230 22754 4306
rect 12752 3794 12847 4230
rect 22627 3794 22754 4230
rect 5764 -101 7026 51
rect 8038 -96 9059 742
rect 12752 -16 22754 3794
rect 23642 3678 23812 5711
rect 23642 3626 23669 3678
rect 23721 3626 23733 3678
rect 23785 3626 23812 3678
rect 23642 3612 23812 3626
rect 24362 6808 24522 6832
rect 24362 6756 24384 6808
rect 24436 6756 24448 6808
rect 24500 6756 24522 6808
rect 24362 4743 24522 6756
rect 24362 4691 24379 4743
rect 24431 4691 24443 4743
rect 24495 4691 24522 4743
rect 24362 3513 24522 4691
rect 25142 5758 25302 7492
rect 26182 7485 26212 8421
rect 26348 7485 26382 8421
rect 26182 7479 26222 7485
rect 26338 7479 26382 7485
rect 26182 7452 26382 7479
rect 26678 7591 27004 12902
rect 26678 7265 28213 7591
rect 27887 6865 28213 7265
rect 25142 5706 25159 5758
rect 25211 5706 25223 5758
rect 25275 5706 25302 5758
rect 25142 3678 25302 5706
rect 25852 6828 26012 6842
rect 25852 6776 25874 6828
rect 25926 6776 25938 6828
rect 25990 6776 26012 6828
rect 25852 5242 26012 6776
rect 27887 6813 28035 6865
rect 28087 6813 28213 6865
rect 27887 6801 28213 6813
rect 27887 6749 28035 6801
rect 28087 6749 28213 6801
rect 27887 6737 28213 6749
rect 27887 6685 28035 6737
rect 28087 6685 28213 6737
rect 27887 6673 28213 6685
rect 27887 6621 28035 6673
rect 28087 6621 28213 6673
rect 27887 6609 28213 6621
rect 27887 6557 28035 6609
rect 28087 6557 28213 6609
rect 27887 6545 28213 6557
rect 27887 6493 28035 6545
rect 28087 6493 28213 6545
rect 27887 6467 28213 6493
rect 25852 4812 27012 5242
rect 25852 4753 26012 4812
rect 25852 4701 25869 4753
rect 25921 4701 25933 4753
rect 25985 4701 26012 4753
rect 25852 4672 26012 4701
rect 25142 3626 25164 3678
rect 25216 3626 25228 3678
rect 25280 3626 25302 3678
rect 25142 3602 25302 3626
rect 24362 3461 24384 3513
rect 24436 3461 24448 3513
rect 24500 3461 24522 3513
rect 24362 3422 24522 3461
rect 26652 3463 27012 4812
rect 26652 3091 26705 3463
rect 26949 3091 27012 3463
rect 26652 3072 27012 3091
rect 30216 1514 31478 23901
rect 51356 24713 52618 24874
rect 51356 23957 51466 24713
rect 52478 23957 52618 24713
rect 32436 22882 33698 23039
rect 32436 22126 32580 22882
rect 33592 22126 33698 22882
rect 32436 3678 33698 22126
rect 41242 22950 42102 23039
rect 41242 22094 41324 22950
rect 42020 22094 42102 22950
rect 41242 22015 42102 22094
rect 49198 22948 50460 23040
rect 49198 22128 49288 22948
rect 50364 22128 50460 22948
rect 41500 19216 41794 19249
rect 41500 19036 41523 19216
rect 41767 19036 41794 19216
rect 43556 19204 43762 19252
rect 43556 19166 43599 19204
rect 41500 19003 41794 19036
rect 43554 19088 43599 19166
rect 43715 19166 43762 19204
rect 43715 19088 43764 19166
rect 43554 19008 43764 19088
rect 42873 18849 43003 18855
rect 43382 18849 43512 18855
rect 43556 18849 43762 19008
rect 43897 18849 44027 18851
rect 42873 18847 45000 18849
rect 42873 18825 45057 18847
rect 42873 18773 42910 18825
rect 42962 18773 43419 18825
rect 43471 18821 45057 18825
rect 43471 18773 43934 18821
rect 42873 18769 43934 18773
rect 43986 18817 45057 18821
rect 43986 18813 44964 18817
rect 43986 18769 44453 18813
rect 42873 18761 44453 18769
rect 44505 18765 44964 18813
rect 45016 18765 45057 18817
rect 44505 18761 45057 18765
rect 42873 18709 42910 18761
rect 42962 18709 43419 18761
rect 43471 18757 45057 18761
rect 43471 18709 43934 18757
rect 42873 18705 43934 18709
rect 43986 18753 45057 18757
rect 43986 18749 44964 18753
rect 43986 18705 44453 18749
rect 42873 18697 44453 18705
rect 44505 18701 44964 18749
rect 45016 18701 45057 18753
rect 44505 18697 45057 18701
rect 42873 18645 42910 18697
rect 42962 18645 43419 18697
rect 43471 18693 45057 18697
rect 43471 18645 43934 18693
rect 42873 18641 43934 18645
rect 43986 18689 45057 18693
rect 43986 18685 44964 18689
rect 43986 18641 44453 18685
rect 42873 18633 44453 18641
rect 44505 18637 44964 18685
rect 45016 18637 45057 18689
rect 44505 18633 45057 18637
rect 42873 18614 45057 18633
rect 42891 18611 45057 18614
rect 43556 18610 43762 18611
rect 43897 18610 44027 18611
rect 44416 18602 44546 18611
rect 44927 18606 45057 18611
rect 39316 18300 39496 18344
rect 39316 18248 39348 18300
rect 39400 18248 39412 18300
rect 39464 18248 39496 18300
rect 39316 18204 39496 18248
rect 45530 18215 46586 18320
rect 45530 18213 45616 18215
rect 46472 18213 46586 18215
rect 39346 17925 39476 18204
rect 39346 17873 39385 17925
rect 39437 17873 39476 17925
rect 39346 17834 39476 17873
rect 39656 17117 39966 17144
rect 44673 17123 44803 17124
rect 45530 17123 45602 18213
rect 42633 17118 45602 17123
rect 39656 17087 39726 17117
rect 39906 17087 39966 17117
rect 39656 17031 39708 17087
rect 39924 17031 39966 17087
rect 39656 17001 39726 17031
rect 39906 17001 39966 17031
rect 39656 16974 39966 17001
rect 42621 17100 45602 17118
rect 42621 17088 42722 17100
rect 42621 17036 42658 17088
rect 42710 17044 42722 17088
rect 42778 17094 45602 17100
rect 42778 17091 44710 17094
rect 42778 17090 44188 17091
rect 42778 17084 43672 17090
rect 42778 17044 43158 17084
rect 42710 17036 43158 17044
rect 42621 17032 43158 17036
rect 43210 17038 43672 17084
rect 43724 17039 44188 17090
rect 44240 17042 44710 17091
rect 44762 17088 45602 17094
rect 44762 17042 45216 17088
rect 44240 17039 45216 17042
rect 43724 17038 45216 17039
rect 43210 17036 45216 17038
rect 45268 17036 45602 17088
rect 43210 17032 45602 17036
rect 42621 17030 45602 17032
rect 42621 17027 44710 17030
rect 42621 17026 44188 17027
rect 42621 17024 43672 17026
rect 42621 16972 42658 17024
rect 42710 17020 43672 17024
rect 42710 16972 42722 17020
rect 42621 16964 42722 16972
rect 42778 16968 43158 17020
rect 43210 16974 43672 17020
rect 43724 16975 44188 17026
rect 44240 16978 44710 17027
rect 44762 17024 45602 17030
rect 44762 16978 45216 17024
rect 44240 16975 45216 16978
rect 43724 16974 45216 16975
rect 43210 16972 45216 16974
rect 45268 16972 45602 17024
rect 43210 16968 45602 16972
rect 42778 16966 45602 16968
rect 42778 16964 44710 16966
rect 42621 16963 44710 16964
rect 42621 16962 44188 16963
rect 42621 16960 43672 16962
rect 39156 16855 39396 16934
rect 42621 16908 42658 16960
rect 42710 16956 43672 16960
rect 42710 16940 43158 16956
rect 42710 16908 42722 16940
rect 42621 16884 42722 16908
rect 42778 16904 43158 16940
rect 43210 16910 43672 16956
rect 43724 16911 44188 16962
rect 44240 16914 44710 16963
rect 44762 16960 45602 16966
rect 44762 16914 45216 16960
rect 44240 16911 45216 16914
rect 43724 16910 45216 16911
rect 43210 16908 45216 16910
rect 45268 16908 45602 16960
rect 43210 16904 45602 16908
rect 42778 16884 45602 16904
rect 42621 16881 45602 16884
rect 46486 16881 46586 18213
rect 42621 16879 45616 16881
rect 46472 16879 46586 16881
rect 42621 16878 46586 16879
rect 42621 16877 42836 16878
rect 42674 16863 42836 16877
rect 43121 16873 43251 16878
rect 45179 16877 45309 16878
rect 39156 16803 39223 16855
rect 39275 16803 39287 16855
rect 39339 16803 39396 16855
rect 45530 16814 46586 16878
rect 39156 15578 39396 16803
rect 40126 15694 40366 16094
rect 40126 15642 40155 15694
rect 40207 15642 40219 15694
rect 40271 15642 40283 15694
rect 40335 15642 40366 15694
rect 40126 15624 40366 15642
rect 38640 15572 40757 15578
rect 38598 15559 40757 15572
rect 38598 15518 40796 15559
rect 38598 15466 38645 15518
rect 38697 15505 40796 15518
rect 38697 15466 39656 15505
rect 38598 15454 39656 15466
rect 38598 15402 38645 15454
rect 38697 15453 39656 15454
rect 39708 15453 40693 15505
rect 40745 15453 40796 15505
rect 38697 15441 40796 15453
rect 38697 15402 39656 15441
rect 38598 15390 39656 15402
rect 38598 15338 38645 15390
rect 38697 15389 39656 15390
rect 39708 15389 40693 15441
rect 40745 15389 40796 15441
rect 38697 15377 40796 15389
rect 38697 15338 39656 15377
rect 38598 15325 39656 15338
rect 39708 15325 40693 15377
rect 40745 15325 40796 15377
rect 35134 15217 36242 15292
rect 38598 15286 40796 15325
rect 38640 15282 40796 15286
rect 39156 15274 39396 15282
rect 39609 15273 39759 15282
rect 40646 15273 40796 15282
rect 35134 14281 35207 15217
rect 36143 14764 36242 15217
rect 36143 14760 41512 14764
rect 36143 14719 41526 14760
rect 36143 14281 41281 14719
rect 35134 14263 41281 14281
rect 41497 14263 41526 14719
rect 35134 14214 41526 14263
rect 35690 14212 41526 14214
rect 39111 13877 39261 13880
rect 40141 13877 40291 13890
rect 38129 13869 40291 13877
rect 38092 13847 40291 13869
rect 38092 13826 39708 13847
rect 38092 13815 39158 13826
rect 38092 13763 38139 13815
rect 38191 13774 39158 13815
rect 39210 13774 39708 13826
rect 38191 13763 39708 13774
rect 38092 13762 39708 13763
rect 38092 13751 39158 13762
rect 38092 13699 38139 13751
rect 38191 13710 39158 13751
rect 39210 13710 39708 13762
rect 38191 13699 39708 13710
rect 38092 13698 39708 13699
rect 38092 13687 39158 13698
rect 38092 13635 38139 13687
rect 38191 13646 39158 13687
rect 39210 13646 39708 13698
rect 38191 13635 39708 13646
rect 38092 13631 39708 13635
rect 39924 13836 40291 13847
rect 39924 13784 40188 13836
rect 40240 13784 40291 13836
rect 39924 13772 40291 13784
rect 39924 13720 40188 13772
rect 40240 13720 40291 13772
rect 39924 13708 40291 13720
rect 39924 13656 40188 13708
rect 40240 13656 40291 13708
rect 39924 13631 40291 13656
rect 38092 13604 40291 13631
rect 38092 13591 40240 13604
rect 38092 13583 38242 13591
rect 37112 13549 37678 13582
rect 37112 13547 37167 13549
rect 37623 13547 37678 13549
rect 37112 13175 37145 13547
rect 37645 13175 37678 13547
rect 41653 13573 41818 13625
rect 41653 13571 41704 13573
rect 41760 13571 41818 13573
rect 38720 13519 38894 13537
rect 38720 13463 38737 13519
rect 38793 13517 38817 13519
rect 38799 13465 38811 13517
rect 38793 13463 38817 13465
rect 38873 13463 38894 13519
rect 38720 13451 38894 13463
rect 37112 13173 37167 13175
rect 37623 13173 37678 13175
rect 37112 13142 37678 13173
rect 41653 13199 41674 13571
rect 41790 13199 41818 13571
rect 41653 13197 41704 13199
rect 41760 13197 41818 13199
rect 41653 13154 41818 13197
rect 37001 11516 41743 11523
rect 37001 11464 37026 11516
rect 37078 11484 41743 11516
rect 37078 11483 41367 11484
rect 37078 11464 37541 11483
rect 37001 11452 37541 11464
rect 37001 11400 37026 11452
rect 37078 11431 37541 11452
rect 37593 11482 38574 11483
rect 37593 11431 38058 11482
rect 37078 11430 38058 11431
rect 38110 11431 38574 11482
rect 38626 11482 41367 11483
rect 38626 11481 39606 11482
rect 38626 11431 39090 11481
rect 38110 11430 39090 11431
rect 37078 11429 39090 11430
rect 39142 11430 39606 11481
rect 39658 11481 40638 11482
rect 39658 11430 40122 11481
rect 39142 11429 40122 11430
rect 40174 11430 40638 11481
rect 40690 11430 41154 11482
rect 41206 11430 41367 11482
rect 40174 11429 41367 11430
rect 37078 11428 41367 11429
rect 41423 11428 41447 11484
rect 41503 11482 41743 11484
rect 41503 11430 41670 11482
rect 41722 11430 41743 11482
rect 41503 11428 41743 11430
rect 37078 11400 41743 11428
rect 37001 11390 41743 11400
rect 36736 11239 41996 11251
rect 36736 11238 39349 11239
rect 36736 11236 37284 11238
rect 36736 11184 36768 11236
rect 36820 11186 37284 11236
rect 37336 11186 37800 11238
rect 37852 11237 38832 11238
rect 37852 11186 38316 11237
rect 36820 11185 38316 11186
rect 38368 11186 38832 11237
rect 38884 11187 39349 11238
rect 39401 11238 41996 11239
rect 39401 11237 40896 11238
rect 39401 11236 40379 11237
rect 39401 11206 39864 11236
rect 39401 11187 39560 11206
rect 38884 11186 39560 11187
rect 38368 11185 39560 11186
rect 36820 11184 39560 11185
rect 36736 11175 39560 11184
rect 36736 11174 39349 11175
rect 36736 11172 37284 11174
rect 36736 11120 36768 11172
rect 36820 11122 37284 11172
rect 37336 11122 37800 11174
rect 37852 11173 38832 11174
rect 37852 11122 38316 11173
rect 36820 11121 38316 11122
rect 38368 11122 38832 11173
rect 38884 11123 39349 11174
rect 39401 11150 39560 11175
rect 39616 11150 39640 11206
rect 39696 11184 39864 11206
rect 39916 11185 40379 11236
rect 40431 11186 40896 11237
rect 40948 11237 41996 11238
rect 40948 11186 41412 11237
rect 40431 11185 41412 11186
rect 41464 11185 41928 11237
rect 41980 11185 41996 11237
rect 39916 11184 41996 11185
rect 39696 11174 41996 11184
rect 39696 11173 40896 11174
rect 39696 11172 40379 11173
rect 39696 11150 39864 11172
rect 39401 11123 39864 11150
rect 38884 11122 39864 11123
rect 38368 11121 39864 11122
rect 36820 11120 39864 11121
rect 39916 11121 40379 11172
rect 40431 11122 40896 11173
rect 40948 11173 41996 11174
rect 40948 11122 41412 11173
rect 40431 11121 41412 11122
rect 41464 11121 41928 11173
rect 41980 11121 41996 11173
rect 39916 11120 41996 11121
rect 36736 11109 41996 11120
rect 38504 10228 40667 10245
rect 38504 10176 38527 10228
rect 38579 10227 40667 10228
rect 38579 10225 39559 10227
rect 38579 10197 39043 10225
rect 38579 10176 38742 10197
rect 38504 10164 38742 10176
rect 38504 10112 38527 10164
rect 38579 10141 38742 10164
rect 38798 10141 38822 10197
rect 38878 10173 39043 10197
rect 39095 10175 39559 10225
rect 39611 10226 40667 10227
rect 39611 10225 40590 10226
rect 39611 10175 40076 10225
rect 39095 10173 40076 10175
rect 40128 10174 40590 10225
rect 40642 10174 40667 10226
rect 40128 10173 40667 10174
rect 38878 10163 40667 10173
rect 38878 10161 39559 10163
rect 38878 10141 39043 10161
rect 38579 10112 39043 10141
rect 38504 10109 39043 10112
rect 39095 10111 39559 10161
rect 39611 10162 40667 10163
rect 39611 10161 40590 10162
rect 39611 10111 40076 10161
rect 39095 10109 40076 10111
rect 40128 10110 40590 10161
rect 40642 10110 40667 10162
rect 40128 10109 40667 10110
rect 38504 10093 40667 10109
rect 38257 9888 40918 9914
rect 38257 9878 38563 9888
rect 38257 9826 38270 9878
rect 38322 9832 38563 9878
rect 38619 9879 40918 9888
rect 38619 9877 39300 9879
rect 38619 9832 38787 9877
rect 38322 9826 38787 9832
rect 38257 9825 38787 9826
rect 38839 9827 39300 9877
rect 39352 9878 40850 9879
rect 39352 9827 39818 9878
rect 38839 9826 39818 9827
rect 39870 9826 40335 9878
rect 40387 9827 40850 9878
rect 40902 9827 40918 9879
rect 40387 9826 40918 9827
rect 38839 9825 40918 9826
rect 38257 9815 40918 9825
rect 38257 9814 39300 9815
rect 38257 9762 38270 9814
rect 38322 9813 39300 9814
rect 38322 9808 38787 9813
rect 38322 9762 38563 9808
rect 38257 9752 38563 9762
rect 38619 9761 38787 9808
rect 38839 9763 39300 9813
rect 39352 9814 40850 9815
rect 39352 9763 39818 9814
rect 38839 9762 39818 9763
rect 39870 9762 40335 9814
rect 40387 9763 40850 9814
rect 40902 9763 40918 9815
rect 40387 9762 40918 9763
rect 38839 9761 40918 9762
rect 38619 9752 40918 9761
rect 38257 9729 40918 9752
rect 43358 9815 44648 9970
rect 43358 9800 43495 9815
rect 43358 7824 43469 9800
rect 43358 7779 43495 7824
rect 44507 7779 44648 9815
rect 43358 7672 44648 7779
rect 38275 7548 42010 7561
rect 38275 7526 41930 7548
rect 38275 7515 38562 7526
rect 38275 7463 38319 7515
rect 38371 7470 38562 7515
rect 38618 7514 41930 7526
rect 38618 7470 41417 7514
rect 38371 7463 41417 7470
rect 38275 7462 41417 7463
rect 41469 7496 41930 7514
rect 41982 7496 42010 7548
rect 41469 7484 42010 7496
rect 41469 7462 41930 7484
rect 38275 7451 41930 7462
rect 38275 7399 38319 7451
rect 38371 7450 41930 7451
rect 38371 7446 41417 7450
rect 38371 7399 38562 7446
rect 38275 7390 38562 7399
rect 38618 7398 41417 7446
rect 41469 7432 41930 7450
rect 41982 7432 42010 7484
rect 41469 7420 42010 7432
rect 41469 7398 41930 7420
rect 38618 7390 41930 7398
rect 38275 7368 41930 7390
rect 41982 7368 42010 7420
rect 38275 7356 42010 7368
rect 38802 7112 40994 7125
rect 38802 7060 38835 7112
rect 38887 7111 40994 7112
rect 38887 7110 40383 7111
rect 38887 7060 39351 7110
rect 38802 7058 39351 7060
rect 39403 7086 40383 7110
rect 39403 7058 39561 7086
rect 38802 7048 39561 7058
rect 38802 6996 38835 7048
rect 38887 7046 39561 7048
rect 38887 6996 39351 7046
rect 38802 6994 39351 6996
rect 39403 6994 39561 7046
rect 38802 6984 39561 6994
rect 38802 6932 38835 6984
rect 38887 6982 39561 6984
rect 38887 6932 39351 6982
rect 38802 6930 39351 6932
rect 39403 6950 39561 6982
rect 39697 7078 40383 7086
rect 39697 7026 39866 7078
rect 39918 7059 40383 7078
rect 40435 7109 40994 7111
rect 40435 7059 40898 7109
rect 39918 7057 40898 7059
rect 40950 7057 40994 7109
rect 39918 7047 40994 7057
rect 39918 7026 40383 7047
rect 39697 7014 40383 7026
rect 39697 6962 39866 7014
rect 39918 6995 40383 7014
rect 40435 7045 40994 7047
rect 40435 6995 40898 7045
rect 39918 6993 40898 6995
rect 40950 6993 40994 7045
rect 39918 6983 40994 6993
rect 39918 6962 40383 6983
rect 39697 6950 40383 6962
rect 39403 6931 40383 6950
rect 40435 6981 40994 6983
rect 40435 6931 40898 6981
rect 39403 6930 40898 6931
rect 38802 6929 40898 6930
rect 40950 6929 40994 6981
rect 38802 6918 40994 6929
rect 37595 6638 42208 6651
rect 37595 6636 38060 6638
rect 37595 6584 37612 6636
rect 37664 6586 38060 6636
rect 38112 6637 42208 6638
rect 38112 6586 38577 6637
rect 37664 6585 38577 6586
rect 38629 6636 39607 6637
rect 38629 6585 39093 6636
rect 37664 6584 39093 6585
rect 39145 6585 39607 6636
rect 39659 6636 40640 6637
rect 39659 6585 40125 6636
rect 39145 6584 40125 6585
rect 40177 6585 40640 6636
rect 40692 6585 41157 6637
rect 41209 6585 41673 6637
rect 41725 6635 42208 6637
rect 41725 6585 42127 6635
rect 40177 6584 42127 6585
rect 37595 6583 42127 6584
rect 42179 6583 42208 6635
rect 37595 6574 42208 6583
rect 37595 6572 38060 6574
rect 37595 6520 37612 6572
rect 37664 6522 38060 6572
rect 38112 6573 42208 6574
rect 38112 6522 38577 6573
rect 37664 6521 38577 6522
rect 38629 6572 39607 6573
rect 38629 6521 39093 6572
rect 37664 6520 39093 6521
rect 39145 6521 39607 6572
rect 39659 6572 40640 6573
rect 39659 6521 40125 6572
rect 39145 6520 40125 6521
rect 40177 6521 40640 6572
rect 40692 6521 41157 6573
rect 41209 6521 41673 6573
rect 41725 6571 42208 6573
rect 41725 6521 42127 6571
rect 40177 6520 42127 6521
rect 37595 6519 42127 6520
rect 42179 6519 42208 6571
rect 37595 6510 42208 6519
rect 37595 6508 38060 6510
rect 37595 6456 37612 6508
rect 37664 6458 38060 6508
rect 38112 6509 42208 6510
rect 38112 6458 38577 6509
rect 37664 6457 38577 6458
rect 38629 6508 39607 6509
rect 38629 6457 39093 6508
rect 37664 6456 39093 6457
rect 39145 6457 39607 6508
rect 39659 6508 40640 6509
rect 39659 6457 40125 6508
rect 39145 6456 40125 6457
rect 40177 6457 40640 6508
rect 40692 6457 41157 6509
rect 41209 6457 41673 6509
rect 41725 6507 42208 6509
rect 41725 6457 42127 6507
rect 40177 6456 42127 6457
rect 37595 6455 42127 6456
rect 42179 6455 42208 6507
rect 37595 6443 42208 6455
rect 41739 6442 42208 6443
rect 32436 2922 32541 3678
rect 33553 2922 33698 3678
rect 32436 2811 33698 2922
rect 49198 3634 50460 22128
rect 49198 2942 49314 3634
rect 50326 2942 50460 3634
rect 49198 2814 50460 2942
rect 30216 758 30400 1514
rect 31284 758 31478 1514
rect 30216 644 31478 758
rect 51356 1493 52618 23957
rect 53360 18574 55010 19136
rect 53360 16518 53650 18574
rect 54506 16518 55010 18574
rect 53360 16110 55010 16518
rect 53214 10282 55944 10672
rect 53214 7186 53542 10282
rect 55278 7186 55944 10282
rect 53214 6898 55944 7186
rect 51356 801 51487 1493
rect 52435 801 52618 1493
rect 51356 649 52618 801
rect 8038 -1044 8106 -96
rect 8990 -1044 9059 -96
rect 8038 -1082 9059 -1044
rect 12750 -172 22754 -16
rect 12750 -992 12843 -172
rect 22623 -534 22754 -172
rect 22623 -992 22752 -534
rect 12750 -1080 22752 -992
<< via2 >>
rect -10189 24654 -9253 25430
rect -115 24520 821 25216
rect -4268 22182 -3572 22200
rect -4268 21362 -4266 22182
rect -4266 21362 -3574 22182
rect -3574 21362 -3572 22182
rect -4268 21344 -3572 21362
rect -4055 18308 -3839 18444
rect -5884 16281 -5866 16337
rect -5866 16281 -5828 16337
rect -5804 16281 -5748 16337
rect -5724 16281 -5686 16337
rect -5686 16281 -5668 16337
rect -2870 16294 -2814 16350
rect -2870 16214 -2814 16270
rect -2870 16134 -2814 16190
rect 45 16183 181 16319
rect -4224 15042 -4214 15178
rect -4214 15042 -4098 15178
rect -4098 15042 -4088 15178
rect -5884 12881 -5668 13097
rect -3888 12821 -3832 12823
rect -6855 12767 -6799 12769
rect -6775 12767 -6719 12769
rect -6855 12715 -6845 12767
rect -6845 12715 -6799 12767
rect -6775 12715 -6729 12767
rect -6729 12715 -6719 12767
rect -6855 12713 -6799 12715
rect -6775 12713 -6719 12715
rect -5333 12626 -4797 12644
rect -5333 12446 -5315 12626
rect -5315 12446 -4815 12626
rect -4815 12446 -4797 12626
rect -5333 12428 -4797 12446
rect -3888 12767 -3832 12821
rect -3888 12687 -3832 12743
rect -3888 12607 -3832 12663
rect -3888 12527 -3832 12583
rect -3888 12449 -3832 12503
rect -3888 12447 -3832 12449
rect -4225 10678 -4169 10734
rect -4145 10678 -4089 10734
rect -9962 9942 -9426 10478
rect -6032 10400 -5976 10456
rect -5952 10400 -5896 10456
rect -6850 9391 -6794 9447
rect -6770 9391 -6714 9447
rect -7029 9082 -6973 9138
rect -7029 9002 -6973 9058
rect -7030 6720 -6974 6776
rect -7030 6640 -6974 6696
rect -6031 6200 -5895 6336
rect 27929 16262 27939 16798
rect 27939 16262 28055 16798
rect 28055 16262 28065 16798
rect 29243 15215 29379 15217
rect 29243 14843 29253 15215
rect 29253 14843 29369 15215
rect 29369 14843 29379 15215
rect 29243 14841 29379 14843
rect 27809 13803 28105 14099
rect 13282 10561 13578 10857
rect 13268 9054 13564 9350
rect 17545 11376 17921 11462
rect 17545 11326 17626 11376
rect 17626 11326 17678 11376
rect 17678 11326 17921 11376
rect 21127 9044 21137 9340
rect 21137 9044 21253 9340
rect 21253 9044 21263 9340
rect 17726 8340 18182 8636
rect 26212 7485 26222 8421
rect 26222 7485 26338 8421
rect 26338 7485 26348 8421
rect 41324 22932 42020 22950
rect 41324 22112 41326 22932
rect 41326 22112 42018 22932
rect 42018 22112 42020 22932
rect 41324 22094 42020 22112
rect 41537 19058 41753 19194
rect 45616 18213 46472 18215
rect 39708 17031 39726 17087
rect 39726 17031 39764 17087
rect 39788 17031 39844 17087
rect 39868 17031 39906 17087
rect 39906 17031 39924 17087
rect 42722 17044 42778 17100
rect 42722 16964 42778 17020
rect 42722 16884 42778 16940
rect 45616 16881 46472 18213
rect 45616 16879 46472 16881
rect 35207 14281 36143 15217
rect 41281 14263 41497 14719
rect 39708 13631 39924 13847
rect 37167 13547 37623 13549
rect 37167 13175 37623 13547
rect 41704 13571 41760 13573
rect 38737 13517 38793 13519
rect 38817 13517 38873 13519
rect 38737 13465 38747 13517
rect 38747 13465 38793 13517
rect 38817 13465 38863 13517
rect 38863 13465 38873 13517
rect 38737 13463 38793 13465
rect 38817 13463 38873 13465
rect 37167 13173 37623 13175
rect 41704 13517 41760 13571
rect 41704 13437 41760 13493
rect 41704 13357 41760 13413
rect 41704 13277 41760 13333
rect 41704 13199 41760 13253
rect 41704 13197 41760 13199
rect 41367 11428 41423 11484
rect 41447 11428 41503 11484
rect 39560 11150 39616 11206
rect 39640 11150 39696 11206
rect 38742 10141 38798 10197
rect 38822 10141 38878 10197
rect 38563 9832 38619 9888
rect 38563 9752 38619 9808
rect 43469 7824 43495 9800
rect 43495 7824 44485 9800
rect 38562 7470 38618 7526
rect 38562 7390 38618 7446
rect 39561 6950 39697 7086
rect 53650 16518 54506 18574
rect 53542 7186 55278 10282
<< metal3 >>
rect -10354 25430 -8968 25616
rect -10354 24654 -10189 25430
rect -9253 24654 -8968 25430
rect -10354 24520 -8968 24654
rect -268 25356 966 25380
rect -268 25216 970 25356
rect -268 24520 -115 25216
rect 821 24520 970 25216
rect -10050 10478 -9270 24520
rect -268 24374 970 24520
rect -268 24366 966 24374
rect -4350 22200 -3490 22289
rect -4350 22164 -4268 22200
rect -3572 22164 -3490 22200
rect -4350 21380 -4272 22164
rect -3568 21380 -3490 22164
rect -4350 21344 -4268 21380
rect -3572 21344 -3490 21380
rect -4350 21265 -3490 21344
rect -4092 18448 -3798 18499
rect -4092 18304 -4059 18448
rect -3835 18304 -3798 18448
rect -4092 18253 -3798 18304
rect -5936 16337 -5626 16394
rect 14 16377 674 24366
rect 41242 22950 42102 23039
rect 41242 22914 41324 22950
rect 42020 22914 42102 22950
rect 41242 22130 41320 22914
rect 42024 22130 42102 22914
rect 41242 22094 41324 22130
rect 42020 22094 42102 22130
rect 41242 22015 42102 22094
rect 41500 19198 41794 19249
rect 41500 19054 41533 19198
rect 41757 19054 41794 19198
rect 41500 19003 41794 19054
rect 53360 18574 55010 19136
rect 53360 18316 53650 18574
rect 45538 18215 53650 18316
rect 39656 17087 39966 17144
rect 39656 17031 39708 17087
rect 39764 17031 39788 17087
rect 39844 17031 39868 17087
rect 39924 17031 39966 17087
rect 42674 17100 42836 17123
rect 42674 17044 42722 17100
rect 42778 17044 42836 17100
rect 42674 17042 42836 17044
rect -5936 16281 -5884 16337
rect -5828 16281 -5804 16337
rect -5748 16281 -5724 16337
rect -5668 16281 -5626 16337
rect -2918 16350 -2756 16373
rect -2918 16294 -2870 16350
rect -2814 16294 -2756 16350
rect -2918 16292 -2756 16294
rect -5936 13097 -5626 16281
rect -5936 12881 -5884 13097
rect -5668 12881 -5626 13097
rect -5936 12844 -5626 12881
rect -4245 16270 -2756 16292
rect -4245 16214 -2870 16270
rect -2814 16214 -2756 16270
rect -4245 16190 -2756 16214
rect -4245 16134 -2870 16190
rect -2814 16134 -2756 16190
rect -4245 16113 -2756 16134
rect -15 16319 674 16377
rect -15 16183 45 16319
rect 181 16183 674 16319
rect -15 16127 674 16183
rect -4245 15178 -4066 16113
rect -13 16070 674 16127
rect 27888 16798 28098 16828
rect 27888 16262 27929 16798
rect 28065 16262 28098 16798
rect 27888 16222 28098 16262
rect -13 15718 242 16070
rect -4245 15042 -4224 15178
rect -4088 15081 -4066 15178
rect -3106 15698 1894 15718
rect -3106 15634 -3078 15698
rect -3014 15634 -2998 15698
rect -2934 15634 -2918 15698
rect -2854 15634 -2838 15698
rect -2774 15634 -2758 15698
rect -2694 15634 -2678 15698
rect -2614 15634 -2598 15698
rect -2534 15634 -2518 15698
rect -2454 15634 -2438 15698
rect -2374 15634 -2358 15698
rect -2294 15634 -2278 15698
rect -2214 15634 -2198 15698
rect -2134 15634 -2118 15698
rect -2054 15634 -2038 15698
rect -1974 15634 -1958 15698
rect -1894 15634 -1878 15698
rect -1814 15634 -1798 15698
rect -1734 15634 -1718 15698
rect -1654 15634 -1638 15698
rect -1574 15634 -1558 15698
rect -1494 15634 -1478 15698
rect -1414 15634 -1398 15698
rect -1334 15634 -1318 15698
rect -1254 15634 -1238 15698
rect -1174 15634 -1158 15698
rect -1094 15634 -1078 15698
rect -1014 15634 -998 15698
rect -934 15634 -918 15698
rect -854 15634 -838 15698
rect -774 15634 -758 15698
rect -694 15634 -678 15698
rect -614 15634 -598 15698
rect -534 15634 -518 15698
rect -454 15634 -438 15698
rect -374 15634 -358 15698
rect -294 15634 -278 15698
rect -214 15634 -198 15698
rect -134 15634 -118 15698
rect -54 15634 -38 15698
rect 26 15634 42 15698
rect 106 15634 122 15698
rect 186 15634 202 15698
rect 266 15634 282 15698
rect 346 15634 362 15698
rect 426 15634 442 15698
rect 506 15634 522 15698
rect 586 15634 602 15698
rect 666 15634 682 15698
rect 746 15634 762 15698
rect 826 15634 842 15698
rect 906 15634 922 15698
rect 986 15634 1002 15698
rect 1066 15634 1082 15698
rect 1146 15634 1162 15698
rect 1226 15634 1242 15698
rect 1306 15634 1322 15698
rect 1386 15634 1402 15698
rect 1466 15634 1482 15698
rect 1546 15634 1562 15698
rect 1626 15634 1642 15698
rect 1706 15634 1722 15698
rect 1786 15634 1802 15698
rect 1866 15634 1894 15698
rect -4088 15042 -4068 15081
rect -10050 9942 -9962 10478
rect -9426 9942 -9270 10478
rect -10050 9880 -9270 9942
rect -6870 12769 -6695 12806
rect -6870 12713 -6855 12769
rect -6799 12713 -6775 12769
rect -6719 12713 -6695 12769
rect -6870 9447 -6695 12713
rect -5381 12644 -4755 12675
rect -5381 12428 -5333 12644
rect -4797 12428 -4755 12644
rect -6870 9391 -6850 9447
rect -6794 9391 -6770 9447
rect -6714 9391 -6695 9447
rect -6870 9343 -6695 9391
rect -6051 10456 -5873 10501
rect -6051 10400 -6032 10456
rect -5976 10400 -5952 10456
rect -5896 10400 -5873 10456
rect -7063 9138 -6938 9164
rect -7063 9082 -7029 9138
rect -6973 9082 -6938 9138
rect -7063 9058 -6938 9082
rect -7063 9002 -7029 9058
rect -6973 9002 -6938 9058
rect -7063 6776 -6938 9002
rect -7063 6720 -7030 6776
rect -6974 6720 -6938 6776
rect -7063 6696 -6938 6720
rect -7063 6640 -7030 6696
rect -6974 6640 -6938 6696
rect -7063 6606 -6938 6640
rect -6051 6336 -5873 10400
rect -5381 9940 -4755 12428
rect -4245 12269 -4068 15042
rect -3939 12827 -3774 12875
rect -3939 12763 -3892 12827
rect -3828 12763 -3774 12827
rect -3939 12747 -3774 12763
rect -3939 12683 -3892 12747
rect -3828 12683 -3774 12747
rect -3939 12667 -3774 12683
rect -3939 12603 -3892 12667
rect -3828 12603 -3774 12667
rect -3939 12587 -3774 12603
rect -3939 12523 -3892 12587
rect -3828 12523 -3774 12587
rect -3939 12507 -3774 12523
rect -3939 12443 -3892 12507
rect -3828 12443 -3774 12507
rect -3939 12404 -3774 12443
rect -4245 10734 -4066 12269
rect -4245 10678 -4225 10734
rect -4169 10678 -4145 10734
rect -4089 10678 -4066 10734
rect -4245 10640 -4066 10678
rect -3106 10619 1894 15634
rect 27888 14686 28096 16222
rect 29188 15217 36230 15292
rect 29188 14841 29243 15217
rect 29379 14841 35207 15217
rect 29188 14740 35207 14841
rect 26178 14478 28096 14686
rect 17510 11462 17962 11498
rect 17510 11326 17545 11462
rect 17921 11326 17962 11462
rect 17510 11290 17962 11326
rect 13198 10938 13662 10942
rect 17618 10938 17958 11290
rect 13198 10857 17962 10938
rect 13198 10561 13282 10857
rect 13578 10561 17962 10857
rect 13198 10496 17962 10561
rect -5381 9923 -1248 9940
rect -5381 9314 -1215 9923
rect -1937 8856 -1215 9314
rect 13194 9398 13644 9424
rect 13194 9350 21302 9398
rect 13194 9054 13268 9350
rect 13564 9340 21302 9350
rect 13564 9054 21127 9340
rect 13194 9044 21127 9054
rect 21263 9044 21302 9340
rect 13194 8994 21302 9044
rect 13194 8988 13644 8994
rect -1937 8636 18226 8856
rect -1937 8340 17726 8636
rect 18182 8340 18226 8636
rect -1937 8134 18226 8340
rect 26178 8421 26386 14478
rect 35134 14281 35207 14740
rect 36143 14281 36230 15217
rect 35134 14214 36230 14281
rect 27750 14099 34680 14168
rect 27750 13803 27809 14099
rect 28105 13803 34680 14099
rect 27750 13728 34680 13803
rect 34240 13582 34680 13728
rect 39656 13847 39966 17031
rect 41347 17020 42836 17042
rect 41347 16964 42722 17020
rect 42778 16964 42836 17020
rect 41347 16940 42836 16964
rect 41347 16884 42722 16940
rect 42778 16884 42836 16940
rect 41347 16863 42836 16884
rect 45538 16879 45616 18215
rect 46472 16879 53650 18215
rect 41347 15831 41526 16863
rect 45538 16792 53650 16879
rect 45579 16468 45834 16792
rect 53360 16518 53650 16792
rect 54506 16518 55010 18574
rect 42486 16448 47486 16468
rect 42486 16384 42514 16448
rect 42578 16384 42594 16448
rect 42658 16384 42674 16448
rect 42738 16384 42754 16448
rect 42818 16384 42834 16448
rect 42898 16384 42914 16448
rect 42978 16384 42994 16448
rect 43058 16384 43074 16448
rect 43138 16384 43154 16448
rect 43218 16384 43234 16448
rect 43298 16384 43314 16448
rect 43378 16384 43394 16448
rect 43458 16384 43474 16448
rect 43538 16384 43554 16448
rect 43618 16384 43634 16448
rect 43698 16384 43714 16448
rect 43778 16384 43794 16448
rect 43858 16384 43874 16448
rect 43938 16384 43954 16448
rect 44018 16384 44034 16448
rect 44098 16384 44114 16448
rect 44178 16384 44194 16448
rect 44258 16384 44274 16448
rect 44338 16384 44354 16448
rect 44418 16384 44434 16448
rect 44498 16384 44514 16448
rect 44578 16384 44594 16448
rect 44658 16384 44674 16448
rect 44738 16384 44754 16448
rect 44818 16384 44834 16448
rect 44898 16384 44914 16448
rect 44978 16384 44994 16448
rect 45058 16384 45074 16448
rect 45138 16384 45154 16448
rect 45218 16384 45234 16448
rect 45298 16384 45314 16448
rect 45378 16384 45394 16448
rect 45458 16384 45474 16448
rect 45538 16384 45554 16448
rect 45618 16384 45634 16448
rect 45698 16384 45714 16448
rect 45778 16384 45794 16448
rect 45858 16384 45874 16448
rect 45938 16384 45954 16448
rect 46018 16384 46034 16448
rect 46098 16384 46114 16448
rect 46178 16384 46194 16448
rect 46258 16384 46274 16448
rect 46338 16384 46354 16448
rect 46418 16384 46434 16448
rect 46498 16384 46514 16448
rect 46578 16384 46594 16448
rect 46658 16384 46674 16448
rect 46738 16384 46754 16448
rect 46818 16384 46834 16448
rect 46898 16384 46914 16448
rect 46978 16384 46994 16448
rect 47058 16384 47074 16448
rect 47138 16384 47154 16448
rect 47218 16384 47234 16448
rect 47298 16384 47314 16448
rect 47378 16384 47394 16448
rect 47458 16384 47486 16448
rect 41347 14764 41524 15831
rect 41246 14719 41526 14764
rect 41246 14263 41281 14719
rect 41497 14263 41526 14719
rect 41246 14212 41526 14263
rect 39656 13631 39708 13847
rect 39924 13631 39966 13847
rect 39656 13594 39966 13631
rect 34240 13549 37678 13582
rect 34240 13173 37167 13549
rect 37623 13173 37678 13549
rect 34240 13142 37678 13173
rect 38722 13519 38897 13556
rect 38722 13463 38737 13519
rect 38793 13463 38817 13519
rect 38873 13463 38897 13519
rect 38722 10197 38897 13463
rect 41347 13019 41524 14212
rect 41653 13577 41818 13625
rect 41653 13513 41700 13577
rect 41764 13513 41818 13577
rect 41653 13497 41818 13513
rect 41653 13433 41700 13497
rect 41764 13433 41818 13497
rect 41653 13417 41818 13433
rect 41653 13353 41700 13417
rect 41764 13353 41818 13417
rect 41653 13337 41818 13353
rect 41653 13273 41700 13337
rect 41764 13273 41818 13337
rect 41653 13257 41818 13273
rect 41653 13193 41700 13257
rect 41764 13193 41818 13257
rect 41653 13154 41818 13193
rect 41347 11484 41526 13019
rect 41347 11428 41367 11484
rect 41423 11428 41447 11484
rect 41503 11428 41526 11484
rect 41347 11390 41526 11428
rect 42486 11369 47486 16384
rect 53360 16110 55010 16518
rect 38722 10141 38742 10197
rect 38798 10141 38822 10197
rect 38878 10141 38897 10197
rect 38722 10093 38897 10141
rect 39541 11206 39719 11251
rect 39541 11150 39560 11206
rect 39616 11150 39640 11206
rect 39696 11150 39719 11206
rect 26178 7485 26212 8421
rect 26348 7485 26386 8421
rect 26178 7452 26386 7485
rect 38529 9888 38654 9914
rect 38529 9832 38563 9888
rect 38619 9832 38654 9888
rect 38529 9808 38654 9832
rect 38529 9752 38563 9808
rect 38619 9752 38654 9808
rect 38529 7526 38654 9752
rect 38529 7470 38562 7526
rect 38618 7470 38654 7526
rect 38529 7446 38654 7470
rect 38529 7390 38562 7446
rect 38618 7390 38654 7446
rect 38529 7356 38654 7390
rect 39541 7086 39719 11150
rect 53214 10282 55944 10672
rect 53214 9974 53542 10282
rect 43366 9800 53542 9974
rect 43366 7824 43469 9800
rect 44485 7824 53542 9800
rect 43366 7664 53542 7824
rect 39541 6950 39561 7086
rect 39697 6950 39719 7086
rect 39541 6918 39719 6950
rect 53214 7186 53542 7664
rect 55278 7186 55944 10282
rect 53214 6898 55944 7186
rect -6051 6200 -6031 6336
rect -5895 6200 -5873 6336
rect -6051 6168 -5873 6200
<< via3 >>
rect -4272 21380 -4268 22164
rect -4268 21380 -3572 22164
rect -3572 21380 -3568 22164
rect -4059 18444 -3835 18448
rect -4059 18308 -4055 18444
rect -4055 18308 -3839 18444
rect -3839 18308 -3835 18444
rect -4059 18304 -3835 18308
rect 41320 22130 41324 22914
rect 41324 22130 42020 22914
rect 42020 22130 42024 22914
rect 41533 19194 41757 19198
rect 41533 19058 41537 19194
rect 41537 19058 41753 19194
rect 41753 19058 41757 19194
rect 41533 19054 41757 19058
rect -3078 15634 -3014 15698
rect -2998 15634 -2934 15698
rect -2918 15634 -2854 15698
rect -2838 15634 -2774 15698
rect -2758 15634 -2694 15698
rect -2678 15634 -2614 15698
rect -2598 15634 -2534 15698
rect -2518 15634 -2454 15698
rect -2438 15634 -2374 15698
rect -2358 15634 -2294 15698
rect -2278 15634 -2214 15698
rect -2198 15634 -2134 15698
rect -2118 15634 -2054 15698
rect -2038 15634 -1974 15698
rect -1958 15634 -1894 15698
rect -1878 15634 -1814 15698
rect -1798 15634 -1734 15698
rect -1718 15634 -1654 15698
rect -1638 15634 -1574 15698
rect -1558 15634 -1494 15698
rect -1478 15634 -1414 15698
rect -1398 15634 -1334 15698
rect -1318 15634 -1254 15698
rect -1238 15634 -1174 15698
rect -1158 15634 -1094 15698
rect -1078 15634 -1014 15698
rect -998 15634 -934 15698
rect -918 15634 -854 15698
rect -838 15634 -774 15698
rect -758 15634 -694 15698
rect -678 15634 -614 15698
rect -598 15634 -534 15698
rect -518 15634 -454 15698
rect -438 15634 -374 15698
rect -358 15634 -294 15698
rect -278 15634 -214 15698
rect -198 15634 -134 15698
rect -118 15634 -54 15698
rect -38 15634 26 15698
rect 42 15634 106 15698
rect 122 15634 186 15698
rect 202 15634 266 15698
rect 282 15634 346 15698
rect 362 15634 426 15698
rect 442 15634 506 15698
rect 522 15634 586 15698
rect 602 15634 666 15698
rect 682 15634 746 15698
rect 762 15634 826 15698
rect 842 15634 906 15698
rect 922 15634 986 15698
rect 1002 15634 1066 15698
rect 1082 15634 1146 15698
rect 1162 15634 1226 15698
rect 1242 15634 1306 15698
rect 1322 15634 1386 15698
rect 1402 15634 1466 15698
rect 1482 15634 1546 15698
rect 1562 15634 1626 15698
rect 1642 15634 1706 15698
rect 1722 15634 1786 15698
rect 1802 15634 1866 15698
rect -3892 12823 -3828 12827
rect -3892 12767 -3888 12823
rect -3888 12767 -3832 12823
rect -3832 12767 -3828 12823
rect -3892 12763 -3828 12767
rect -3892 12743 -3828 12747
rect -3892 12687 -3888 12743
rect -3888 12687 -3832 12743
rect -3832 12687 -3828 12743
rect -3892 12683 -3828 12687
rect -3892 12663 -3828 12667
rect -3892 12607 -3888 12663
rect -3888 12607 -3832 12663
rect -3832 12607 -3828 12663
rect -3892 12603 -3828 12607
rect -3892 12583 -3828 12587
rect -3892 12527 -3888 12583
rect -3888 12527 -3832 12583
rect -3832 12527 -3828 12583
rect -3892 12523 -3828 12527
rect -3892 12503 -3828 12507
rect -3892 12447 -3888 12503
rect -3888 12447 -3832 12503
rect -3832 12447 -3828 12503
rect -3892 12443 -3828 12447
rect 42514 16384 42578 16448
rect 42594 16384 42658 16448
rect 42674 16384 42738 16448
rect 42754 16384 42818 16448
rect 42834 16384 42898 16448
rect 42914 16384 42978 16448
rect 42994 16384 43058 16448
rect 43074 16384 43138 16448
rect 43154 16384 43218 16448
rect 43234 16384 43298 16448
rect 43314 16384 43378 16448
rect 43394 16384 43458 16448
rect 43474 16384 43538 16448
rect 43554 16384 43618 16448
rect 43634 16384 43698 16448
rect 43714 16384 43778 16448
rect 43794 16384 43858 16448
rect 43874 16384 43938 16448
rect 43954 16384 44018 16448
rect 44034 16384 44098 16448
rect 44114 16384 44178 16448
rect 44194 16384 44258 16448
rect 44274 16384 44338 16448
rect 44354 16384 44418 16448
rect 44434 16384 44498 16448
rect 44514 16384 44578 16448
rect 44594 16384 44658 16448
rect 44674 16384 44738 16448
rect 44754 16384 44818 16448
rect 44834 16384 44898 16448
rect 44914 16384 44978 16448
rect 44994 16384 45058 16448
rect 45074 16384 45138 16448
rect 45154 16384 45218 16448
rect 45234 16384 45298 16448
rect 45314 16384 45378 16448
rect 45394 16384 45458 16448
rect 45474 16384 45538 16448
rect 45554 16384 45618 16448
rect 45634 16384 45698 16448
rect 45714 16384 45778 16448
rect 45794 16384 45858 16448
rect 45874 16384 45938 16448
rect 45954 16384 46018 16448
rect 46034 16384 46098 16448
rect 46114 16384 46178 16448
rect 46194 16384 46258 16448
rect 46274 16384 46338 16448
rect 46354 16384 46418 16448
rect 46434 16384 46498 16448
rect 46514 16384 46578 16448
rect 46594 16384 46658 16448
rect 46674 16384 46738 16448
rect 46754 16384 46818 16448
rect 46834 16384 46898 16448
rect 46914 16384 46978 16448
rect 46994 16384 47058 16448
rect 47074 16384 47138 16448
rect 47154 16384 47218 16448
rect 47234 16384 47298 16448
rect 47314 16384 47378 16448
rect 47394 16384 47458 16448
rect 41700 13573 41764 13577
rect 41700 13517 41704 13573
rect 41704 13517 41760 13573
rect 41760 13517 41764 13573
rect 41700 13513 41764 13517
rect 41700 13493 41764 13497
rect 41700 13437 41704 13493
rect 41704 13437 41760 13493
rect 41760 13437 41764 13493
rect 41700 13433 41764 13437
rect 41700 13413 41764 13417
rect 41700 13357 41704 13413
rect 41704 13357 41760 13413
rect 41760 13357 41764 13413
rect 41700 13353 41764 13357
rect 41700 13333 41764 13337
rect 41700 13277 41704 13333
rect 41704 13277 41760 13333
rect 41760 13277 41764 13333
rect 41700 13273 41764 13277
rect 41700 13253 41764 13257
rect 41700 13197 41704 13253
rect 41704 13197 41760 13253
rect 41760 13197 41764 13253
rect 41700 13193 41764 13197
<< mimcap >>
rect 42586 16221 47386 16269
rect -3006 15471 1794 15519
rect -3006 10767 -2958 15471
rect 1746 10767 1794 15471
rect 42586 11517 42634 16221
rect 47338 11517 47386 16221
rect 42586 11469 47386 11517
rect -3006 10719 1794 10767
<< mimcapcontact >>
rect -2958 10767 1746 15471
rect 42634 11517 47338 16221
<< metal4 >>
rect 41502 23039 41792 23040
rect 41242 22914 42102 23039
rect -4090 22289 -3800 22290
rect -4350 22164 -3490 22289
rect -4350 21380 -4272 22164
rect -3568 21380 -3490 22164
rect 41242 22130 41320 22914
rect 42024 22130 42102 22914
rect 41242 22015 42102 22130
rect -4350 21265 -3490 21380
rect -4090 18448 -3800 21265
rect 41502 19198 41792 22015
rect 41502 19054 41533 19198
rect 41757 19054 41792 19198
rect 41502 19007 41792 19054
rect -4090 18304 -4059 18448
rect -3835 18304 -3800 18448
rect -4090 18257 -3800 18304
rect 42498 16448 47474 16464
rect 42498 16384 42514 16448
rect 42578 16384 42594 16448
rect 42658 16384 42674 16448
rect 42738 16384 42754 16448
rect 42818 16384 42834 16448
rect 42898 16384 42914 16448
rect 42978 16384 42994 16448
rect 43058 16384 43074 16448
rect 43138 16384 43154 16448
rect 43218 16384 43234 16448
rect 43298 16384 43314 16448
rect 43378 16384 43394 16448
rect 43458 16384 43474 16448
rect 43538 16384 43554 16448
rect 43618 16384 43634 16448
rect 43698 16384 43714 16448
rect 43778 16384 43794 16448
rect 43858 16384 43874 16448
rect 43938 16384 43954 16448
rect 44018 16384 44034 16448
rect 44098 16384 44114 16448
rect 44178 16384 44194 16448
rect 44258 16384 44274 16448
rect 44338 16384 44354 16448
rect 44418 16384 44434 16448
rect 44498 16384 44514 16448
rect 44578 16384 44594 16448
rect 44658 16384 44674 16448
rect 44738 16384 44754 16448
rect 44818 16384 44834 16448
rect 44898 16384 44914 16448
rect 44978 16384 44994 16448
rect 45058 16384 45074 16448
rect 45138 16384 45154 16448
rect 45218 16384 45234 16448
rect 45298 16384 45314 16448
rect 45378 16384 45394 16448
rect 45458 16384 45474 16448
rect 45538 16384 45554 16448
rect 45618 16384 45634 16448
rect 45698 16384 45714 16448
rect 45778 16384 45794 16448
rect 45858 16384 45874 16448
rect 45938 16384 45954 16448
rect 46018 16384 46034 16448
rect 46098 16384 46114 16448
rect 46178 16384 46194 16448
rect 46258 16384 46274 16448
rect 46338 16384 46354 16448
rect 46418 16384 46434 16448
rect 46498 16384 46514 16448
rect 46578 16384 46594 16448
rect 46658 16384 46674 16448
rect 46738 16384 46754 16448
rect 46818 16384 46834 16448
rect 46898 16384 46914 16448
rect 46978 16384 46994 16448
rect 47058 16384 47074 16448
rect 47138 16384 47154 16448
rect 47218 16384 47234 16448
rect 47298 16384 47314 16448
rect 47378 16384 47394 16448
rect 47458 16384 47474 16448
rect 42498 16368 47474 16384
rect 42625 16221 47347 16230
rect -3094 15698 1882 15714
rect -3094 15634 -3078 15698
rect -3014 15634 -2998 15698
rect -2934 15634 -2918 15698
rect -2854 15634 -2838 15698
rect -2774 15634 -2758 15698
rect -2694 15634 -2678 15698
rect -2614 15634 -2598 15698
rect -2534 15634 -2518 15698
rect -2454 15634 -2438 15698
rect -2374 15634 -2358 15698
rect -2294 15634 -2278 15698
rect -2214 15634 -2198 15698
rect -2134 15634 -2118 15698
rect -2054 15634 -2038 15698
rect -1974 15634 -1958 15698
rect -1894 15634 -1878 15698
rect -1814 15634 -1798 15698
rect -1734 15634 -1718 15698
rect -1654 15634 -1638 15698
rect -1574 15634 -1558 15698
rect -1494 15634 -1478 15698
rect -1414 15634 -1398 15698
rect -1334 15634 -1318 15698
rect -1254 15634 -1238 15698
rect -1174 15634 -1158 15698
rect -1094 15634 -1078 15698
rect -1014 15634 -998 15698
rect -934 15634 -918 15698
rect -854 15634 -838 15698
rect -774 15634 -758 15698
rect -694 15634 -678 15698
rect -614 15634 -598 15698
rect -534 15634 -518 15698
rect -454 15634 -438 15698
rect -374 15634 -358 15698
rect -294 15634 -278 15698
rect -214 15634 -198 15698
rect -134 15634 -118 15698
rect -54 15634 -38 15698
rect 26 15634 42 15698
rect 106 15634 122 15698
rect 186 15634 202 15698
rect 266 15634 282 15698
rect 346 15634 362 15698
rect 426 15634 442 15698
rect 506 15634 522 15698
rect 586 15634 602 15698
rect 666 15634 682 15698
rect 746 15634 762 15698
rect 826 15634 842 15698
rect 906 15634 922 15698
rect 986 15634 1002 15698
rect 1066 15634 1082 15698
rect 1146 15634 1162 15698
rect 1226 15634 1242 15698
rect 1306 15634 1322 15698
rect 1386 15634 1402 15698
rect 1466 15634 1482 15698
rect 1546 15634 1562 15698
rect 1626 15634 1642 15698
rect 1706 15634 1722 15698
rect 1786 15634 1802 15698
rect 1866 15634 1882 15698
rect -3094 15618 1882 15634
rect -2967 15471 1755 15480
rect -3939 12855 -3774 12875
rect -2967 12855 -2958 15471
rect -3939 12827 -2958 12855
rect -3939 12763 -3892 12827
rect -3828 12763 -2958 12827
rect -3939 12747 -2958 12763
rect -3939 12683 -3892 12747
rect -3828 12683 -2958 12747
rect -3939 12667 -2958 12683
rect -3939 12603 -3892 12667
rect -3828 12603 -2958 12667
rect -3939 12587 -2958 12603
rect -3939 12523 -3892 12587
rect -3828 12523 -2958 12587
rect -3939 12507 -2958 12523
rect -3939 12443 -3892 12507
rect -3828 12443 -2958 12507
rect -3939 12404 -2958 12443
rect -2967 10767 -2958 12404
rect 1746 10767 1755 15471
rect 41653 13605 41818 13625
rect 42625 13605 42634 16221
rect 41653 13577 42634 13605
rect 41653 13513 41700 13577
rect 41764 13513 42634 13577
rect 41653 13497 42634 13513
rect 41653 13433 41700 13497
rect 41764 13433 42634 13497
rect 41653 13417 42634 13433
rect 41653 13353 41700 13417
rect 41764 13353 42634 13417
rect 41653 13337 42634 13353
rect 41653 13273 41700 13337
rect 41764 13273 42634 13337
rect 41653 13257 42634 13273
rect 41653 13193 41700 13257
rect 41764 13193 42634 13257
rect 41653 13154 42634 13193
rect 42625 11517 42634 13154
rect 47338 11517 47347 16221
rect 42625 11508 47347 11517
rect -2967 10758 1755 10767
<< labels >>
flabel metal1 s 26368 22558 26368 22558 0 FreeSans 10000 0 0 0 VDD
port 1 nsew
flabel metal1 s 26430 24258 26430 24258 0 FreeSans 10000 0 0 0 VSS
port 2 nsew
flabel metal3 s 45742 16738 45742 16738 0 FreeSans 10000 0 0 0 Vfinal
port 3 nsew
flabel metal1 s 38112 10752 38112 10752 0 FreeSans 10000 0 0 0 IBIAS
port 4 nsew
flabel metal1 s -7552 9972 -7552 9972 0 FreeSans 10000 0 0 0 IBIAS2
port 5 nsew
flabel metal3 s 92 15942 92 15942 0 FreeSans 10000 0 0 0 VBGR1
port 6 nsew
<< end >>
