magic
tech sky130B
magscale 1 2
timestamp 1667543118
<< nwell >>
rect -3138 -3138 3138 3138
<< pwell >>
rect -3266 3180 3266 3266
rect -3266 -3180 -3180 3180
rect 3180 -3180 3266 3180
rect -3266 -3266 3266 -3180
<< psubdiff >>
rect -3240 3206 -3111 3240
rect -3077 3206 -3043 3240
rect -3009 3206 -2975 3240
rect -2941 3206 -2907 3240
rect -2873 3206 -2839 3240
rect -2805 3206 -2771 3240
rect -2737 3206 -2703 3240
rect -2669 3206 -2635 3240
rect -2601 3206 -2567 3240
rect -2533 3206 -2499 3240
rect -2465 3206 -2431 3240
rect -2397 3206 -2363 3240
rect -2329 3206 -2295 3240
rect -2261 3206 -2227 3240
rect -2193 3206 -2159 3240
rect -2125 3206 -2091 3240
rect -2057 3206 -2023 3240
rect -1989 3206 -1955 3240
rect -1921 3206 -1887 3240
rect -1853 3206 -1819 3240
rect -1785 3206 -1751 3240
rect -1717 3206 -1683 3240
rect -1649 3206 -1615 3240
rect -1581 3206 -1547 3240
rect -1513 3206 -1479 3240
rect -1445 3206 -1411 3240
rect -1377 3206 -1343 3240
rect -1309 3206 -1275 3240
rect -1241 3206 -1207 3240
rect -1173 3206 -1139 3240
rect -1105 3206 -1071 3240
rect -1037 3206 -1003 3240
rect -969 3206 -935 3240
rect -901 3206 -867 3240
rect -833 3206 -799 3240
rect -765 3206 -731 3240
rect -697 3206 -663 3240
rect -629 3206 -595 3240
rect -561 3206 -527 3240
rect -493 3206 -459 3240
rect -425 3206 -391 3240
rect -357 3206 -323 3240
rect -289 3206 -255 3240
rect -221 3206 -187 3240
rect -153 3206 -119 3240
rect -85 3206 -51 3240
rect -17 3206 17 3240
rect 51 3206 85 3240
rect 119 3206 153 3240
rect 187 3206 221 3240
rect 255 3206 289 3240
rect 323 3206 357 3240
rect 391 3206 425 3240
rect 459 3206 493 3240
rect 527 3206 561 3240
rect 595 3206 629 3240
rect 663 3206 697 3240
rect 731 3206 765 3240
rect 799 3206 833 3240
rect 867 3206 901 3240
rect 935 3206 969 3240
rect 1003 3206 1037 3240
rect 1071 3206 1105 3240
rect 1139 3206 1173 3240
rect 1207 3206 1241 3240
rect 1275 3206 1309 3240
rect 1343 3206 1377 3240
rect 1411 3206 1445 3240
rect 1479 3206 1513 3240
rect 1547 3206 1581 3240
rect 1615 3206 1649 3240
rect 1683 3206 1717 3240
rect 1751 3206 1785 3240
rect 1819 3206 1853 3240
rect 1887 3206 1921 3240
rect 1955 3206 1989 3240
rect 2023 3206 2057 3240
rect 2091 3206 2125 3240
rect 2159 3206 2193 3240
rect 2227 3206 2261 3240
rect 2295 3206 2329 3240
rect 2363 3206 2397 3240
rect 2431 3206 2465 3240
rect 2499 3206 2533 3240
rect 2567 3206 2601 3240
rect 2635 3206 2669 3240
rect 2703 3206 2737 3240
rect 2771 3206 2805 3240
rect 2839 3206 2873 3240
rect 2907 3206 2941 3240
rect 2975 3206 3009 3240
rect 3043 3206 3077 3240
rect 3111 3206 3240 3240
rect -3240 3111 -3206 3206
rect 3206 3111 3240 3206
rect -3240 3043 -3206 3077
rect -3240 2975 -3206 3009
rect -3240 2907 -3206 2941
rect -3240 2839 -3206 2873
rect -3240 2771 -3206 2805
rect -3240 2703 -3206 2737
rect -3240 2635 -3206 2669
rect -3240 2567 -3206 2601
rect -3240 2499 -3206 2533
rect -3240 2431 -3206 2465
rect -3240 2363 -3206 2397
rect -3240 2295 -3206 2329
rect -3240 2227 -3206 2261
rect -3240 2159 -3206 2193
rect -3240 2091 -3206 2125
rect -3240 2023 -3206 2057
rect -3240 1955 -3206 1989
rect -3240 1887 -3206 1921
rect -3240 1819 -3206 1853
rect -3240 1751 -3206 1785
rect -3240 1683 -3206 1717
rect -3240 1615 -3206 1649
rect -3240 1547 -3206 1581
rect -3240 1479 -3206 1513
rect -3240 1411 -3206 1445
rect -3240 1343 -3206 1377
rect -3240 1275 -3206 1309
rect -3240 1207 -3206 1241
rect -3240 1139 -3206 1173
rect -3240 1071 -3206 1105
rect -3240 1003 -3206 1037
rect -3240 935 -3206 969
rect -3240 867 -3206 901
rect -3240 799 -3206 833
rect -3240 731 -3206 765
rect -3240 663 -3206 697
rect -3240 595 -3206 629
rect -3240 527 -3206 561
rect -3240 459 -3206 493
rect -3240 391 -3206 425
rect -3240 323 -3206 357
rect -3240 255 -3206 289
rect -3240 187 -3206 221
rect -3240 119 -3206 153
rect -3240 51 -3206 85
rect -3240 -17 -3206 17
rect -3240 -85 -3206 -51
rect -3240 -153 -3206 -119
rect -3240 -221 -3206 -187
rect -3240 -289 -3206 -255
rect -3240 -357 -3206 -323
rect -3240 -425 -3206 -391
rect -3240 -493 -3206 -459
rect -3240 -561 -3206 -527
rect -3240 -629 -3206 -595
rect -3240 -697 -3206 -663
rect -3240 -765 -3206 -731
rect -3240 -833 -3206 -799
rect -3240 -901 -3206 -867
rect -3240 -969 -3206 -935
rect -3240 -1037 -3206 -1003
rect -3240 -1105 -3206 -1071
rect -3240 -1173 -3206 -1139
rect -3240 -1241 -3206 -1207
rect -3240 -1309 -3206 -1275
rect -3240 -1377 -3206 -1343
rect -3240 -1445 -3206 -1411
rect -3240 -1513 -3206 -1479
rect -3240 -1581 -3206 -1547
rect -3240 -1649 -3206 -1615
rect -3240 -1717 -3206 -1683
rect -3240 -1785 -3206 -1751
rect -3240 -1853 -3206 -1819
rect -3240 -1921 -3206 -1887
rect -3240 -1989 -3206 -1955
rect -3240 -2057 -3206 -2023
rect -3240 -2125 -3206 -2091
rect -3240 -2193 -3206 -2159
rect -3240 -2261 -3206 -2227
rect -3240 -2329 -3206 -2295
rect -3240 -2397 -3206 -2363
rect -3240 -2465 -3206 -2431
rect -3240 -2533 -3206 -2499
rect -3240 -2601 -3206 -2567
rect -3240 -2669 -3206 -2635
rect -3240 -2737 -3206 -2703
rect -3240 -2805 -3206 -2771
rect -3240 -2873 -3206 -2839
rect -3240 -2941 -3206 -2907
rect -3240 -3009 -3206 -2975
rect -3240 -3077 -3206 -3043
rect 3206 3043 3240 3077
rect 3206 2975 3240 3009
rect 3206 2907 3240 2941
rect 3206 2839 3240 2873
rect 3206 2771 3240 2805
rect 3206 2703 3240 2737
rect 3206 2635 3240 2669
rect 3206 2567 3240 2601
rect 3206 2499 3240 2533
rect 3206 2431 3240 2465
rect 3206 2363 3240 2397
rect 3206 2295 3240 2329
rect 3206 2227 3240 2261
rect 3206 2159 3240 2193
rect 3206 2091 3240 2125
rect 3206 2023 3240 2057
rect 3206 1955 3240 1989
rect 3206 1887 3240 1921
rect 3206 1819 3240 1853
rect 3206 1751 3240 1785
rect 3206 1683 3240 1717
rect 3206 1615 3240 1649
rect 3206 1547 3240 1581
rect 3206 1479 3240 1513
rect 3206 1411 3240 1445
rect 3206 1343 3240 1377
rect 3206 1275 3240 1309
rect 3206 1207 3240 1241
rect 3206 1139 3240 1173
rect 3206 1071 3240 1105
rect 3206 1003 3240 1037
rect 3206 935 3240 969
rect 3206 867 3240 901
rect 3206 799 3240 833
rect 3206 731 3240 765
rect 3206 663 3240 697
rect 3206 595 3240 629
rect 3206 527 3240 561
rect 3206 459 3240 493
rect 3206 391 3240 425
rect 3206 323 3240 357
rect 3206 255 3240 289
rect 3206 187 3240 221
rect 3206 119 3240 153
rect 3206 51 3240 85
rect 3206 -17 3240 17
rect 3206 -85 3240 -51
rect 3206 -153 3240 -119
rect 3206 -221 3240 -187
rect 3206 -289 3240 -255
rect 3206 -357 3240 -323
rect 3206 -425 3240 -391
rect 3206 -493 3240 -459
rect 3206 -561 3240 -527
rect 3206 -629 3240 -595
rect 3206 -697 3240 -663
rect 3206 -765 3240 -731
rect 3206 -833 3240 -799
rect 3206 -901 3240 -867
rect 3206 -969 3240 -935
rect 3206 -1037 3240 -1003
rect 3206 -1105 3240 -1071
rect 3206 -1173 3240 -1139
rect 3206 -1241 3240 -1207
rect 3206 -1309 3240 -1275
rect 3206 -1377 3240 -1343
rect 3206 -1445 3240 -1411
rect 3206 -1513 3240 -1479
rect 3206 -1581 3240 -1547
rect 3206 -1649 3240 -1615
rect 3206 -1717 3240 -1683
rect 3206 -1785 3240 -1751
rect 3206 -1853 3240 -1819
rect 3206 -1921 3240 -1887
rect 3206 -1989 3240 -1955
rect 3206 -2057 3240 -2023
rect 3206 -2125 3240 -2091
rect 3206 -2193 3240 -2159
rect 3206 -2261 3240 -2227
rect 3206 -2329 3240 -2295
rect 3206 -2397 3240 -2363
rect 3206 -2465 3240 -2431
rect 3206 -2533 3240 -2499
rect 3206 -2601 3240 -2567
rect 3206 -2669 3240 -2635
rect 3206 -2737 3240 -2703
rect 3206 -2805 3240 -2771
rect 3206 -2873 3240 -2839
rect 3206 -2941 3240 -2907
rect 3206 -3009 3240 -2975
rect 3206 -3077 3240 -3043
rect -3240 -3206 -3206 -3111
rect 3206 -3206 3240 -3111
rect -3240 -3240 -3111 -3206
rect -3077 -3240 -3043 -3206
rect -3009 -3240 -2975 -3206
rect -2941 -3240 -2907 -3206
rect -2873 -3240 -2839 -3206
rect -2805 -3240 -2771 -3206
rect -2737 -3240 -2703 -3206
rect -2669 -3240 -2635 -3206
rect -2601 -3240 -2567 -3206
rect -2533 -3240 -2499 -3206
rect -2465 -3240 -2431 -3206
rect -2397 -3240 -2363 -3206
rect -2329 -3240 -2295 -3206
rect -2261 -3240 -2227 -3206
rect -2193 -3240 -2159 -3206
rect -2125 -3240 -2091 -3206
rect -2057 -3240 -2023 -3206
rect -1989 -3240 -1955 -3206
rect -1921 -3240 -1887 -3206
rect -1853 -3240 -1819 -3206
rect -1785 -3240 -1751 -3206
rect -1717 -3240 -1683 -3206
rect -1649 -3240 -1615 -3206
rect -1581 -3240 -1547 -3206
rect -1513 -3240 -1479 -3206
rect -1445 -3240 -1411 -3206
rect -1377 -3240 -1343 -3206
rect -1309 -3240 -1275 -3206
rect -1241 -3240 -1207 -3206
rect -1173 -3240 -1139 -3206
rect -1105 -3240 -1071 -3206
rect -1037 -3240 -1003 -3206
rect -969 -3240 -935 -3206
rect -901 -3240 -867 -3206
rect -833 -3240 -799 -3206
rect -765 -3240 -731 -3206
rect -697 -3240 -663 -3206
rect -629 -3240 -595 -3206
rect -561 -3240 -527 -3206
rect -493 -3240 -459 -3206
rect -425 -3240 -391 -3206
rect -357 -3240 -323 -3206
rect -289 -3240 -255 -3206
rect -221 -3240 -187 -3206
rect -153 -3240 -119 -3206
rect -85 -3240 -51 -3206
rect -17 -3240 17 -3206
rect 51 -3240 85 -3206
rect 119 -3240 153 -3206
rect 187 -3240 221 -3206
rect 255 -3240 289 -3206
rect 323 -3240 357 -3206
rect 391 -3240 425 -3206
rect 459 -3240 493 -3206
rect 527 -3240 561 -3206
rect 595 -3240 629 -3206
rect 663 -3240 697 -3206
rect 731 -3240 765 -3206
rect 799 -3240 833 -3206
rect 867 -3240 901 -3206
rect 935 -3240 969 -3206
rect 1003 -3240 1037 -3206
rect 1071 -3240 1105 -3206
rect 1139 -3240 1173 -3206
rect 1207 -3240 1241 -3206
rect 1275 -3240 1309 -3206
rect 1343 -3240 1377 -3206
rect 1411 -3240 1445 -3206
rect 1479 -3240 1513 -3206
rect 1547 -3240 1581 -3206
rect 1615 -3240 1649 -3206
rect 1683 -3240 1717 -3206
rect 1751 -3240 1785 -3206
rect 1819 -3240 1853 -3206
rect 1887 -3240 1921 -3206
rect 1955 -3240 1989 -3206
rect 2023 -3240 2057 -3206
rect 2091 -3240 2125 -3206
rect 2159 -3240 2193 -3206
rect 2227 -3240 2261 -3206
rect 2295 -3240 2329 -3206
rect 2363 -3240 2397 -3206
rect 2431 -3240 2465 -3206
rect 2499 -3240 2533 -3206
rect 2567 -3240 2601 -3206
rect 2635 -3240 2669 -3206
rect 2703 -3240 2737 -3206
rect 2771 -3240 2805 -3206
rect 2839 -3240 2873 -3206
rect 2907 -3240 2941 -3206
rect 2975 -3240 3009 -3206
rect 3043 -3240 3077 -3206
rect 3111 -3240 3240 -3206
<< nsubdiff >>
rect -3102 3068 -2975 3102
rect -2941 3068 -2907 3102
rect -2873 3068 -2839 3102
rect -2805 3068 -2771 3102
rect -2737 3068 -2703 3102
rect -2669 3068 -2635 3102
rect -2601 3068 -2567 3102
rect -2533 3068 -2499 3102
rect -2465 3068 -2431 3102
rect -2397 3068 -2363 3102
rect -2329 3068 -2295 3102
rect -2261 3068 -2227 3102
rect -2193 3068 -2159 3102
rect -2125 3068 -2091 3102
rect -2057 3068 -2023 3102
rect -1989 3068 -1955 3102
rect -1921 3068 -1887 3102
rect -1853 3068 -1819 3102
rect -1785 3068 -1751 3102
rect -1717 3068 -1683 3102
rect -1649 3068 -1615 3102
rect -1581 3068 -1547 3102
rect -1513 3068 -1479 3102
rect -1445 3068 -1411 3102
rect -1377 3068 -1343 3102
rect -1309 3068 -1275 3102
rect -1241 3068 -1207 3102
rect -1173 3068 -1139 3102
rect -1105 3068 -1071 3102
rect -1037 3068 -1003 3102
rect -969 3068 -935 3102
rect -901 3068 -867 3102
rect -833 3068 -799 3102
rect -765 3068 -731 3102
rect -697 3068 -663 3102
rect -629 3068 -595 3102
rect -561 3068 -527 3102
rect -493 3068 -459 3102
rect -425 3068 -391 3102
rect -357 3068 -323 3102
rect -289 3068 -255 3102
rect -221 3068 -187 3102
rect -153 3068 -119 3102
rect -85 3068 -51 3102
rect -17 3068 17 3102
rect 51 3068 85 3102
rect 119 3068 153 3102
rect 187 3068 221 3102
rect 255 3068 289 3102
rect 323 3068 357 3102
rect 391 3068 425 3102
rect 459 3068 493 3102
rect 527 3068 561 3102
rect 595 3068 629 3102
rect 663 3068 697 3102
rect 731 3068 765 3102
rect 799 3068 833 3102
rect 867 3068 901 3102
rect 935 3068 969 3102
rect 1003 3068 1037 3102
rect 1071 3068 1105 3102
rect 1139 3068 1173 3102
rect 1207 3068 1241 3102
rect 1275 3068 1309 3102
rect 1343 3068 1377 3102
rect 1411 3068 1445 3102
rect 1479 3068 1513 3102
rect 1547 3068 1581 3102
rect 1615 3068 1649 3102
rect 1683 3068 1717 3102
rect 1751 3068 1785 3102
rect 1819 3068 1853 3102
rect 1887 3068 1921 3102
rect 1955 3068 1989 3102
rect 2023 3068 2057 3102
rect 2091 3068 2125 3102
rect 2159 3068 2193 3102
rect 2227 3068 2261 3102
rect 2295 3068 2329 3102
rect 2363 3068 2397 3102
rect 2431 3068 2465 3102
rect 2499 3068 2533 3102
rect 2567 3068 2601 3102
rect 2635 3068 2669 3102
rect 2703 3068 2737 3102
rect 2771 3068 2805 3102
rect 2839 3068 2873 3102
rect 2907 3068 2941 3102
rect 2975 3068 3102 3102
rect -3102 2975 -3068 3068
rect -3102 2907 -3068 2941
rect -3102 2839 -3068 2873
rect -3102 2771 -3068 2805
rect -3102 2703 -3068 2737
rect -3102 2635 -3068 2669
rect -3102 2567 -3068 2601
rect -3102 2499 -3068 2533
rect -3102 2431 -3068 2465
rect -3102 2363 -3068 2397
rect -3102 2295 -3068 2329
rect -3102 2227 -3068 2261
rect -3102 2159 -3068 2193
rect -3102 2091 -3068 2125
rect -3102 2023 -3068 2057
rect -3102 1955 -3068 1989
rect -3102 1887 -3068 1921
rect -3102 1819 -3068 1853
rect -3102 1751 -3068 1785
rect -3102 1683 -3068 1717
rect -3102 1615 -3068 1649
rect -3102 1547 -3068 1581
rect -3102 1479 -3068 1513
rect -3102 1411 -3068 1445
rect -3102 1343 -3068 1377
rect -3102 1275 -3068 1309
rect -3102 1207 -3068 1241
rect -3102 1139 -3068 1173
rect -3102 1071 -3068 1105
rect -3102 1003 -3068 1037
rect -3102 935 -3068 969
rect -3102 867 -3068 901
rect -3102 799 -3068 833
rect -3102 731 -3068 765
rect -3102 663 -3068 697
rect -3102 595 -3068 629
rect -3102 527 -3068 561
rect -3102 459 -3068 493
rect -3102 391 -3068 425
rect -3102 323 -3068 357
rect -3102 255 -3068 289
rect -3102 187 -3068 221
rect -3102 119 -3068 153
rect -3102 51 -3068 85
rect -3102 -17 -3068 17
rect -3102 -85 -3068 -51
rect -3102 -153 -3068 -119
rect -3102 -221 -3068 -187
rect -3102 -289 -3068 -255
rect -3102 -357 -3068 -323
rect -3102 -425 -3068 -391
rect -3102 -493 -3068 -459
rect -3102 -561 -3068 -527
rect -3102 -629 -3068 -595
rect -3102 -697 -3068 -663
rect -3102 -765 -3068 -731
rect -3102 -833 -3068 -799
rect -3102 -901 -3068 -867
rect -3102 -969 -3068 -935
rect -3102 -1037 -3068 -1003
rect -3102 -1105 -3068 -1071
rect -3102 -1173 -3068 -1139
rect -3102 -1241 -3068 -1207
rect -3102 -1309 -3068 -1275
rect -3102 -1377 -3068 -1343
rect -3102 -1445 -3068 -1411
rect -3102 -1513 -3068 -1479
rect -3102 -1581 -3068 -1547
rect -3102 -1649 -3068 -1615
rect -3102 -1717 -3068 -1683
rect -3102 -1785 -3068 -1751
rect -3102 -1853 -3068 -1819
rect -3102 -1921 -3068 -1887
rect -3102 -1989 -3068 -1955
rect -3102 -2057 -3068 -2023
rect -3102 -2125 -3068 -2091
rect -3102 -2193 -3068 -2159
rect -3102 -2261 -3068 -2227
rect -3102 -2329 -3068 -2295
rect -3102 -2397 -3068 -2363
rect -3102 -2465 -3068 -2431
rect -3102 -2533 -3068 -2499
rect -3102 -2601 -3068 -2567
rect -3102 -2669 -3068 -2635
rect -3102 -2737 -3068 -2703
rect -3102 -2805 -3068 -2771
rect -3102 -2873 -3068 -2839
rect -3102 -2941 -3068 -2907
rect -3102 -3068 -3068 -2975
rect 3068 2975 3102 3068
rect 3068 2907 3102 2941
rect 3068 2839 3102 2873
rect 3068 2771 3102 2805
rect 3068 2703 3102 2737
rect 3068 2635 3102 2669
rect 3068 2567 3102 2601
rect 3068 2499 3102 2533
rect 3068 2431 3102 2465
rect 3068 2363 3102 2397
rect 3068 2295 3102 2329
rect 3068 2227 3102 2261
rect 3068 2159 3102 2193
rect 3068 2091 3102 2125
rect 3068 2023 3102 2057
rect 3068 1955 3102 1989
rect 3068 1887 3102 1921
rect 3068 1819 3102 1853
rect 3068 1751 3102 1785
rect 3068 1683 3102 1717
rect 3068 1615 3102 1649
rect 3068 1547 3102 1581
rect 3068 1479 3102 1513
rect 3068 1411 3102 1445
rect 3068 1343 3102 1377
rect 3068 1275 3102 1309
rect 3068 1207 3102 1241
rect 3068 1139 3102 1173
rect 3068 1071 3102 1105
rect 3068 1003 3102 1037
rect 3068 935 3102 969
rect 3068 867 3102 901
rect 3068 799 3102 833
rect 3068 731 3102 765
rect 3068 663 3102 697
rect 3068 595 3102 629
rect 3068 527 3102 561
rect 3068 459 3102 493
rect 3068 391 3102 425
rect 3068 323 3102 357
rect 3068 255 3102 289
rect 3068 187 3102 221
rect 3068 119 3102 153
rect 3068 51 3102 85
rect 3068 -17 3102 17
rect 3068 -85 3102 -51
rect 3068 -153 3102 -119
rect 3068 -221 3102 -187
rect 3068 -289 3102 -255
rect 3068 -357 3102 -323
rect 3068 -425 3102 -391
rect 3068 -493 3102 -459
rect 3068 -561 3102 -527
rect 3068 -629 3102 -595
rect 3068 -697 3102 -663
rect 3068 -765 3102 -731
rect 3068 -833 3102 -799
rect 3068 -901 3102 -867
rect 3068 -969 3102 -935
rect 3068 -1037 3102 -1003
rect 3068 -1105 3102 -1071
rect 3068 -1173 3102 -1139
rect 3068 -1241 3102 -1207
rect 3068 -1309 3102 -1275
rect 3068 -1377 3102 -1343
rect 3068 -1445 3102 -1411
rect 3068 -1513 3102 -1479
rect 3068 -1581 3102 -1547
rect 3068 -1649 3102 -1615
rect 3068 -1717 3102 -1683
rect 3068 -1785 3102 -1751
rect 3068 -1853 3102 -1819
rect 3068 -1921 3102 -1887
rect 3068 -1989 3102 -1955
rect 3068 -2057 3102 -2023
rect 3068 -2125 3102 -2091
rect 3068 -2193 3102 -2159
rect 3068 -2261 3102 -2227
rect 3068 -2329 3102 -2295
rect 3068 -2397 3102 -2363
rect 3068 -2465 3102 -2431
rect 3068 -2533 3102 -2499
rect 3068 -2601 3102 -2567
rect 3068 -2669 3102 -2635
rect 3068 -2737 3102 -2703
rect 3068 -2805 3102 -2771
rect 3068 -2873 3102 -2839
rect 3068 -2941 3102 -2907
rect 3068 -3068 3102 -2975
rect -3102 -3102 -2975 -3068
rect -2941 -3102 -2907 -3068
rect -2873 -3102 -2839 -3068
rect -2805 -3102 -2771 -3068
rect -2737 -3102 -2703 -3068
rect -2669 -3102 -2635 -3068
rect -2601 -3102 -2567 -3068
rect -2533 -3102 -2499 -3068
rect -2465 -3102 -2431 -3068
rect -2397 -3102 -2363 -3068
rect -2329 -3102 -2295 -3068
rect -2261 -3102 -2227 -3068
rect -2193 -3102 -2159 -3068
rect -2125 -3102 -2091 -3068
rect -2057 -3102 -2023 -3068
rect -1989 -3102 -1955 -3068
rect -1921 -3102 -1887 -3068
rect -1853 -3102 -1819 -3068
rect -1785 -3102 -1751 -3068
rect -1717 -3102 -1683 -3068
rect -1649 -3102 -1615 -3068
rect -1581 -3102 -1547 -3068
rect -1513 -3102 -1479 -3068
rect -1445 -3102 -1411 -3068
rect -1377 -3102 -1343 -3068
rect -1309 -3102 -1275 -3068
rect -1241 -3102 -1207 -3068
rect -1173 -3102 -1139 -3068
rect -1105 -3102 -1071 -3068
rect -1037 -3102 -1003 -3068
rect -969 -3102 -935 -3068
rect -901 -3102 -867 -3068
rect -833 -3102 -799 -3068
rect -765 -3102 -731 -3068
rect -697 -3102 -663 -3068
rect -629 -3102 -595 -3068
rect -561 -3102 -527 -3068
rect -493 -3102 -459 -3068
rect -425 -3102 -391 -3068
rect -357 -3102 -323 -3068
rect -289 -3102 -255 -3068
rect -221 -3102 -187 -3068
rect -153 -3102 -119 -3068
rect -85 -3102 -51 -3068
rect -17 -3102 17 -3068
rect 51 -3102 85 -3068
rect 119 -3102 153 -3068
rect 187 -3102 221 -3068
rect 255 -3102 289 -3068
rect 323 -3102 357 -3068
rect 391 -3102 425 -3068
rect 459 -3102 493 -3068
rect 527 -3102 561 -3068
rect 595 -3102 629 -3068
rect 663 -3102 697 -3068
rect 731 -3102 765 -3068
rect 799 -3102 833 -3068
rect 867 -3102 901 -3068
rect 935 -3102 969 -3068
rect 1003 -3102 1037 -3068
rect 1071 -3102 1105 -3068
rect 1139 -3102 1173 -3068
rect 1207 -3102 1241 -3068
rect 1275 -3102 1309 -3068
rect 1343 -3102 1377 -3068
rect 1411 -3102 1445 -3068
rect 1479 -3102 1513 -3068
rect 1547 -3102 1581 -3068
rect 1615 -3102 1649 -3068
rect 1683 -3102 1717 -3068
rect 1751 -3102 1785 -3068
rect 1819 -3102 1853 -3068
rect 1887 -3102 1921 -3068
rect 1955 -3102 1989 -3068
rect 2023 -3102 2057 -3068
rect 2091 -3102 2125 -3068
rect 2159 -3102 2193 -3068
rect 2227 -3102 2261 -3068
rect 2295 -3102 2329 -3068
rect 2363 -3102 2397 -3068
rect 2431 -3102 2465 -3068
rect 2499 -3102 2533 -3068
rect 2567 -3102 2601 -3068
rect 2635 -3102 2669 -3068
rect 2703 -3102 2737 -3068
rect 2771 -3102 2805 -3068
rect 2839 -3102 2873 -3068
rect 2907 -3102 2941 -3068
rect 2975 -3102 3102 -3068
<< psubdiffcont >>
rect -3111 3206 -3077 3240
rect -3043 3206 -3009 3240
rect -2975 3206 -2941 3240
rect -2907 3206 -2873 3240
rect -2839 3206 -2805 3240
rect -2771 3206 -2737 3240
rect -2703 3206 -2669 3240
rect -2635 3206 -2601 3240
rect -2567 3206 -2533 3240
rect -2499 3206 -2465 3240
rect -2431 3206 -2397 3240
rect -2363 3206 -2329 3240
rect -2295 3206 -2261 3240
rect -2227 3206 -2193 3240
rect -2159 3206 -2125 3240
rect -2091 3206 -2057 3240
rect -2023 3206 -1989 3240
rect -1955 3206 -1921 3240
rect -1887 3206 -1853 3240
rect -1819 3206 -1785 3240
rect -1751 3206 -1717 3240
rect -1683 3206 -1649 3240
rect -1615 3206 -1581 3240
rect -1547 3206 -1513 3240
rect -1479 3206 -1445 3240
rect -1411 3206 -1377 3240
rect -1343 3206 -1309 3240
rect -1275 3206 -1241 3240
rect -1207 3206 -1173 3240
rect -1139 3206 -1105 3240
rect -1071 3206 -1037 3240
rect -1003 3206 -969 3240
rect -935 3206 -901 3240
rect -867 3206 -833 3240
rect -799 3206 -765 3240
rect -731 3206 -697 3240
rect -663 3206 -629 3240
rect -595 3206 -561 3240
rect -527 3206 -493 3240
rect -459 3206 -425 3240
rect -391 3206 -357 3240
rect -323 3206 -289 3240
rect -255 3206 -221 3240
rect -187 3206 -153 3240
rect -119 3206 -85 3240
rect -51 3206 -17 3240
rect 17 3206 51 3240
rect 85 3206 119 3240
rect 153 3206 187 3240
rect 221 3206 255 3240
rect 289 3206 323 3240
rect 357 3206 391 3240
rect 425 3206 459 3240
rect 493 3206 527 3240
rect 561 3206 595 3240
rect 629 3206 663 3240
rect 697 3206 731 3240
rect 765 3206 799 3240
rect 833 3206 867 3240
rect 901 3206 935 3240
rect 969 3206 1003 3240
rect 1037 3206 1071 3240
rect 1105 3206 1139 3240
rect 1173 3206 1207 3240
rect 1241 3206 1275 3240
rect 1309 3206 1343 3240
rect 1377 3206 1411 3240
rect 1445 3206 1479 3240
rect 1513 3206 1547 3240
rect 1581 3206 1615 3240
rect 1649 3206 1683 3240
rect 1717 3206 1751 3240
rect 1785 3206 1819 3240
rect 1853 3206 1887 3240
rect 1921 3206 1955 3240
rect 1989 3206 2023 3240
rect 2057 3206 2091 3240
rect 2125 3206 2159 3240
rect 2193 3206 2227 3240
rect 2261 3206 2295 3240
rect 2329 3206 2363 3240
rect 2397 3206 2431 3240
rect 2465 3206 2499 3240
rect 2533 3206 2567 3240
rect 2601 3206 2635 3240
rect 2669 3206 2703 3240
rect 2737 3206 2771 3240
rect 2805 3206 2839 3240
rect 2873 3206 2907 3240
rect 2941 3206 2975 3240
rect 3009 3206 3043 3240
rect 3077 3206 3111 3240
rect -3240 3077 -3206 3111
rect -3240 3009 -3206 3043
rect -3240 2941 -3206 2975
rect -3240 2873 -3206 2907
rect -3240 2805 -3206 2839
rect -3240 2737 -3206 2771
rect -3240 2669 -3206 2703
rect -3240 2601 -3206 2635
rect -3240 2533 -3206 2567
rect -3240 2465 -3206 2499
rect -3240 2397 -3206 2431
rect -3240 2329 -3206 2363
rect -3240 2261 -3206 2295
rect -3240 2193 -3206 2227
rect -3240 2125 -3206 2159
rect -3240 2057 -3206 2091
rect -3240 1989 -3206 2023
rect -3240 1921 -3206 1955
rect -3240 1853 -3206 1887
rect -3240 1785 -3206 1819
rect -3240 1717 -3206 1751
rect -3240 1649 -3206 1683
rect -3240 1581 -3206 1615
rect -3240 1513 -3206 1547
rect -3240 1445 -3206 1479
rect -3240 1377 -3206 1411
rect -3240 1309 -3206 1343
rect -3240 1241 -3206 1275
rect -3240 1173 -3206 1207
rect -3240 1105 -3206 1139
rect -3240 1037 -3206 1071
rect -3240 969 -3206 1003
rect -3240 901 -3206 935
rect -3240 833 -3206 867
rect -3240 765 -3206 799
rect -3240 697 -3206 731
rect -3240 629 -3206 663
rect -3240 561 -3206 595
rect -3240 493 -3206 527
rect -3240 425 -3206 459
rect -3240 357 -3206 391
rect -3240 289 -3206 323
rect -3240 221 -3206 255
rect -3240 153 -3206 187
rect -3240 85 -3206 119
rect -3240 17 -3206 51
rect -3240 -51 -3206 -17
rect -3240 -119 -3206 -85
rect -3240 -187 -3206 -153
rect -3240 -255 -3206 -221
rect -3240 -323 -3206 -289
rect -3240 -391 -3206 -357
rect -3240 -459 -3206 -425
rect -3240 -527 -3206 -493
rect -3240 -595 -3206 -561
rect -3240 -663 -3206 -629
rect -3240 -731 -3206 -697
rect -3240 -799 -3206 -765
rect -3240 -867 -3206 -833
rect -3240 -935 -3206 -901
rect -3240 -1003 -3206 -969
rect -3240 -1071 -3206 -1037
rect -3240 -1139 -3206 -1105
rect -3240 -1207 -3206 -1173
rect -3240 -1275 -3206 -1241
rect -3240 -1343 -3206 -1309
rect -3240 -1411 -3206 -1377
rect -3240 -1479 -3206 -1445
rect -3240 -1547 -3206 -1513
rect -3240 -1615 -3206 -1581
rect -3240 -1683 -3206 -1649
rect -3240 -1751 -3206 -1717
rect -3240 -1819 -3206 -1785
rect -3240 -1887 -3206 -1853
rect -3240 -1955 -3206 -1921
rect -3240 -2023 -3206 -1989
rect -3240 -2091 -3206 -2057
rect -3240 -2159 -3206 -2125
rect -3240 -2227 -3206 -2193
rect -3240 -2295 -3206 -2261
rect -3240 -2363 -3206 -2329
rect -3240 -2431 -3206 -2397
rect -3240 -2499 -3206 -2465
rect -3240 -2567 -3206 -2533
rect -3240 -2635 -3206 -2601
rect -3240 -2703 -3206 -2669
rect -3240 -2771 -3206 -2737
rect -3240 -2839 -3206 -2805
rect -3240 -2907 -3206 -2873
rect -3240 -2975 -3206 -2941
rect -3240 -3043 -3206 -3009
rect -3240 -3111 -3206 -3077
rect 3206 3077 3240 3111
rect 3206 3009 3240 3043
rect 3206 2941 3240 2975
rect 3206 2873 3240 2907
rect 3206 2805 3240 2839
rect 3206 2737 3240 2771
rect 3206 2669 3240 2703
rect 3206 2601 3240 2635
rect 3206 2533 3240 2567
rect 3206 2465 3240 2499
rect 3206 2397 3240 2431
rect 3206 2329 3240 2363
rect 3206 2261 3240 2295
rect 3206 2193 3240 2227
rect 3206 2125 3240 2159
rect 3206 2057 3240 2091
rect 3206 1989 3240 2023
rect 3206 1921 3240 1955
rect 3206 1853 3240 1887
rect 3206 1785 3240 1819
rect 3206 1717 3240 1751
rect 3206 1649 3240 1683
rect 3206 1581 3240 1615
rect 3206 1513 3240 1547
rect 3206 1445 3240 1479
rect 3206 1377 3240 1411
rect 3206 1309 3240 1343
rect 3206 1241 3240 1275
rect 3206 1173 3240 1207
rect 3206 1105 3240 1139
rect 3206 1037 3240 1071
rect 3206 969 3240 1003
rect 3206 901 3240 935
rect 3206 833 3240 867
rect 3206 765 3240 799
rect 3206 697 3240 731
rect 3206 629 3240 663
rect 3206 561 3240 595
rect 3206 493 3240 527
rect 3206 425 3240 459
rect 3206 357 3240 391
rect 3206 289 3240 323
rect 3206 221 3240 255
rect 3206 153 3240 187
rect 3206 85 3240 119
rect 3206 17 3240 51
rect 3206 -51 3240 -17
rect 3206 -119 3240 -85
rect 3206 -187 3240 -153
rect 3206 -255 3240 -221
rect 3206 -323 3240 -289
rect 3206 -391 3240 -357
rect 3206 -459 3240 -425
rect 3206 -527 3240 -493
rect 3206 -595 3240 -561
rect 3206 -663 3240 -629
rect 3206 -731 3240 -697
rect 3206 -799 3240 -765
rect 3206 -867 3240 -833
rect 3206 -935 3240 -901
rect 3206 -1003 3240 -969
rect 3206 -1071 3240 -1037
rect 3206 -1139 3240 -1105
rect 3206 -1207 3240 -1173
rect 3206 -1275 3240 -1241
rect 3206 -1343 3240 -1309
rect 3206 -1411 3240 -1377
rect 3206 -1479 3240 -1445
rect 3206 -1547 3240 -1513
rect 3206 -1615 3240 -1581
rect 3206 -1683 3240 -1649
rect 3206 -1751 3240 -1717
rect 3206 -1819 3240 -1785
rect 3206 -1887 3240 -1853
rect 3206 -1955 3240 -1921
rect 3206 -2023 3240 -1989
rect 3206 -2091 3240 -2057
rect 3206 -2159 3240 -2125
rect 3206 -2227 3240 -2193
rect 3206 -2295 3240 -2261
rect 3206 -2363 3240 -2329
rect 3206 -2431 3240 -2397
rect 3206 -2499 3240 -2465
rect 3206 -2567 3240 -2533
rect 3206 -2635 3240 -2601
rect 3206 -2703 3240 -2669
rect 3206 -2771 3240 -2737
rect 3206 -2839 3240 -2805
rect 3206 -2907 3240 -2873
rect 3206 -2975 3240 -2941
rect 3206 -3043 3240 -3009
rect 3206 -3111 3240 -3077
rect -3111 -3240 -3077 -3206
rect -3043 -3240 -3009 -3206
rect -2975 -3240 -2941 -3206
rect -2907 -3240 -2873 -3206
rect -2839 -3240 -2805 -3206
rect -2771 -3240 -2737 -3206
rect -2703 -3240 -2669 -3206
rect -2635 -3240 -2601 -3206
rect -2567 -3240 -2533 -3206
rect -2499 -3240 -2465 -3206
rect -2431 -3240 -2397 -3206
rect -2363 -3240 -2329 -3206
rect -2295 -3240 -2261 -3206
rect -2227 -3240 -2193 -3206
rect -2159 -3240 -2125 -3206
rect -2091 -3240 -2057 -3206
rect -2023 -3240 -1989 -3206
rect -1955 -3240 -1921 -3206
rect -1887 -3240 -1853 -3206
rect -1819 -3240 -1785 -3206
rect -1751 -3240 -1717 -3206
rect -1683 -3240 -1649 -3206
rect -1615 -3240 -1581 -3206
rect -1547 -3240 -1513 -3206
rect -1479 -3240 -1445 -3206
rect -1411 -3240 -1377 -3206
rect -1343 -3240 -1309 -3206
rect -1275 -3240 -1241 -3206
rect -1207 -3240 -1173 -3206
rect -1139 -3240 -1105 -3206
rect -1071 -3240 -1037 -3206
rect -1003 -3240 -969 -3206
rect -935 -3240 -901 -3206
rect -867 -3240 -833 -3206
rect -799 -3240 -765 -3206
rect -731 -3240 -697 -3206
rect -663 -3240 -629 -3206
rect -595 -3240 -561 -3206
rect -527 -3240 -493 -3206
rect -459 -3240 -425 -3206
rect -391 -3240 -357 -3206
rect -323 -3240 -289 -3206
rect -255 -3240 -221 -3206
rect -187 -3240 -153 -3206
rect -119 -3240 -85 -3206
rect -51 -3240 -17 -3206
rect 17 -3240 51 -3206
rect 85 -3240 119 -3206
rect 153 -3240 187 -3206
rect 221 -3240 255 -3206
rect 289 -3240 323 -3206
rect 357 -3240 391 -3206
rect 425 -3240 459 -3206
rect 493 -3240 527 -3206
rect 561 -3240 595 -3206
rect 629 -3240 663 -3206
rect 697 -3240 731 -3206
rect 765 -3240 799 -3206
rect 833 -3240 867 -3206
rect 901 -3240 935 -3206
rect 969 -3240 1003 -3206
rect 1037 -3240 1071 -3206
rect 1105 -3240 1139 -3206
rect 1173 -3240 1207 -3206
rect 1241 -3240 1275 -3206
rect 1309 -3240 1343 -3206
rect 1377 -3240 1411 -3206
rect 1445 -3240 1479 -3206
rect 1513 -3240 1547 -3206
rect 1581 -3240 1615 -3206
rect 1649 -3240 1683 -3206
rect 1717 -3240 1751 -3206
rect 1785 -3240 1819 -3206
rect 1853 -3240 1887 -3206
rect 1921 -3240 1955 -3206
rect 1989 -3240 2023 -3206
rect 2057 -3240 2091 -3206
rect 2125 -3240 2159 -3206
rect 2193 -3240 2227 -3206
rect 2261 -3240 2295 -3206
rect 2329 -3240 2363 -3206
rect 2397 -3240 2431 -3206
rect 2465 -3240 2499 -3206
rect 2533 -3240 2567 -3206
rect 2601 -3240 2635 -3206
rect 2669 -3240 2703 -3206
rect 2737 -3240 2771 -3206
rect 2805 -3240 2839 -3206
rect 2873 -3240 2907 -3206
rect 2941 -3240 2975 -3206
rect 3009 -3240 3043 -3206
rect 3077 -3240 3111 -3206
<< nsubdiffcont >>
rect -2975 3068 -2941 3102
rect -2907 3068 -2873 3102
rect -2839 3068 -2805 3102
rect -2771 3068 -2737 3102
rect -2703 3068 -2669 3102
rect -2635 3068 -2601 3102
rect -2567 3068 -2533 3102
rect -2499 3068 -2465 3102
rect -2431 3068 -2397 3102
rect -2363 3068 -2329 3102
rect -2295 3068 -2261 3102
rect -2227 3068 -2193 3102
rect -2159 3068 -2125 3102
rect -2091 3068 -2057 3102
rect -2023 3068 -1989 3102
rect -1955 3068 -1921 3102
rect -1887 3068 -1853 3102
rect -1819 3068 -1785 3102
rect -1751 3068 -1717 3102
rect -1683 3068 -1649 3102
rect -1615 3068 -1581 3102
rect -1547 3068 -1513 3102
rect -1479 3068 -1445 3102
rect -1411 3068 -1377 3102
rect -1343 3068 -1309 3102
rect -1275 3068 -1241 3102
rect -1207 3068 -1173 3102
rect -1139 3068 -1105 3102
rect -1071 3068 -1037 3102
rect -1003 3068 -969 3102
rect -935 3068 -901 3102
rect -867 3068 -833 3102
rect -799 3068 -765 3102
rect -731 3068 -697 3102
rect -663 3068 -629 3102
rect -595 3068 -561 3102
rect -527 3068 -493 3102
rect -459 3068 -425 3102
rect -391 3068 -357 3102
rect -323 3068 -289 3102
rect -255 3068 -221 3102
rect -187 3068 -153 3102
rect -119 3068 -85 3102
rect -51 3068 -17 3102
rect 17 3068 51 3102
rect 85 3068 119 3102
rect 153 3068 187 3102
rect 221 3068 255 3102
rect 289 3068 323 3102
rect 357 3068 391 3102
rect 425 3068 459 3102
rect 493 3068 527 3102
rect 561 3068 595 3102
rect 629 3068 663 3102
rect 697 3068 731 3102
rect 765 3068 799 3102
rect 833 3068 867 3102
rect 901 3068 935 3102
rect 969 3068 1003 3102
rect 1037 3068 1071 3102
rect 1105 3068 1139 3102
rect 1173 3068 1207 3102
rect 1241 3068 1275 3102
rect 1309 3068 1343 3102
rect 1377 3068 1411 3102
rect 1445 3068 1479 3102
rect 1513 3068 1547 3102
rect 1581 3068 1615 3102
rect 1649 3068 1683 3102
rect 1717 3068 1751 3102
rect 1785 3068 1819 3102
rect 1853 3068 1887 3102
rect 1921 3068 1955 3102
rect 1989 3068 2023 3102
rect 2057 3068 2091 3102
rect 2125 3068 2159 3102
rect 2193 3068 2227 3102
rect 2261 3068 2295 3102
rect 2329 3068 2363 3102
rect 2397 3068 2431 3102
rect 2465 3068 2499 3102
rect 2533 3068 2567 3102
rect 2601 3068 2635 3102
rect 2669 3068 2703 3102
rect 2737 3068 2771 3102
rect 2805 3068 2839 3102
rect 2873 3068 2907 3102
rect 2941 3068 2975 3102
rect -3102 2941 -3068 2975
rect -3102 2873 -3068 2907
rect -3102 2805 -3068 2839
rect -3102 2737 -3068 2771
rect -3102 2669 -3068 2703
rect -3102 2601 -3068 2635
rect -3102 2533 -3068 2567
rect -3102 2465 -3068 2499
rect -3102 2397 -3068 2431
rect -3102 2329 -3068 2363
rect -3102 2261 -3068 2295
rect -3102 2193 -3068 2227
rect -3102 2125 -3068 2159
rect -3102 2057 -3068 2091
rect -3102 1989 -3068 2023
rect -3102 1921 -3068 1955
rect -3102 1853 -3068 1887
rect -3102 1785 -3068 1819
rect -3102 1717 -3068 1751
rect -3102 1649 -3068 1683
rect -3102 1581 -3068 1615
rect -3102 1513 -3068 1547
rect -3102 1445 -3068 1479
rect -3102 1377 -3068 1411
rect -3102 1309 -3068 1343
rect -3102 1241 -3068 1275
rect -3102 1173 -3068 1207
rect -3102 1105 -3068 1139
rect -3102 1037 -3068 1071
rect -3102 969 -3068 1003
rect -3102 901 -3068 935
rect -3102 833 -3068 867
rect -3102 765 -3068 799
rect -3102 697 -3068 731
rect -3102 629 -3068 663
rect -3102 561 -3068 595
rect -3102 493 -3068 527
rect -3102 425 -3068 459
rect -3102 357 -3068 391
rect -3102 289 -3068 323
rect -3102 221 -3068 255
rect -3102 153 -3068 187
rect -3102 85 -3068 119
rect -3102 17 -3068 51
rect -3102 -51 -3068 -17
rect -3102 -119 -3068 -85
rect -3102 -187 -3068 -153
rect -3102 -255 -3068 -221
rect -3102 -323 -3068 -289
rect -3102 -391 -3068 -357
rect -3102 -459 -3068 -425
rect -3102 -527 -3068 -493
rect -3102 -595 -3068 -561
rect -3102 -663 -3068 -629
rect -3102 -731 -3068 -697
rect -3102 -799 -3068 -765
rect -3102 -867 -3068 -833
rect -3102 -935 -3068 -901
rect -3102 -1003 -3068 -969
rect -3102 -1071 -3068 -1037
rect -3102 -1139 -3068 -1105
rect -3102 -1207 -3068 -1173
rect -3102 -1275 -3068 -1241
rect -3102 -1343 -3068 -1309
rect -3102 -1411 -3068 -1377
rect -3102 -1479 -3068 -1445
rect -3102 -1547 -3068 -1513
rect -3102 -1615 -3068 -1581
rect -3102 -1683 -3068 -1649
rect -3102 -1751 -3068 -1717
rect -3102 -1819 -3068 -1785
rect -3102 -1887 -3068 -1853
rect -3102 -1955 -3068 -1921
rect -3102 -2023 -3068 -1989
rect -3102 -2091 -3068 -2057
rect -3102 -2159 -3068 -2125
rect -3102 -2227 -3068 -2193
rect -3102 -2295 -3068 -2261
rect -3102 -2363 -3068 -2329
rect -3102 -2431 -3068 -2397
rect -3102 -2499 -3068 -2465
rect -3102 -2567 -3068 -2533
rect -3102 -2635 -3068 -2601
rect -3102 -2703 -3068 -2669
rect -3102 -2771 -3068 -2737
rect -3102 -2839 -3068 -2805
rect -3102 -2907 -3068 -2873
rect -3102 -2975 -3068 -2941
rect 3068 2941 3102 2975
rect 3068 2873 3102 2907
rect 3068 2805 3102 2839
rect 3068 2737 3102 2771
rect 3068 2669 3102 2703
rect 3068 2601 3102 2635
rect 3068 2533 3102 2567
rect 3068 2465 3102 2499
rect 3068 2397 3102 2431
rect 3068 2329 3102 2363
rect 3068 2261 3102 2295
rect 3068 2193 3102 2227
rect 3068 2125 3102 2159
rect 3068 2057 3102 2091
rect 3068 1989 3102 2023
rect 3068 1921 3102 1955
rect 3068 1853 3102 1887
rect 3068 1785 3102 1819
rect 3068 1717 3102 1751
rect 3068 1649 3102 1683
rect 3068 1581 3102 1615
rect 3068 1513 3102 1547
rect 3068 1445 3102 1479
rect 3068 1377 3102 1411
rect 3068 1309 3102 1343
rect 3068 1241 3102 1275
rect 3068 1173 3102 1207
rect 3068 1105 3102 1139
rect 3068 1037 3102 1071
rect 3068 969 3102 1003
rect 3068 901 3102 935
rect 3068 833 3102 867
rect 3068 765 3102 799
rect 3068 697 3102 731
rect 3068 629 3102 663
rect 3068 561 3102 595
rect 3068 493 3102 527
rect 3068 425 3102 459
rect 3068 357 3102 391
rect 3068 289 3102 323
rect 3068 221 3102 255
rect 3068 153 3102 187
rect 3068 85 3102 119
rect 3068 17 3102 51
rect 3068 -51 3102 -17
rect 3068 -119 3102 -85
rect 3068 -187 3102 -153
rect 3068 -255 3102 -221
rect 3068 -323 3102 -289
rect 3068 -391 3102 -357
rect 3068 -459 3102 -425
rect 3068 -527 3102 -493
rect 3068 -595 3102 -561
rect 3068 -663 3102 -629
rect 3068 -731 3102 -697
rect 3068 -799 3102 -765
rect 3068 -867 3102 -833
rect 3068 -935 3102 -901
rect 3068 -1003 3102 -969
rect 3068 -1071 3102 -1037
rect 3068 -1139 3102 -1105
rect 3068 -1207 3102 -1173
rect 3068 -1275 3102 -1241
rect 3068 -1343 3102 -1309
rect 3068 -1411 3102 -1377
rect 3068 -1479 3102 -1445
rect 3068 -1547 3102 -1513
rect 3068 -1615 3102 -1581
rect 3068 -1683 3102 -1649
rect 3068 -1751 3102 -1717
rect 3068 -1819 3102 -1785
rect 3068 -1887 3102 -1853
rect 3068 -1955 3102 -1921
rect 3068 -2023 3102 -1989
rect 3068 -2091 3102 -2057
rect 3068 -2159 3102 -2125
rect 3068 -2227 3102 -2193
rect 3068 -2295 3102 -2261
rect 3068 -2363 3102 -2329
rect 3068 -2431 3102 -2397
rect 3068 -2499 3102 -2465
rect 3068 -2567 3102 -2533
rect 3068 -2635 3102 -2601
rect 3068 -2703 3102 -2669
rect 3068 -2771 3102 -2737
rect 3068 -2839 3102 -2805
rect 3068 -2907 3102 -2873
rect 3068 -2975 3102 -2941
rect -2975 -3102 -2941 -3068
rect -2907 -3102 -2873 -3068
rect -2839 -3102 -2805 -3068
rect -2771 -3102 -2737 -3068
rect -2703 -3102 -2669 -3068
rect -2635 -3102 -2601 -3068
rect -2567 -3102 -2533 -3068
rect -2499 -3102 -2465 -3068
rect -2431 -3102 -2397 -3068
rect -2363 -3102 -2329 -3068
rect -2295 -3102 -2261 -3068
rect -2227 -3102 -2193 -3068
rect -2159 -3102 -2125 -3068
rect -2091 -3102 -2057 -3068
rect -2023 -3102 -1989 -3068
rect -1955 -3102 -1921 -3068
rect -1887 -3102 -1853 -3068
rect -1819 -3102 -1785 -3068
rect -1751 -3102 -1717 -3068
rect -1683 -3102 -1649 -3068
rect -1615 -3102 -1581 -3068
rect -1547 -3102 -1513 -3068
rect -1479 -3102 -1445 -3068
rect -1411 -3102 -1377 -3068
rect -1343 -3102 -1309 -3068
rect -1275 -3102 -1241 -3068
rect -1207 -3102 -1173 -3068
rect -1139 -3102 -1105 -3068
rect -1071 -3102 -1037 -3068
rect -1003 -3102 -969 -3068
rect -935 -3102 -901 -3068
rect -867 -3102 -833 -3068
rect -799 -3102 -765 -3068
rect -731 -3102 -697 -3068
rect -663 -3102 -629 -3068
rect -595 -3102 -561 -3068
rect -527 -3102 -493 -3068
rect -459 -3102 -425 -3068
rect -391 -3102 -357 -3068
rect -323 -3102 -289 -3068
rect -255 -3102 -221 -3068
rect -187 -3102 -153 -3068
rect -119 -3102 -85 -3068
rect -51 -3102 -17 -3068
rect 17 -3102 51 -3068
rect 85 -3102 119 -3068
rect 153 -3102 187 -3068
rect 221 -3102 255 -3068
rect 289 -3102 323 -3068
rect 357 -3102 391 -3068
rect 425 -3102 459 -3068
rect 493 -3102 527 -3068
rect 561 -3102 595 -3068
rect 629 -3102 663 -3068
rect 697 -3102 731 -3068
rect 765 -3102 799 -3068
rect 833 -3102 867 -3068
rect 901 -3102 935 -3068
rect 969 -3102 1003 -3068
rect 1037 -3102 1071 -3068
rect 1105 -3102 1139 -3068
rect 1173 -3102 1207 -3068
rect 1241 -3102 1275 -3068
rect 1309 -3102 1343 -3068
rect 1377 -3102 1411 -3068
rect 1445 -3102 1479 -3068
rect 1513 -3102 1547 -3068
rect 1581 -3102 1615 -3068
rect 1649 -3102 1683 -3068
rect 1717 -3102 1751 -3068
rect 1785 -3102 1819 -3068
rect 1853 -3102 1887 -3068
rect 1921 -3102 1955 -3068
rect 1989 -3102 2023 -3068
rect 2057 -3102 2091 -3068
rect 2125 -3102 2159 -3068
rect 2193 -3102 2227 -3068
rect 2261 -3102 2295 -3068
rect 2329 -3102 2363 -3068
rect 2397 -3102 2431 -3068
rect 2465 -3102 2499 -3068
rect 2533 -3102 2567 -3068
rect 2601 -3102 2635 -3068
rect 2669 -3102 2703 -3068
rect 2737 -3102 2771 -3068
rect 2805 -3102 2839 -3068
rect 2873 -3102 2907 -3068
rect 2941 -3102 2975 -3068
<< pdiode >>
rect -3000 2975 3000 3000
rect -3000 -2975 -2975 2975
rect 2975 -2975 3000 2975
rect -3000 -3000 3000 -2975
<< pdiodec >>
rect -2975 -2975 2975 2975
<< locali >>
rect -3240 3206 -3111 3240
rect -3077 3206 -3043 3240
rect -3009 3206 -2975 3240
rect -2941 3206 -2907 3240
rect -2873 3206 -2839 3240
rect -2805 3206 -2771 3240
rect -2737 3206 -2703 3240
rect -2669 3206 -2635 3240
rect -2601 3206 -2567 3240
rect -2533 3206 -2499 3240
rect -2465 3206 -2431 3240
rect -2397 3206 -2363 3240
rect -2329 3206 -2295 3240
rect -2261 3206 -2227 3240
rect -2193 3206 -2159 3240
rect -2125 3206 -2091 3240
rect -2057 3206 -2023 3240
rect -1989 3206 -1955 3240
rect -1921 3206 -1887 3240
rect -1853 3206 -1819 3240
rect -1785 3206 -1751 3240
rect -1717 3206 -1683 3240
rect -1649 3206 -1615 3240
rect -1581 3206 -1547 3240
rect -1513 3206 -1479 3240
rect -1445 3206 -1411 3240
rect -1377 3206 -1343 3240
rect -1309 3206 -1275 3240
rect -1241 3206 -1207 3240
rect -1173 3206 -1139 3240
rect -1105 3206 -1071 3240
rect -1037 3206 -1003 3240
rect -969 3206 -935 3240
rect -901 3206 -867 3240
rect -833 3206 -799 3240
rect -765 3206 -731 3240
rect -697 3206 -663 3240
rect -629 3206 -595 3240
rect -561 3206 -527 3240
rect -493 3206 -459 3240
rect -425 3206 -391 3240
rect -357 3206 -323 3240
rect -289 3206 -255 3240
rect -221 3206 -187 3240
rect -153 3206 -119 3240
rect -85 3206 -51 3240
rect -17 3206 17 3240
rect 51 3206 85 3240
rect 119 3206 153 3240
rect 187 3206 221 3240
rect 255 3206 289 3240
rect 323 3206 357 3240
rect 391 3206 425 3240
rect 459 3206 493 3240
rect 527 3206 561 3240
rect 595 3206 629 3240
rect 663 3206 697 3240
rect 731 3206 765 3240
rect 799 3206 833 3240
rect 867 3206 901 3240
rect 935 3206 969 3240
rect 1003 3206 1037 3240
rect 1071 3206 1105 3240
rect 1139 3206 1173 3240
rect 1207 3206 1241 3240
rect 1275 3206 1309 3240
rect 1343 3206 1377 3240
rect 1411 3206 1445 3240
rect 1479 3206 1513 3240
rect 1547 3206 1581 3240
rect 1615 3206 1649 3240
rect 1683 3206 1717 3240
rect 1751 3206 1785 3240
rect 1819 3206 1853 3240
rect 1887 3206 1921 3240
rect 1955 3206 1989 3240
rect 2023 3206 2057 3240
rect 2091 3206 2125 3240
rect 2159 3206 2193 3240
rect 2227 3206 2261 3240
rect 2295 3206 2329 3240
rect 2363 3206 2397 3240
rect 2431 3206 2465 3240
rect 2499 3206 2533 3240
rect 2567 3206 2601 3240
rect 2635 3206 2669 3240
rect 2703 3206 2737 3240
rect 2771 3206 2805 3240
rect 2839 3206 2873 3240
rect 2907 3206 2941 3240
rect 2975 3206 3009 3240
rect 3043 3206 3077 3240
rect 3111 3206 3240 3240
rect -3240 3111 -3206 3206
rect 3206 3111 3240 3206
rect -3240 3043 -3206 3077
rect -3240 2975 -3206 3009
rect -3240 2907 -3206 2941
rect -3240 2839 -3206 2873
rect -3240 2771 -3206 2805
rect -3240 2703 -3206 2737
rect -3240 2635 -3206 2669
rect -3240 2567 -3206 2601
rect -3240 2499 -3206 2533
rect -3240 2431 -3206 2465
rect -3240 2363 -3206 2397
rect -3240 2295 -3206 2329
rect -3240 2227 -3206 2261
rect -3240 2159 -3206 2193
rect -3240 2091 -3206 2125
rect -3240 2023 -3206 2057
rect -3240 1955 -3206 1989
rect -3240 1887 -3206 1921
rect -3240 1819 -3206 1853
rect -3240 1751 -3206 1785
rect -3240 1683 -3206 1717
rect -3240 1615 -3206 1649
rect -3240 1547 -3206 1581
rect -3240 1479 -3206 1513
rect -3240 1411 -3206 1445
rect -3240 1343 -3206 1377
rect -3240 1275 -3206 1309
rect -3240 1207 -3206 1241
rect -3240 1139 -3206 1173
rect -3240 1071 -3206 1105
rect -3240 1003 -3206 1037
rect -3240 935 -3206 969
rect -3240 867 -3206 901
rect -3240 799 -3206 833
rect -3240 731 -3206 765
rect -3240 663 -3206 697
rect -3240 595 -3206 629
rect -3240 527 -3206 561
rect -3240 459 -3206 493
rect -3240 391 -3206 425
rect -3240 323 -3206 357
rect -3240 255 -3206 289
rect -3240 187 -3206 221
rect -3240 119 -3206 153
rect -3240 51 -3206 85
rect -3240 -17 -3206 17
rect -3240 -85 -3206 -51
rect -3240 -153 -3206 -119
rect -3240 -221 -3206 -187
rect -3240 -289 -3206 -255
rect -3240 -357 -3206 -323
rect -3240 -425 -3206 -391
rect -3240 -493 -3206 -459
rect -3240 -561 -3206 -527
rect -3240 -629 -3206 -595
rect -3240 -697 -3206 -663
rect -3240 -765 -3206 -731
rect -3240 -833 -3206 -799
rect -3240 -901 -3206 -867
rect -3240 -969 -3206 -935
rect -3240 -1037 -3206 -1003
rect -3240 -1105 -3206 -1071
rect -3240 -1173 -3206 -1139
rect -3240 -1241 -3206 -1207
rect -3240 -1309 -3206 -1275
rect -3240 -1377 -3206 -1343
rect -3240 -1445 -3206 -1411
rect -3240 -1513 -3206 -1479
rect -3240 -1581 -3206 -1547
rect -3240 -1649 -3206 -1615
rect -3240 -1717 -3206 -1683
rect -3240 -1785 -3206 -1751
rect -3240 -1853 -3206 -1819
rect -3240 -1921 -3206 -1887
rect -3240 -1989 -3206 -1955
rect -3240 -2057 -3206 -2023
rect -3240 -2125 -3206 -2091
rect -3240 -2193 -3206 -2159
rect -3240 -2261 -3206 -2227
rect -3240 -2329 -3206 -2295
rect -3240 -2397 -3206 -2363
rect -3240 -2465 -3206 -2431
rect -3240 -2533 -3206 -2499
rect -3240 -2601 -3206 -2567
rect -3240 -2669 -3206 -2635
rect -3240 -2737 -3206 -2703
rect -3240 -2805 -3206 -2771
rect -3240 -2873 -3206 -2839
rect -3240 -2941 -3206 -2907
rect -3240 -3009 -3206 -2975
rect -3240 -3077 -3206 -3043
rect -3102 3068 -2975 3102
rect -2941 3068 -2907 3102
rect -2873 3068 -2839 3102
rect -2805 3068 -2771 3102
rect -2737 3068 -2703 3102
rect -2669 3068 -2635 3102
rect -2601 3068 -2567 3102
rect -2533 3068 -2499 3102
rect -2465 3068 -2431 3102
rect -2397 3068 -2363 3102
rect -2329 3068 -2295 3102
rect -2261 3068 -2227 3102
rect -2193 3068 -2159 3102
rect -2125 3068 -2091 3102
rect -2057 3068 -2023 3102
rect -1989 3068 -1955 3102
rect -1921 3068 -1887 3102
rect -1853 3068 -1819 3102
rect -1785 3068 -1751 3102
rect -1717 3068 -1683 3102
rect -1649 3068 -1615 3102
rect -1581 3068 -1547 3102
rect -1513 3068 -1479 3102
rect -1445 3068 -1411 3102
rect -1377 3068 -1343 3102
rect -1309 3068 -1275 3102
rect -1241 3068 -1207 3102
rect -1173 3068 -1139 3102
rect -1105 3068 -1071 3102
rect -1037 3068 -1003 3102
rect -969 3068 -935 3102
rect -901 3068 -867 3102
rect -833 3068 -799 3102
rect -765 3068 -731 3102
rect -697 3068 -663 3102
rect -629 3068 -595 3102
rect -561 3068 -527 3102
rect -493 3068 -459 3102
rect -425 3068 -391 3102
rect -357 3068 -323 3102
rect -289 3068 -255 3102
rect -221 3068 -187 3102
rect -153 3068 -119 3102
rect -85 3068 -51 3102
rect -17 3068 17 3102
rect 51 3068 85 3102
rect 119 3068 153 3102
rect 187 3068 221 3102
rect 255 3068 289 3102
rect 323 3068 357 3102
rect 391 3068 425 3102
rect 459 3068 493 3102
rect 527 3068 561 3102
rect 595 3068 629 3102
rect 663 3068 697 3102
rect 731 3068 765 3102
rect 799 3068 833 3102
rect 867 3068 901 3102
rect 935 3068 969 3102
rect 1003 3068 1037 3102
rect 1071 3068 1105 3102
rect 1139 3068 1173 3102
rect 1207 3068 1241 3102
rect 1275 3068 1309 3102
rect 1343 3068 1377 3102
rect 1411 3068 1445 3102
rect 1479 3068 1513 3102
rect 1547 3068 1581 3102
rect 1615 3068 1649 3102
rect 1683 3068 1717 3102
rect 1751 3068 1785 3102
rect 1819 3068 1853 3102
rect 1887 3068 1921 3102
rect 1955 3068 1989 3102
rect 2023 3068 2057 3102
rect 2091 3068 2125 3102
rect 2159 3068 2193 3102
rect 2227 3068 2261 3102
rect 2295 3068 2329 3102
rect 2363 3068 2397 3102
rect 2431 3068 2465 3102
rect 2499 3068 2533 3102
rect 2567 3068 2601 3102
rect 2635 3068 2669 3102
rect 2703 3068 2737 3102
rect 2771 3068 2805 3102
rect 2839 3068 2873 3102
rect 2907 3068 2941 3102
rect 2975 3068 3102 3102
rect -3102 2975 -3068 3068
rect -3102 2907 -3068 2941
rect -3102 2839 -3068 2873
rect -3102 2771 -3068 2805
rect -3102 2703 -3068 2737
rect -3102 2635 -3068 2669
rect -3102 2567 -3068 2601
rect -3102 2499 -3068 2533
rect -3102 2431 -3068 2465
rect -3102 2363 -3068 2397
rect -3102 2295 -3068 2329
rect -3102 2227 -3068 2261
rect -3102 2159 -3068 2193
rect -3102 2091 -3068 2125
rect -3102 2023 -3068 2057
rect -3102 1955 -3068 1989
rect -3102 1887 -3068 1921
rect -3102 1819 -3068 1853
rect -3102 1751 -3068 1785
rect -3102 1683 -3068 1717
rect -3102 1615 -3068 1649
rect -3102 1547 -3068 1581
rect -3102 1479 -3068 1513
rect -3102 1411 -3068 1445
rect -3102 1343 -3068 1377
rect -3102 1275 -3068 1309
rect -3102 1207 -3068 1241
rect -3102 1139 -3068 1173
rect -3102 1071 -3068 1105
rect -3102 1003 -3068 1037
rect -3102 935 -3068 969
rect -3102 867 -3068 901
rect -3102 799 -3068 833
rect -3102 731 -3068 765
rect -3102 663 -3068 697
rect -3102 595 -3068 629
rect -3102 527 -3068 561
rect -3102 459 -3068 493
rect -3102 391 -3068 425
rect -3102 323 -3068 357
rect -3102 255 -3068 289
rect -3102 187 -3068 221
rect -3102 119 -3068 153
rect -3102 51 -3068 85
rect -3102 -17 -3068 17
rect -3102 -85 -3068 -51
rect -3102 -153 -3068 -119
rect -3102 -221 -3068 -187
rect -3102 -289 -3068 -255
rect -3102 -357 -3068 -323
rect -3102 -425 -3068 -391
rect -3102 -493 -3068 -459
rect -3102 -561 -3068 -527
rect -3102 -629 -3068 -595
rect -3102 -697 -3068 -663
rect -3102 -765 -3068 -731
rect -3102 -833 -3068 -799
rect -3102 -901 -3068 -867
rect -3102 -969 -3068 -935
rect -3102 -1037 -3068 -1003
rect -3102 -1105 -3068 -1071
rect -3102 -1173 -3068 -1139
rect -3102 -1241 -3068 -1207
rect -3102 -1309 -3068 -1275
rect -3102 -1377 -3068 -1343
rect -3102 -1445 -3068 -1411
rect -3102 -1513 -3068 -1479
rect -3102 -1581 -3068 -1547
rect -3102 -1649 -3068 -1615
rect -3102 -1717 -3068 -1683
rect -3102 -1785 -3068 -1751
rect -3102 -1853 -3068 -1819
rect -3102 -1921 -3068 -1887
rect -3102 -1989 -3068 -1955
rect -3102 -2057 -3068 -2023
rect -3102 -2125 -3068 -2091
rect -3102 -2193 -3068 -2159
rect -3102 -2261 -3068 -2227
rect -3102 -2329 -3068 -2295
rect -3102 -2397 -3068 -2363
rect -3102 -2465 -3068 -2431
rect -3102 -2533 -3068 -2499
rect -3102 -2601 -3068 -2567
rect -3102 -2669 -3068 -2635
rect -3102 -2737 -3068 -2703
rect -3102 -2805 -3068 -2771
rect -3102 -2873 -3068 -2839
rect -3102 -2941 -3068 -2907
rect -3102 -3068 -3068 -2975
rect -3004 2975 3004 2988
rect -3004 -2975 -2975 2975
rect 2975 -2975 3004 2975
rect -3004 -2988 3004 -2975
rect 3068 2975 3102 3068
rect 3068 2907 3102 2941
rect 3068 2839 3102 2873
rect 3068 2771 3102 2805
rect 3068 2703 3102 2737
rect 3068 2635 3102 2669
rect 3068 2567 3102 2601
rect 3068 2499 3102 2533
rect 3068 2431 3102 2465
rect 3068 2363 3102 2397
rect 3068 2295 3102 2329
rect 3068 2227 3102 2261
rect 3068 2159 3102 2193
rect 3068 2091 3102 2125
rect 3068 2023 3102 2057
rect 3068 1955 3102 1989
rect 3068 1887 3102 1921
rect 3068 1819 3102 1853
rect 3068 1751 3102 1785
rect 3068 1683 3102 1717
rect 3068 1615 3102 1649
rect 3068 1547 3102 1581
rect 3068 1479 3102 1513
rect 3068 1411 3102 1445
rect 3068 1343 3102 1377
rect 3068 1275 3102 1309
rect 3068 1207 3102 1241
rect 3068 1139 3102 1173
rect 3068 1071 3102 1105
rect 3068 1003 3102 1037
rect 3068 935 3102 969
rect 3068 867 3102 901
rect 3068 799 3102 833
rect 3068 731 3102 765
rect 3068 663 3102 697
rect 3068 595 3102 629
rect 3068 527 3102 561
rect 3068 459 3102 493
rect 3068 391 3102 425
rect 3068 323 3102 357
rect 3068 255 3102 289
rect 3068 187 3102 221
rect 3068 119 3102 153
rect 3068 51 3102 85
rect 3068 -17 3102 17
rect 3068 -85 3102 -51
rect 3068 -153 3102 -119
rect 3068 -221 3102 -187
rect 3068 -289 3102 -255
rect 3068 -357 3102 -323
rect 3068 -425 3102 -391
rect 3068 -493 3102 -459
rect 3068 -561 3102 -527
rect 3068 -629 3102 -595
rect 3068 -697 3102 -663
rect 3068 -765 3102 -731
rect 3068 -833 3102 -799
rect 3068 -901 3102 -867
rect 3068 -969 3102 -935
rect 3068 -1037 3102 -1003
rect 3068 -1105 3102 -1071
rect 3068 -1173 3102 -1139
rect 3068 -1241 3102 -1207
rect 3068 -1309 3102 -1275
rect 3068 -1377 3102 -1343
rect 3068 -1445 3102 -1411
rect 3068 -1513 3102 -1479
rect 3068 -1581 3102 -1547
rect 3068 -1649 3102 -1615
rect 3068 -1717 3102 -1683
rect 3068 -1785 3102 -1751
rect 3068 -1853 3102 -1819
rect 3068 -1921 3102 -1887
rect 3068 -1989 3102 -1955
rect 3068 -2057 3102 -2023
rect 3068 -2125 3102 -2091
rect 3068 -2193 3102 -2159
rect 3068 -2261 3102 -2227
rect 3068 -2329 3102 -2295
rect 3068 -2397 3102 -2363
rect 3068 -2465 3102 -2431
rect 3068 -2533 3102 -2499
rect 3068 -2601 3102 -2567
rect 3068 -2669 3102 -2635
rect 3068 -2737 3102 -2703
rect 3068 -2805 3102 -2771
rect 3068 -2873 3102 -2839
rect 3068 -2941 3102 -2907
rect 3068 -3068 3102 -2975
rect -3102 -3102 -2975 -3068
rect -2941 -3102 -2907 -3068
rect -2873 -3102 -2839 -3068
rect -2805 -3102 -2771 -3068
rect -2737 -3102 -2703 -3068
rect -2669 -3102 -2635 -3068
rect -2601 -3102 -2567 -3068
rect -2533 -3102 -2499 -3068
rect -2465 -3102 -2431 -3068
rect -2397 -3102 -2363 -3068
rect -2329 -3102 -2295 -3068
rect -2261 -3102 -2227 -3068
rect -2193 -3102 -2159 -3068
rect -2125 -3102 -2091 -3068
rect -2057 -3102 -2023 -3068
rect -1989 -3102 -1955 -3068
rect -1921 -3102 -1887 -3068
rect -1853 -3102 -1819 -3068
rect -1785 -3102 -1751 -3068
rect -1717 -3102 -1683 -3068
rect -1649 -3102 -1615 -3068
rect -1581 -3102 -1547 -3068
rect -1513 -3102 -1479 -3068
rect -1445 -3102 -1411 -3068
rect -1377 -3102 -1343 -3068
rect -1309 -3102 -1275 -3068
rect -1241 -3102 -1207 -3068
rect -1173 -3102 -1139 -3068
rect -1105 -3102 -1071 -3068
rect -1037 -3102 -1003 -3068
rect -969 -3102 -935 -3068
rect -901 -3102 -867 -3068
rect -833 -3102 -799 -3068
rect -765 -3102 -731 -3068
rect -697 -3102 -663 -3068
rect -629 -3102 -595 -3068
rect -561 -3102 -527 -3068
rect -493 -3102 -459 -3068
rect -425 -3102 -391 -3068
rect -357 -3102 -323 -3068
rect -289 -3102 -255 -3068
rect -221 -3102 -187 -3068
rect -153 -3102 -119 -3068
rect -85 -3102 -51 -3068
rect -17 -3102 17 -3068
rect 51 -3102 85 -3068
rect 119 -3102 153 -3068
rect 187 -3102 221 -3068
rect 255 -3102 289 -3068
rect 323 -3102 357 -3068
rect 391 -3102 425 -3068
rect 459 -3102 493 -3068
rect 527 -3102 561 -3068
rect 595 -3102 629 -3068
rect 663 -3102 697 -3068
rect 731 -3102 765 -3068
rect 799 -3102 833 -3068
rect 867 -3102 901 -3068
rect 935 -3102 969 -3068
rect 1003 -3102 1037 -3068
rect 1071 -3102 1105 -3068
rect 1139 -3102 1173 -3068
rect 1207 -3102 1241 -3068
rect 1275 -3102 1309 -3068
rect 1343 -3102 1377 -3068
rect 1411 -3102 1445 -3068
rect 1479 -3102 1513 -3068
rect 1547 -3102 1581 -3068
rect 1615 -3102 1649 -3068
rect 1683 -3102 1717 -3068
rect 1751 -3102 1785 -3068
rect 1819 -3102 1853 -3068
rect 1887 -3102 1921 -3068
rect 1955 -3102 1989 -3068
rect 2023 -3102 2057 -3068
rect 2091 -3102 2125 -3068
rect 2159 -3102 2193 -3068
rect 2227 -3102 2261 -3068
rect 2295 -3102 2329 -3068
rect 2363 -3102 2397 -3068
rect 2431 -3102 2465 -3068
rect 2499 -3102 2533 -3068
rect 2567 -3102 2601 -3068
rect 2635 -3102 2669 -3068
rect 2703 -3102 2737 -3068
rect 2771 -3102 2805 -3068
rect 2839 -3102 2873 -3068
rect 2907 -3102 2941 -3068
rect 2975 -3102 3102 -3068
rect 3206 3043 3240 3077
rect 3206 2975 3240 3009
rect 3206 2907 3240 2941
rect 3206 2839 3240 2873
rect 3206 2771 3240 2805
rect 3206 2703 3240 2737
rect 3206 2635 3240 2669
rect 3206 2567 3240 2601
rect 3206 2499 3240 2533
rect 3206 2431 3240 2465
rect 3206 2363 3240 2397
rect 3206 2295 3240 2329
rect 3206 2227 3240 2261
rect 3206 2159 3240 2193
rect 3206 2091 3240 2125
rect 3206 2023 3240 2057
rect 3206 1955 3240 1989
rect 3206 1887 3240 1921
rect 3206 1819 3240 1853
rect 3206 1751 3240 1785
rect 3206 1683 3240 1717
rect 3206 1615 3240 1649
rect 3206 1547 3240 1581
rect 3206 1479 3240 1513
rect 3206 1411 3240 1445
rect 3206 1343 3240 1377
rect 3206 1275 3240 1309
rect 3206 1207 3240 1241
rect 3206 1139 3240 1173
rect 3206 1071 3240 1105
rect 3206 1003 3240 1037
rect 3206 935 3240 969
rect 3206 867 3240 901
rect 3206 799 3240 833
rect 3206 731 3240 765
rect 3206 663 3240 697
rect 3206 595 3240 629
rect 3206 527 3240 561
rect 3206 459 3240 493
rect 3206 391 3240 425
rect 3206 323 3240 357
rect 3206 255 3240 289
rect 3206 187 3240 221
rect 3206 119 3240 153
rect 3206 51 3240 85
rect 3206 -17 3240 17
rect 3206 -85 3240 -51
rect 3206 -153 3240 -119
rect 3206 -221 3240 -187
rect 3206 -289 3240 -255
rect 3206 -357 3240 -323
rect 3206 -425 3240 -391
rect 3206 -493 3240 -459
rect 3206 -561 3240 -527
rect 3206 -629 3240 -595
rect 3206 -697 3240 -663
rect 3206 -765 3240 -731
rect 3206 -833 3240 -799
rect 3206 -901 3240 -867
rect 3206 -969 3240 -935
rect 3206 -1037 3240 -1003
rect 3206 -1105 3240 -1071
rect 3206 -1173 3240 -1139
rect 3206 -1241 3240 -1207
rect 3206 -1309 3240 -1275
rect 3206 -1377 3240 -1343
rect 3206 -1445 3240 -1411
rect 3206 -1513 3240 -1479
rect 3206 -1581 3240 -1547
rect 3206 -1649 3240 -1615
rect 3206 -1717 3240 -1683
rect 3206 -1785 3240 -1751
rect 3206 -1853 3240 -1819
rect 3206 -1921 3240 -1887
rect 3206 -1989 3240 -1955
rect 3206 -2057 3240 -2023
rect 3206 -2125 3240 -2091
rect 3206 -2193 3240 -2159
rect 3206 -2261 3240 -2227
rect 3206 -2329 3240 -2295
rect 3206 -2397 3240 -2363
rect 3206 -2465 3240 -2431
rect 3206 -2533 3240 -2499
rect 3206 -2601 3240 -2567
rect 3206 -2669 3240 -2635
rect 3206 -2737 3240 -2703
rect 3206 -2805 3240 -2771
rect 3206 -2873 3240 -2839
rect 3206 -2941 3240 -2907
rect 3206 -3009 3240 -2975
rect 3206 -3077 3240 -3043
rect -3240 -3206 -3206 -3111
rect 3206 -3206 3240 -3111
rect -3240 -3240 -3111 -3206
rect -3077 -3240 -3043 -3206
rect -3009 -3240 -2975 -3206
rect -2941 -3240 -2907 -3206
rect -2873 -3240 -2839 -3206
rect -2805 -3240 -2771 -3206
rect -2737 -3240 -2703 -3206
rect -2669 -3240 -2635 -3206
rect -2601 -3240 -2567 -3206
rect -2533 -3240 -2499 -3206
rect -2465 -3240 -2431 -3206
rect -2397 -3240 -2363 -3206
rect -2329 -3240 -2295 -3206
rect -2261 -3240 -2227 -3206
rect -2193 -3240 -2159 -3206
rect -2125 -3240 -2091 -3206
rect -2057 -3240 -2023 -3206
rect -1989 -3240 -1955 -3206
rect -1921 -3240 -1887 -3206
rect -1853 -3240 -1819 -3206
rect -1785 -3240 -1751 -3206
rect -1717 -3240 -1683 -3206
rect -1649 -3240 -1615 -3206
rect -1581 -3240 -1547 -3206
rect -1513 -3240 -1479 -3206
rect -1445 -3240 -1411 -3206
rect -1377 -3240 -1343 -3206
rect -1309 -3240 -1275 -3206
rect -1241 -3240 -1207 -3206
rect -1173 -3240 -1139 -3206
rect -1105 -3240 -1071 -3206
rect -1037 -3240 -1003 -3206
rect -969 -3240 -935 -3206
rect -901 -3240 -867 -3206
rect -833 -3240 -799 -3206
rect -765 -3240 -731 -3206
rect -697 -3240 -663 -3206
rect -629 -3240 -595 -3206
rect -561 -3240 -527 -3206
rect -493 -3240 -459 -3206
rect -425 -3240 -391 -3206
rect -357 -3240 -323 -3206
rect -289 -3240 -255 -3206
rect -221 -3240 -187 -3206
rect -153 -3240 -119 -3206
rect -85 -3240 -51 -3206
rect -17 -3240 17 -3206
rect 51 -3240 85 -3206
rect 119 -3240 153 -3206
rect 187 -3240 221 -3206
rect 255 -3240 289 -3206
rect 323 -3240 357 -3206
rect 391 -3240 425 -3206
rect 459 -3240 493 -3206
rect 527 -3240 561 -3206
rect 595 -3240 629 -3206
rect 663 -3240 697 -3206
rect 731 -3240 765 -3206
rect 799 -3240 833 -3206
rect 867 -3240 901 -3206
rect 935 -3240 969 -3206
rect 1003 -3240 1037 -3206
rect 1071 -3240 1105 -3206
rect 1139 -3240 1173 -3206
rect 1207 -3240 1241 -3206
rect 1275 -3240 1309 -3206
rect 1343 -3240 1377 -3206
rect 1411 -3240 1445 -3206
rect 1479 -3240 1513 -3206
rect 1547 -3240 1581 -3206
rect 1615 -3240 1649 -3206
rect 1683 -3240 1717 -3206
rect 1751 -3240 1785 -3206
rect 1819 -3240 1853 -3206
rect 1887 -3240 1921 -3206
rect 1955 -3240 1989 -3206
rect 2023 -3240 2057 -3206
rect 2091 -3240 2125 -3206
rect 2159 -3240 2193 -3206
rect 2227 -3240 2261 -3206
rect 2295 -3240 2329 -3206
rect 2363 -3240 2397 -3206
rect 2431 -3240 2465 -3206
rect 2499 -3240 2533 -3206
rect 2567 -3240 2601 -3206
rect 2635 -3240 2669 -3206
rect 2703 -3240 2737 -3206
rect 2771 -3240 2805 -3206
rect 2839 -3240 2873 -3206
rect 2907 -3240 2941 -3206
rect 2975 -3240 3009 -3206
rect 3043 -3240 3077 -3206
rect 3111 -3240 3240 -3206
<< viali >>
rect -2969 -2969 2969 2969
<< metal1 >>
rect -3000 2969 3000 2994
rect -3000 -2969 -2969 2969
rect 2969 -2969 3000 2969
rect -3000 -2994 3000 -2969
<< properties >>
string FIXED_BBOX -3084 -3084 3084 3084
<< end >>
