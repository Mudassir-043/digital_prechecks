magic
tech sky130B
magscale 1 2
timestamp 1667586985
<< metal4 >>
rect -1349 3039 1349 3080
rect -1349 -3039 1093 3039
rect 1329 -3039 1349 3039
rect -1349 -3080 1349 -3039
<< via4 >>
rect 1093 -3039 1329 3039
<< mimcap2 >>
rect -1269 2960 731 3000
rect -1269 -2960 -1229 2960
rect 691 -2960 731 2960
rect -1269 -3000 731 -2960
<< mimcap2contact >>
rect -1229 -2960 691 2960
<< metal5 >>
rect 1051 3039 1371 3081
rect -1253 2960 715 2984
rect -1253 -2960 -1229 2960
rect 691 -2960 715 2960
rect -1253 -2984 715 -2960
rect 1051 -3039 1093 3039
rect 1329 -3039 1371 3039
rect 1051 -3081 1371 -3039
<< properties >>
string FIXED_BBOX -1349 -3080 811 3080
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 10 l 30 val 615.2 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
