magic
tech sky130B
timestamp 1667596055
<< pwell >>
rect -2069 -2069 2069 2069
<< psubdiff >>
rect -2051 2034 -2003 2051
rect 2003 2034 2051 2051
rect -2051 2003 -2034 2034
rect 2034 2003 2051 2034
rect -2051 -2034 -2034 -2003
rect 2034 -2034 2051 -2003
rect -2051 -2051 -2003 -2034
rect 2003 -2051 2051 -2034
<< psubdiffcont >>
rect -2003 2034 2003 2051
rect -2051 -2003 -2034 2003
rect 2034 -2003 2051 2003
rect -2003 -2051 2003 -2034
<< ndiode >>
rect -2000 1994 2000 2000
rect -2000 -1994 -1994 1994
rect 1994 -1994 2000 1994
rect -2000 -2000 2000 -1994
<< ndiodec >>
rect -1994 -1994 1994 1994
<< locali >>
rect -2051 2034 -2003 2051
rect 2003 2034 2051 2051
rect -2051 2003 -2034 2034
rect 2034 2003 2051 2034
rect -2002 -1994 -1994 1994
rect 1994 -1994 2002 1994
rect -2051 -2034 -2034 -2003
rect 2034 -2034 2051 -2003
rect -2051 -2051 -2003 -2034
rect 2003 -2051 2051 -2034
<< viali >>
rect -1994 -1994 1994 1994
<< metal1 >>
rect -2000 1994 2000 1997
rect -2000 -1994 -1994 1994
rect 1994 -1994 2000 1994
rect -2000 -1997 2000 -1994
<< properties >>
string FIXED_BBOX -2042 -2042 2042 2042
string gencell sky130_fd_pr__diode_pw2nd_05v5
string library sky130
string parameters w 40 l 40 area 1.6k peri 160.0 nx 1 ny 1 dummy 0 lmin 0.45 wmin 0.45 elc 1 erc 1 etc 1 ebc 1 doverlap 0 compatible {sky130_fd_pr__diode_pw2nd_05v5 sky130_fd_pr__diode_pw2nd_05v5_lvt  sky130_fd_pr__diode_pw2nd_05v5_nvt sky130_fd_pr__diode_pw2nd_11v0} full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
