magic
tech sky130B
timestamp 1667595866
<< pwell >>
rect -1069 -1069 1069 1069
<< psubdiff >>
rect -1051 1034 -1003 1051
rect 1003 1034 1051 1051
rect -1051 1003 -1034 1034
rect 1034 1003 1051 1034
rect -1051 -1034 -1034 -1003
rect 1034 -1034 1051 -1003
rect -1051 -1051 -1003 -1034
rect 1003 -1051 1051 -1034
<< psubdiffcont >>
rect -1003 1034 1003 1051
rect -1051 -1003 -1034 1003
rect 1034 -1003 1051 1003
rect -1003 -1051 1003 -1034
<< ndiode >>
rect -1000 994 1000 1000
rect -1000 -994 -994 994
rect 994 -994 1000 994
rect -1000 -1000 1000 -994
<< ndiodec >>
rect -994 -994 994 994
<< locali >>
rect -1051 1034 -1003 1051
rect 1003 1034 1051 1051
rect -1051 1003 -1034 1034
rect 1034 1003 1051 1034
rect -1002 -994 -994 994
rect 994 -994 1002 994
rect -1051 -1034 -1034 -1003
rect 1034 -1034 1051 -1003
rect -1051 -1051 -1003 -1034
rect 1003 -1051 1051 -1034
<< viali >>
rect -994 -994 994 994
<< metal1 >>
rect -1000 994 1000 997
rect -1000 -994 -994 994
rect 994 -994 1000 994
rect -1000 -997 1000 -994
<< properties >>
string FIXED_BBOX -1042 -1042 1042 1042
string gencell sky130_fd_pr__diode_pw2nd_05v5
string library sky130
string parameters w 20 l 20 area 400.0 peri 80.0 nx 1 ny 1 dummy 0 lmin 0.45 wmin 0.45 elc 1 erc 1 etc 1 ebc 1 doverlap 0 compatible {sky130_fd_pr__diode_pw2nd_05v5 sky130_fd_pr__diode_pw2nd_05v5_lvt  sky130_fd_pr__diode_pw2nd_05v5_nvt sky130_fd_pr__diode_pw2nd_11v0} full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
